magic
tech gf180mcuD
magscale 1 5
timestamp 1702149601
<< obsm1 >>
rect 672 1538 19400 18633
<< metal2 >>
rect 9072 19600 9128 20000
rect 9408 19600 9464 20000
rect 9744 19600 9800 20000
rect 10080 19600 10136 20000
rect 10416 19600 10472 20000
rect 10752 19600 10808 20000
rect 11088 19600 11144 20000
rect 11424 19600 11480 20000
rect 11760 19600 11816 20000
rect 12096 19600 12152 20000
rect 12432 19600 12488 20000
rect 12768 19600 12824 20000
rect 13104 19600 13160 20000
rect 13440 19600 13496 20000
rect 13776 19600 13832 20000
rect 14112 19600 14168 20000
rect 14448 19600 14504 20000
rect 14784 19600 14840 20000
rect 15120 19600 15176 20000
rect 15456 19600 15512 20000
rect 15792 19600 15848 20000
rect 16128 19600 16184 20000
rect 16464 19600 16520 20000
rect 16800 19600 16856 20000
rect 17136 19600 17192 20000
rect 17472 19600 17528 20000
rect 17808 19600 17864 20000
rect 18144 19600 18200 20000
rect 18480 19600 18536 20000
rect 18816 19600 18872 20000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
rect 13104 0 13160 400
rect 13440 0 13496 400
rect 13776 0 13832 400
rect 14112 0 14168 400
rect 14448 0 14504 400
rect 14784 0 14840 400
rect 15120 0 15176 400
rect 15456 0 15512 400
rect 15792 0 15848 400
rect 16128 0 16184 400
rect 16464 0 16520 400
rect 16800 0 16856 400
rect 17136 0 17192 400
rect 17472 0 17528 400
rect 17808 0 17864 400
rect 18144 0 18200 400
rect 18480 0 18536 400
rect 18816 0 18872 400
rect 19152 0 19208 400
rect 19488 0 19544 400
rect 19824 0 19880 400
<< obsm2 >>
rect 742 19570 9042 19871
rect 9158 19570 9378 19871
rect 9494 19570 9714 19871
rect 9830 19570 10050 19871
rect 10166 19570 10386 19871
rect 10502 19570 10722 19871
rect 10838 19570 11058 19871
rect 11174 19570 11394 19871
rect 11510 19570 11730 19871
rect 11846 19570 12066 19871
rect 12182 19570 12402 19871
rect 12518 19570 12738 19871
rect 12854 19570 13074 19871
rect 13190 19570 13410 19871
rect 13526 19570 13746 19871
rect 13862 19570 14082 19871
rect 14198 19570 14418 19871
rect 14534 19570 14754 19871
rect 14870 19570 15090 19871
rect 15206 19570 15426 19871
rect 15542 19570 15762 19871
rect 15878 19570 16098 19871
rect 16214 19570 16434 19871
rect 16550 19570 16770 19871
rect 16886 19570 17106 19871
rect 17222 19570 17442 19871
rect 17558 19570 17778 19871
rect 17894 19570 18114 19871
rect 18230 19570 18450 19871
rect 18566 19570 18786 19871
rect 18902 19570 19866 19871
rect 742 430 19866 19570
rect 758 9 978 430
rect 1094 9 1314 430
rect 1430 9 1650 430
rect 1766 9 1986 430
rect 2102 9 2322 430
rect 2438 9 2658 430
rect 2774 9 2994 430
rect 3110 9 3330 430
rect 3446 9 3666 430
rect 3782 9 4002 430
rect 4118 9 4338 430
rect 4454 9 4674 430
rect 4790 9 5010 430
rect 5126 9 5346 430
rect 5462 9 5682 430
rect 5798 9 6018 430
rect 6134 9 6354 430
rect 6470 9 6690 430
rect 6806 9 7026 430
rect 7142 9 7362 430
rect 7478 9 7698 430
rect 7814 9 8034 430
rect 8150 9 8370 430
rect 8486 9 8706 430
rect 8822 9 9042 430
rect 9158 9 9378 430
rect 9494 9 9714 430
rect 9830 9 10050 430
rect 10166 9 10386 430
rect 10502 9 10722 430
rect 10838 9 11058 430
rect 11174 9 11394 430
rect 11510 9 11730 430
rect 11846 9 12066 430
rect 12182 9 12402 430
rect 12518 9 12738 430
rect 12854 9 13074 430
rect 13190 9 13410 430
rect 13526 9 13746 430
rect 13862 9 14082 430
rect 14198 9 14418 430
rect 14534 9 14754 430
rect 14870 9 15090 430
rect 15206 9 15426 430
rect 15542 9 15762 430
rect 15878 9 16098 430
rect 16214 9 16434 430
rect 16550 9 16770 430
rect 16886 9 17106 430
rect 17222 9 17442 430
rect 17558 9 17778 430
rect 17894 9 18114 430
rect 18230 9 18450 430
rect 18566 9 18786 430
rect 18902 9 19122 430
rect 19238 9 19458 430
rect 19574 9 19794 430
<< metal3 >>
rect 19600 19824 20000 19880
rect 19600 19488 20000 19544
rect 19600 19152 20000 19208
rect 19600 18816 20000 18872
rect 19600 18480 20000 18536
rect 19600 18144 20000 18200
rect 19600 17808 20000 17864
rect 19600 17472 20000 17528
rect 19600 17136 20000 17192
rect 19600 16800 20000 16856
rect 19600 16464 20000 16520
rect 19600 16128 20000 16184
rect 19600 15792 20000 15848
rect 19600 15456 20000 15512
rect 19600 15120 20000 15176
rect 19600 14784 20000 14840
rect 19600 14448 20000 14504
rect 19600 14112 20000 14168
rect 19600 13776 20000 13832
rect 19600 13440 20000 13496
rect 0 13104 400 13160
rect 19600 13104 20000 13160
rect 19600 12768 20000 12824
rect 19600 8400 20000 8456
rect 19600 8064 20000 8120
rect 19600 7728 20000 7784
rect 0 7392 400 7448
rect 19600 7392 20000 7448
rect 19600 7056 20000 7112
rect 19600 6720 20000 6776
rect 19600 6384 20000 6440
rect 19600 6048 20000 6104
rect 19600 5712 20000 5768
rect 19600 5376 20000 5432
rect 19600 5040 20000 5096
rect 19600 4704 20000 4760
rect 19600 4368 20000 4424
rect 19600 4032 20000 4088
rect 19600 3696 20000 3752
rect 19600 3360 20000 3416
rect 19600 3024 20000 3080
rect 19600 2688 20000 2744
rect 19600 2352 20000 2408
rect 19600 2016 20000 2072
rect 19600 1680 20000 1736
rect 19600 1344 20000 1400
rect 19600 1008 20000 1064
rect 19600 672 20000 728
rect 19600 336 20000 392
rect 19600 0 20000 56
<< obsm3 >>
rect 400 19794 19570 19866
rect 400 19574 19871 19794
rect 400 19458 19570 19574
rect 400 19238 19871 19458
rect 400 19122 19570 19238
rect 400 18902 19871 19122
rect 400 18786 19570 18902
rect 400 18566 19871 18786
rect 400 18450 19570 18566
rect 400 18230 19871 18450
rect 400 18114 19570 18230
rect 400 17894 19871 18114
rect 400 17778 19570 17894
rect 400 17558 19871 17778
rect 400 17442 19570 17558
rect 400 17222 19871 17442
rect 400 17106 19570 17222
rect 400 16886 19871 17106
rect 400 16770 19570 16886
rect 400 16550 19871 16770
rect 400 16434 19570 16550
rect 400 16214 19871 16434
rect 400 16098 19570 16214
rect 400 15878 19871 16098
rect 400 15762 19570 15878
rect 400 15542 19871 15762
rect 400 15426 19570 15542
rect 400 15206 19871 15426
rect 400 15090 19570 15206
rect 400 14870 19871 15090
rect 400 14754 19570 14870
rect 400 14534 19871 14754
rect 400 14418 19570 14534
rect 400 14198 19871 14418
rect 400 14082 19570 14198
rect 400 13862 19871 14082
rect 400 13746 19570 13862
rect 400 13526 19871 13746
rect 400 13410 19570 13526
rect 400 13190 19871 13410
rect 430 13074 19570 13190
rect 400 12854 19871 13074
rect 400 12738 19570 12854
rect 400 8486 19871 12738
rect 400 8370 19570 8486
rect 400 8150 19871 8370
rect 400 8034 19570 8150
rect 400 7814 19871 8034
rect 400 7698 19570 7814
rect 400 7478 19871 7698
rect 430 7362 19570 7478
rect 400 7142 19871 7362
rect 400 7026 19570 7142
rect 400 6806 19871 7026
rect 400 6690 19570 6806
rect 400 6470 19871 6690
rect 400 6354 19570 6470
rect 400 6134 19871 6354
rect 400 6018 19570 6134
rect 400 5798 19871 6018
rect 400 5682 19570 5798
rect 400 5462 19871 5682
rect 400 5346 19570 5462
rect 400 5126 19871 5346
rect 400 5010 19570 5126
rect 400 4790 19871 5010
rect 400 4674 19570 4790
rect 400 4454 19871 4674
rect 400 4338 19570 4454
rect 400 4118 19871 4338
rect 400 4002 19570 4118
rect 400 3782 19871 4002
rect 400 3666 19570 3782
rect 400 3446 19871 3666
rect 400 3330 19570 3446
rect 400 3110 19871 3330
rect 400 2994 19570 3110
rect 400 2774 19871 2994
rect 400 2658 19570 2774
rect 400 2438 19871 2658
rect 400 2322 19570 2438
rect 400 2102 19871 2322
rect 400 1986 19570 2102
rect 400 1766 19871 1986
rect 400 1650 19570 1766
rect 400 1430 19871 1650
rect 400 1314 19570 1430
rect 400 1094 19871 1314
rect 400 978 19570 1094
rect 400 758 19871 978
rect 400 642 19570 758
rect 400 422 19871 642
rect 400 306 19570 422
rect 400 86 19871 306
rect 400 14 19570 86
<< metal4 >>
rect 2923 1538 3083 18454
rect 5254 1538 5414 18454
rect 7585 1538 7745 18454
rect 9916 1538 10076 18454
rect 12247 1538 12407 18454
rect 14578 1538 14738 18454
rect 16909 1538 17069 18454
rect 19240 1538 19400 18454
<< obsm4 >>
rect 14854 1508 16879 8335
rect 17099 1508 17626 8335
rect 14854 1017 17626 1508
<< labels >>
rlabel metal2 s 1008 0 1064 400 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
rlabel metal2 s 672 0 728 400 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 2 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 3 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 4 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 5 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 6 nsew signal input
rlabel metal3 s 0 7392 400 7448 6 ccff_head
port 7 nsew signal input
rlabel metal3 s 19600 8400 20000 8456 6 ccff_tail
port 8 nsew signal output
rlabel metal2 s 3024 0 3080 400 6 chanx_left_in[0]
port 9 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 chanx_left_in[10]
port 10 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 chanx_left_in[11]
port 11 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 chanx_left_in[12]
port 12 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 chanx_left_in[13]
port 13 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 chanx_left_in[14]
port 14 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 chanx_left_in[15]
port 15 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 chanx_left_in[16]
port 16 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 chanx_left_in[17]
port 17 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 chanx_left_in[18]
port 18 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 chanx_left_in[19]
port 19 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 chanx_left_in[1]
port 20 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 chanx_left_in[2]
port 21 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 chanx_left_in[3]
port 22 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 chanx_left_in[4]
port 23 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 chanx_left_in[5]
port 24 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 chanx_left_in[6]
port 25 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 chanx_left_in[7]
port 26 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 chanx_left_in[8]
port 27 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 chanx_left_in[9]
port 28 nsew signal input
rlabel metal2 s 13104 19600 13160 20000 6 chanx_left_out[0]
port 29 nsew signal output
rlabel metal2 s 18816 19600 18872 20000 6 chanx_left_out[10]
port 30 nsew signal output
rlabel metal2 s 18144 19600 18200 20000 6 chanx_left_out[11]
port 31 nsew signal output
rlabel metal2 s 17472 19600 17528 20000 6 chanx_left_out[12]
port 32 nsew signal output
rlabel metal3 s 19600 0 20000 56 6 chanx_left_out[13]
port 33 nsew signal output
rlabel metal3 s 19600 12768 20000 12824 6 chanx_left_out[14]
port 34 nsew signal output
rlabel metal2 s 14448 19600 14504 20000 6 chanx_left_out[15]
port 35 nsew signal output
rlabel metal2 s 19824 0 19880 400 6 chanx_left_out[16]
port 36 nsew signal output
rlabel metal3 s 19600 5712 20000 5768 6 chanx_left_out[17]
port 37 nsew signal output
rlabel metal3 s 19600 19824 20000 19880 6 chanx_left_out[18]
port 38 nsew signal output
rlabel metal2 s 16464 19600 16520 20000 6 chanx_left_out[19]
port 39 nsew signal output
rlabel metal3 s 19600 16800 20000 16856 6 chanx_left_out[1]
port 40 nsew signal output
rlabel metal2 s 15792 19600 15848 20000 6 chanx_left_out[2]
port 41 nsew signal output
rlabel metal3 s 19600 2016 20000 2072 6 chanx_left_out[3]
port 42 nsew signal output
rlabel metal2 s 13440 0 13496 400 6 chanx_left_out[4]
port 43 nsew signal output
rlabel metal2 s 17136 19600 17192 20000 6 chanx_left_out[5]
port 44 nsew signal output
rlabel metal3 s 19600 16464 20000 16520 6 chanx_left_out[6]
port 45 nsew signal output
rlabel metal3 s 19600 1680 20000 1736 6 chanx_left_out[7]
port 46 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 chanx_left_out[8]
port 47 nsew signal output
rlabel metal2 s 16800 19600 16856 20000 6 chanx_left_out[9]
port 48 nsew signal output
rlabel metal3 s 19600 13776 20000 13832 6 chany_bottom_in[0]
port 49 nsew signal input
rlabel metal2 s 14112 19600 14168 20000 6 chany_bottom_in[10]
port 50 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 chany_bottom_in[11]
port 51 nsew signal input
rlabel metal2 s 12096 19600 12152 20000 6 chany_bottom_in[12]
port 52 nsew signal input
rlabel metal3 s 19600 1008 20000 1064 6 chany_bottom_in[13]
port 53 nsew signal input
rlabel metal2 s 18480 19600 18536 20000 6 chany_bottom_in[14]
port 54 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 chany_bottom_in[15]
port 55 nsew signal input
rlabel metal2 s 11760 19600 11816 20000 6 chany_bottom_in[16]
port 56 nsew signal input
rlabel metal2 s 9072 19600 9128 20000 6 chany_bottom_in[17]
port 57 nsew signal input
rlabel metal3 s 19600 2688 20000 2744 6 chany_bottom_in[18]
port 58 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 chany_bottom_in[19]
port 59 nsew signal input
rlabel metal3 s 19600 13440 20000 13496 6 chany_bottom_in[1]
port 60 nsew signal input
rlabel metal3 s 19600 14112 20000 14168 6 chany_bottom_in[2]
port 61 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 chany_bottom_in[3]
port 62 nsew signal input
rlabel metal3 s 19600 672 20000 728 6 chany_bottom_in[4]
port 63 nsew signal input
rlabel metal3 s 19600 4368 20000 4424 6 chany_bottom_in[5]
port 64 nsew signal input
rlabel metal3 s 19600 336 20000 392 6 chany_bottom_in[6]
port 65 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 chany_bottom_in[7]
port 66 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 chany_bottom_in[8]
port 67 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 chany_bottom_in[9]
port 68 nsew signal input
rlabel metal3 s 19600 17136 20000 17192 6 chany_bottom_out[0]
port 69 nsew signal output
rlabel metal2 s 15792 0 15848 400 6 chany_bottom_out[10]
port 70 nsew signal output
rlabel metal3 s 19600 13104 20000 13160 6 chany_bottom_out[11]
port 71 nsew signal output
rlabel metal2 s 14784 19600 14840 20000 6 chany_bottom_out[12]
port 72 nsew signal output
rlabel metal2 s 16800 0 16856 400 6 chany_bottom_out[13]
port 73 nsew signal output
rlabel metal3 s 19600 4704 20000 4760 6 chany_bottom_out[14]
port 74 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 chany_bottom_out[15]
port 75 nsew signal output
rlabel metal2 s 10752 19600 10808 20000 6 chany_bottom_out[16]
port 76 nsew signal output
rlabel metal2 s 15456 19600 15512 20000 6 chany_bottom_out[17]
port 77 nsew signal output
rlabel metal3 s 19600 19152 20000 19208 6 chany_bottom_out[18]
port 78 nsew signal output
rlabel metal2 s 10416 19600 10472 20000 6 chany_bottom_out[19]
port 79 nsew signal output
rlabel metal2 s 14112 0 14168 400 6 chany_bottom_out[1]
port 80 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 chany_bottom_out[2]
port 81 nsew signal output
rlabel metal2 s 11088 19600 11144 20000 6 chany_bottom_out[3]
port 82 nsew signal output
rlabel metal3 s 19600 16128 20000 16184 6 chany_bottom_out[4]
port 83 nsew signal output
rlabel metal2 s 14784 0 14840 400 6 chany_bottom_out[5]
port 84 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 chany_bottom_out[6]
port 85 nsew signal output
rlabel metal2 s 12432 19600 12488 20000 6 chany_bottom_out[7]
port 86 nsew signal output
rlabel metal3 s 19600 1344 20000 1400 6 chany_bottom_out[8]
port 87 nsew signal output
rlabel metal3 s 19600 18480 20000 18536 6 chany_bottom_out[9]
port 88 nsew signal output
rlabel metal2 s 13776 0 13832 400 6 chany_top_in[0]
port 89 nsew signal input
rlabel metal3 s 19600 14784 20000 14840 6 chany_top_in[10]
port 90 nsew signal input
rlabel metal3 s 19600 18816 20000 18872 6 chany_top_in[11]
port 91 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 chany_top_in[12]
port 92 nsew signal input
rlabel metal3 s 19600 5376 20000 5432 6 chany_top_in[13]
port 93 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 chany_top_in[14]
port 94 nsew signal input
rlabel metal3 s 19600 3360 20000 3416 6 chany_top_in[15]
port 95 nsew signal input
rlabel metal2 s 15120 19600 15176 20000 6 chany_top_in[16]
port 96 nsew signal input
rlabel metal3 s 19600 17808 20000 17864 6 chany_top_in[17]
port 97 nsew signal input
rlabel metal2 s 9408 19600 9464 20000 6 chany_top_in[18]
port 98 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 chany_top_in[19]
port 99 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 chany_top_in[1]
port 100 nsew signal input
rlabel metal2 s 10080 19600 10136 20000 6 chany_top_in[2]
port 101 nsew signal input
rlabel metal2 s 336 0 392 400 6 chany_top_in[3]
port 102 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 chany_top_in[4]
port 103 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 chany_top_in[5]
port 104 nsew signal input
rlabel metal2 s 11424 19600 11480 20000 6 chany_top_in[6]
port 105 nsew signal input
rlabel metal2 s 17808 19600 17864 20000 6 chany_top_in[7]
port 106 nsew signal input
rlabel metal3 s 19600 14448 20000 14504 6 chany_top_in[8]
port 107 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 chany_top_in[9]
port 108 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 chany_top_out[0]
port 109 nsew signal output
rlabel metal2 s 17472 0 17528 400 6 chany_top_out[10]
port 110 nsew signal output
rlabel metal2 s 13776 19600 13832 20000 6 chany_top_out[11]
port 111 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 chany_top_out[12]
port 112 nsew signal output
rlabel metal2 s 13440 19600 13496 20000 6 chany_top_out[13]
port 113 nsew signal output
rlabel metal3 s 19600 4032 20000 4088 6 chany_top_out[14]
port 114 nsew signal output
rlabel metal2 s 16128 19600 16184 20000 6 chany_top_out[15]
port 115 nsew signal output
rlabel metal3 s 19600 15792 20000 15848 6 chany_top_out[16]
port 116 nsew signal output
rlabel metal2 s 12768 19600 12824 20000 6 chany_top_out[17]
port 117 nsew signal output
rlabel metal2 s 9744 19600 9800 20000 6 chany_top_out[18]
port 118 nsew signal output
rlabel metal3 s 19600 5040 20000 5096 6 chany_top_out[19]
port 119 nsew signal output
rlabel metal3 s 19600 18144 20000 18200 6 chany_top_out[1]
port 120 nsew signal output
rlabel metal3 s 19600 17472 20000 17528 6 chany_top_out[2]
port 121 nsew signal output
rlabel metal3 s 19600 19488 20000 19544 6 chany_top_out[3]
port 122 nsew signal output
rlabel metal3 s 19600 15120 20000 15176 6 chany_top_out[4]
port 123 nsew signal output
rlabel metal3 s 19600 2352 20000 2408 6 chany_top_out[5]
port 124 nsew signal output
rlabel metal3 s 19600 3024 20000 3080 6 chany_top_out[6]
port 125 nsew signal output
rlabel metal3 s 19600 3696 20000 3752 6 chany_top_out[7]
port 126 nsew signal output
rlabel metal3 s 19600 15456 20000 15512 6 chany_top_out[8]
port 127 nsew signal output
rlabel metal2 s 11088 0 11144 400 6 chany_top_out[9]
port 128 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 129 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 130 nsew signal input
rlabel metal2 s 0 0 56 400 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 131 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 132 nsew signal input
rlabel metal3 s 19600 8064 20000 8120 6 pReset
port 133 nsew signal input
rlabel metal3 s 0 13104 400 13160 6 prog_clk
port 134 nsew signal input
rlabel metal3 s 19600 7392 20000 7448 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 135 nsew signal input
rlabel metal3 s 19600 7728 20000 7784 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 136 nsew signal input
rlabel metal3 s 19600 6384 20000 6440 6 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 137 nsew signal input
rlabel metal3 s 19600 6048 20000 6104 6 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 138 nsew signal input
rlabel metal3 s 19600 6720 20000 6776 6 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 139 nsew signal input
rlabel metal3 s 19600 7056 20000 7112 6 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 140 nsew signal input
rlabel metal4 s 2923 1538 3083 18454 6 vdd
port 141 nsew power bidirectional
rlabel metal4 s 7585 1538 7745 18454 6 vdd
port 141 nsew power bidirectional
rlabel metal4 s 12247 1538 12407 18454 6 vdd
port 141 nsew power bidirectional
rlabel metal4 s 16909 1538 17069 18454 6 vdd
port 141 nsew power bidirectional
rlabel metal4 s 5254 1538 5414 18454 6 vss
port 142 nsew ground bidirectional
rlabel metal4 s 9916 1538 10076 18454 6 vss
port 142 nsew ground bidirectional
rlabel metal4 s 14578 1538 14738 18454 6 vss
port 142 nsew ground bidirectional
rlabel metal4 s 19240 1538 19400 18454 6 vss
port 142 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 834138
string GDS_FILE /home/baungarten/Desktop/2x2_FPGA_180nmD/openlane/sb_2__1_/runs/23_12_09_13_19/results/signoff/sb_2__1_.magic.gds
string GDS_START 99688
<< end >>

