// This is the unpowered netlist.
module grid_io_bottom (ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    top_width_0_height_0_subtile_0__pin_inpad_0_,
    top_width_0_height_0_subtile_0__pin_outpad_0_,
    top_width_0_height_0_subtile_1__pin_inpad_0_,
    top_width_0_height_0_subtile_1__pin_outpad_0_,
    top_width_0_height_0_subtile_2__pin_inpad_0_,
    top_width_0_height_0_subtile_2__pin_outpad_0_,
    top_width_0_height_0_subtile_3__pin_inpad_0_,
    top_width_0_height_0_subtile_3__pin_outpad_0_,
    gfpga_pad_GPIO_PAD);
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 output top_width_0_height_0_subtile_0__pin_inpad_0_;
 input top_width_0_height_0_subtile_0__pin_outpad_0_;
 output top_width_0_height_0_subtile_1__pin_inpad_0_;
 input top_width_0_height_0_subtile_1__pin_outpad_0_;
 output top_width_0_height_0_subtile_2__pin_inpad_0_;
 input top_width_0_height_0_subtile_2__pin_outpad_0_;
 output top_width_0_height_0_subtile_3__pin_inpad_0_;
 input top_width_0_height_0_subtile_3__pin_outpad_0_;
 inout [3:0] gfpga_pad_GPIO_PAD;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire clknet_0_prog_clk;
 wire clknet_1_0__leaf_prog_clk;
 wire clknet_1_1__leaf_prog_clk;
 wire \logical_tile_io_mode_io__0.ccff_tail ;
 wire \logical_tile_io_mode_io__1.ccff_tail ;
 wire \logical_tile_io_mode_io__2.ccff_tail ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(top_width_0_height_0_subtile_0__pin_outpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(top_width_0_height_0_subtile_1__pin_outpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(top_width_0_height_0_subtile_2__pin_outpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(top_width_0_height_0_subtile_3__pin_outpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_39 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _04_ (.I(net2),
    .ZN(_00_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05_ (.I(net2),
    .ZN(_01_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06_ (.I(net2),
    .ZN(_02_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07_ (.I(net2),
    .ZN(_03_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _08_ (.D(net1),
    .RN(_00_),
    .CLK(clknet_1_0__leaf_prog_clk),
    .Q(\logical_tile_io_mode_io__0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _09_ (.D(net13),
    .RN(_01_),
    .CLK(clknet_1_0__leaf_prog_clk),
    .Q(\logical_tile_io_mode_io__1.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _10_ (.D(net12),
    .RN(_02_),
    .CLK(clknet_1_1__leaf_prog_clk),
    .Q(\logical_tile_io_mode_io__2.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _11_ (.D(net14),
    .RN(_03_),
    .CLK(clknet_1_1__leaf_prog_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _12_ (.I(net6),
    .Z(gfpga_pad_GPIO_PAD[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _13_ (.I(net5),
    .Z(gfpga_pad_GPIO_PAD[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _14_ (.I(net4),
    .Z(gfpga_pad_GPIO_PAD[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _15_ (.I(net3),
    .Z(gfpga_pad_GPIO_PAD[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16_ (.I(net3),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _17_ (.I(net4),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _18_ (.I(net5),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _19_ (.I(net6),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\logical_tile_io_mode_io__1.ccff_tail ),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\logical_tile_io_mode_io__0.ccff_tail ),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\logical_tile_io_mode_io__2.ccff_tail ),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(pReset),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(top_width_0_height_0_subtile_0__pin_outpad_0_),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(top_width_0_height_0_subtile_1__pin_outpad_0_),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(top_width_0_height_0_subtile_2__pin_outpad_0_),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(top_width_0_height_0_subtile_3__pin_outpad_0_),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output10 (.I(net10),
    .Z(top_width_0_height_0_subtile_2__pin_inpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output11 (.I(net11),
    .Z(top_width_0_height_0_subtile_3__pin_inpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(top_width_0_height_0_subtile_0__pin_inpad_0_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output9 (.I(net9),
    .Z(top_width_0_height_0_subtile_1__pin_inpad_0_));
endmodule

