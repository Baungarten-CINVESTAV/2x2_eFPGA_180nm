magic
tech gf180mcuD
magscale 1 10
timestamp 1702148757
<< metal1 >>
rect 8530 26798 8542 26850
rect 8594 26847 8606 26850
rect 9426 26847 9438 26850
rect 8594 26801 9438 26847
rect 8594 26798 8606 26801
rect 9426 26798 9438 26801
rect 9490 26798 9502 26850
rect 10098 26798 10110 26850
rect 10162 26847 10174 26850
rect 11106 26847 11118 26850
rect 10162 26801 11118 26847
rect 10162 26798 10174 26801
rect 11106 26798 11118 26801
rect 11170 26798 11182 26850
rect 16818 26798 16830 26850
rect 16882 26847 16894 26850
rect 18274 26847 18286 26850
rect 16882 26801 18286 26847
rect 16882 26798 16894 26801
rect 18274 26798 18286 26801
rect 18338 26798 18350 26850
rect 22194 26798 22206 26850
rect 22258 26847 22270 26850
rect 23202 26847 23214 26850
rect 22258 26801 23214 26847
rect 22258 26798 22270 26801
rect 23202 26798 23214 26801
rect 23266 26798 23278 26850
rect 23538 26798 23550 26850
rect 23602 26847 23614 26850
rect 24994 26847 25006 26850
rect 23602 26801 25006 26847
rect 23602 26798 23614 26801
rect 24994 26798 25006 26801
rect 25058 26798 25070 26850
rect 1344 26682 28720 26716
rect 1344 26630 8018 26682
rect 8070 26630 8122 26682
rect 8174 26630 8226 26682
rect 8278 26630 14822 26682
rect 14874 26630 14926 26682
rect 14978 26630 15030 26682
rect 15082 26630 21626 26682
rect 21678 26630 21730 26682
rect 21782 26630 21834 26682
rect 21886 26630 28430 26682
rect 28482 26630 28534 26682
rect 28586 26630 28638 26682
rect 28690 26630 28720 26682
rect 1344 26596 28720 26630
rect 3726 26514 3778 26526
rect 3726 26450 3778 26462
rect 9438 26514 9490 26526
rect 9438 26450 9490 26462
rect 15822 26514 15874 26526
rect 15822 26450 15874 26462
rect 18286 26514 18338 26526
rect 18286 26450 18338 26462
rect 20302 26514 20354 26526
rect 20302 26450 20354 26462
rect 23214 26514 23266 26526
rect 23214 26450 23266 26462
rect 6078 26402 6130 26414
rect 6078 26338 6130 26350
rect 6750 26402 6802 26414
rect 6750 26338 6802 26350
rect 7422 26402 7474 26414
rect 7422 26338 7474 26350
rect 8094 26402 8146 26414
rect 8094 26338 8146 26350
rect 8766 26402 8818 26414
rect 20750 26402 20802 26414
rect 10658 26350 10670 26402
rect 10722 26350 10734 26402
rect 12226 26350 12238 26402
rect 12290 26350 12302 26402
rect 8766 26338 8818 26350
rect 20750 26338 20802 26350
rect 21422 26402 21474 26414
rect 21422 26338 21474 26350
rect 6414 26290 6466 26302
rect 13134 26290 13186 26302
rect 2930 26238 2942 26290
rect 2994 26238 3006 26290
rect 4386 26238 4398 26290
rect 4450 26238 4462 26290
rect 5842 26238 5854 26290
rect 5906 26238 5918 26290
rect 7186 26238 7198 26290
rect 7250 26238 7262 26290
rect 7858 26238 7870 26290
rect 7922 26238 7934 26290
rect 8530 26238 8542 26290
rect 8594 26238 8606 26290
rect 9762 26238 9774 26290
rect 9826 26238 9838 26290
rect 11330 26238 11342 26290
rect 11394 26238 11406 26290
rect 6414 26226 6466 26238
rect 13134 26226 13186 26238
rect 15038 26290 15090 26302
rect 18622 26290 18674 26302
rect 22430 26290 22482 26302
rect 17602 26238 17614 26290
rect 17666 26238 17678 26290
rect 20962 26238 20974 26290
rect 21026 26238 21038 26290
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 15038 26226 15090 26238
rect 18622 26226 18674 26238
rect 22430 26226 22482 26238
rect 24558 26290 24610 26302
rect 26562 26238 26574 26290
rect 26626 26238 26638 26290
rect 24558 26226 24610 26238
rect 3390 26178 3442 26190
rect 1922 26126 1934 26178
rect 1986 26126 1998 26178
rect 13570 26126 13582 26178
rect 13634 26126 13646 26178
rect 19058 26126 19070 26178
rect 19122 26126 19134 26178
rect 24994 26126 25006 26178
rect 25058 26126 25070 26178
rect 27682 26126 27694 26178
rect 27746 26126 27758 26178
rect 3390 26114 3442 26126
rect 1344 25898 28560 25932
rect 1344 25846 4616 25898
rect 4668 25846 4720 25898
rect 4772 25846 4824 25898
rect 4876 25846 11420 25898
rect 11472 25846 11524 25898
rect 11576 25846 11628 25898
rect 11680 25846 18224 25898
rect 18276 25846 18328 25898
rect 18380 25846 18432 25898
rect 18484 25846 25028 25898
rect 25080 25846 25132 25898
rect 25184 25846 25236 25898
rect 25288 25846 28560 25898
rect 1344 25812 28560 25846
rect 15026 25678 15038 25730
rect 15090 25727 15102 25730
rect 15362 25727 15374 25730
rect 15090 25681 15374 25727
rect 15090 25678 15102 25681
rect 15362 25678 15374 25681
rect 15426 25678 15438 25730
rect 1822 25618 1874 25630
rect 1822 25554 1874 25566
rect 5182 25618 5234 25630
rect 5182 25554 5234 25566
rect 6414 25618 6466 25630
rect 6414 25554 6466 25566
rect 6974 25618 7026 25630
rect 6974 25554 7026 25566
rect 7646 25618 7698 25630
rect 7646 25554 7698 25566
rect 8318 25618 8370 25630
rect 15038 25618 15090 25630
rect 11106 25566 11118 25618
rect 11170 25566 11182 25618
rect 12114 25566 12126 25618
rect 12178 25566 12190 25618
rect 8318 25554 8370 25566
rect 15038 25554 15090 25566
rect 15486 25618 15538 25630
rect 15486 25554 15538 25566
rect 17502 25618 17554 25630
rect 17502 25554 17554 25566
rect 18846 25618 18898 25630
rect 18846 25554 18898 25566
rect 20414 25618 20466 25630
rect 20414 25554 20466 25566
rect 20862 25618 20914 25630
rect 23538 25566 23550 25618
rect 23602 25566 23614 25618
rect 25330 25566 25342 25618
rect 25394 25566 25406 25618
rect 20862 25554 20914 25566
rect 3278 25506 3330 25518
rect 3278 25442 3330 25454
rect 3950 25506 4002 25518
rect 3950 25442 4002 25454
rect 5630 25506 5682 25518
rect 16382 25506 16434 25518
rect 15922 25454 15934 25506
rect 15986 25454 15998 25506
rect 5630 25442 5682 25454
rect 16382 25442 16434 25454
rect 17726 25506 17778 25518
rect 17726 25442 17778 25454
rect 19070 25506 19122 25518
rect 19070 25442 19122 25454
rect 21646 25506 21698 25518
rect 21646 25442 21698 25454
rect 5966 25394 6018 25406
rect 5966 25330 6018 25342
rect 13694 25394 13746 25406
rect 13694 25330 13746 25342
rect 14366 25394 14418 25406
rect 14366 25330 14418 25342
rect 21982 25394 22034 25406
rect 21982 25330 22034 25342
rect 23102 25394 23154 25406
rect 23102 25330 23154 25342
rect 26238 25394 26290 25406
rect 26238 25330 26290 25342
rect 2158 25282 2210 25294
rect 2158 25218 2210 25230
rect 2942 25282 2994 25294
rect 2942 25218 2994 25230
rect 3614 25282 3666 25294
rect 3614 25218 3666 25230
rect 4286 25282 4338 25294
rect 4286 25218 4338 25230
rect 10558 25282 10610 25294
rect 10558 25218 10610 25230
rect 11678 25282 11730 25294
rect 11678 25218 11730 25230
rect 15710 25282 15762 25294
rect 15710 25218 15762 25230
rect 16718 25282 16770 25294
rect 16718 25218 16770 25230
rect 18062 25282 18114 25294
rect 18062 25218 18114 25230
rect 19406 25282 19458 25294
rect 19406 25218 19458 25230
rect 21310 25282 21362 25294
rect 21310 25218 21362 25230
rect 24670 25282 24722 25294
rect 24670 25218 24722 25230
rect 26574 25282 26626 25294
rect 26574 25218 26626 25230
rect 26910 25282 26962 25294
rect 26910 25218 26962 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 28254 25282 28306 25294
rect 28254 25218 28306 25230
rect 1344 25114 28720 25148
rect 1344 25062 8018 25114
rect 8070 25062 8122 25114
rect 8174 25062 8226 25114
rect 8278 25062 14822 25114
rect 14874 25062 14926 25114
rect 14978 25062 15030 25114
rect 15082 25062 21626 25114
rect 21678 25062 21730 25114
rect 21782 25062 21834 25114
rect 21886 25062 28430 25114
rect 28482 25062 28534 25114
rect 28586 25062 28638 25114
rect 28690 25062 28720 25114
rect 1344 25028 28720 25062
rect 2158 24946 2210 24958
rect 2158 24882 2210 24894
rect 3614 24946 3666 24958
rect 3614 24882 3666 24894
rect 4622 24946 4674 24958
rect 4622 24882 4674 24894
rect 10110 24946 10162 24958
rect 10110 24882 10162 24894
rect 21198 24946 21250 24958
rect 21198 24882 21250 24894
rect 24110 24946 24162 24958
rect 24110 24882 24162 24894
rect 26126 24946 26178 24958
rect 26126 24882 26178 24894
rect 28142 24946 28194 24958
rect 28142 24882 28194 24894
rect 2942 24834 2994 24846
rect 2942 24770 2994 24782
rect 4958 24834 5010 24846
rect 4958 24770 5010 24782
rect 24670 24834 24722 24846
rect 24670 24770 24722 24782
rect 4286 24722 4338 24734
rect 10894 24722 10946 24734
rect 25342 24722 25394 24734
rect 3826 24670 3838 24722
rect 3890 24670 3902 24722
rect 5170 24670 5182 24722
rect 5234 24670 5246 24722
rect 20962 24670 20974 24722
rect 21026 24670 21038 24722
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 4286 24658 4338 24670
rect 10894 24658 10946 24670
rect 25342 24658 25394 24670
rect 26910 24722 26962 24734
rect 26910 24658 26962 24670
rect 27694 24722 27746 24734
rect 27694 24658 27746 24670
rect 1822 24610 1874 24622
rect 1822 24546 1874 24558
rect 1344 24330 28560 24364
rect 1344 24278 4616 24330
rect 4668 24278 4720 24330
rect 4772 24278 4824 24330
rect 4876 24278 11420 24330
rect 11472 24278 11524 24330
rect 11576 24278 11628 24330
rect 11680 24278 18224 24330
rect 18276 24278 18328 24330
rect 18380 24278 18432 24330
rect 18484 24278 25028 24330
rect 25080 24278 25132 24330
rect 25184 24278 25236 24330
rect 25288 24278 28560 24330
rect 1344 24244 28560 24278
rect 3166 24050 3218 24062
rect 27570 23998 27582 24050
rect 27634 23998 27646 24050
rect 3166 23986 3218 23998
rect 2382 23938 2434 23950
rect 9326 23938 9378 23950
rect 10670 23938 10722 23950
rect 4162 23886 4174 23938
rect 4226 23886 4238 23938
rect 4946 23886 4958 23938
rect 5010 23886 5022 23938
rect 10098 23886 10110 23938
rect 10162 23886 10174 23938
rect 2382 23874 2434 23886
rect 9326 23874 9378 23886
rect 10670 23874 10722 23886
rect 11342 23938 11394 23950
rect 17166 23938 17218 23950
rect 12114 23886 12126 23938
rect 12178 23886 12190 23938
rect 17938 23886 17950 23938
rect 18002 23886 18014 23938
rect 20514 23886 20526 23938
rect 20578 23886 20590 23938
rect 21410 23886 21422 23938
rect 21474 23886 21486 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 11342 23874 11394 23886
rect 17166 23874 17218 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 2046 23762 2098 23774
rect 2718 23826 2770 23838
rect 2718 23762 2770 23774
rect 3950 23826 4002 23838
rect 3950 23762 4002 23774
rect 6078 23826 6130 23838
rect 6078 23762 6130 23774
rect 9662 23826 9714 23838
rect 9662 23762 9714 23774
rect 10334 23826 10386 23838
rect 10334 23762 10386 23774
rect 11006 23826 11058 23838
rect 11006 23762 11058 23774
rect 11678 23826 11730 23838
rect 11678 23762 11730 23774
rect 12350 23826 12402 23838
rect 12350 23762 12402 23774
rect 17502 23826 17554 23838
rect 17502 23762 17554 23774
rect 18174 23826 18226 23838
rect 18174 23762 18226 23774
rect 20750 23826 20802 23838
rect 20750 23762 20802 23774
rect 21646 23826 21698 23838
rect 21646 23762 21698 23774
rect 24334 23826 24386 23838
rect 24334 23762 24386 23774
rect 24782 23826 24834 23838
rect 24782 23762 24834 23774
rect 25454 23826 25506 23838
rect 25454 23762 25506 23774
rect 25790 23826 25842 23838
rect 25790 23762 25842 23774
rect 26126 23826 26178 23838
rect 26126 23762 26178 23774
rect 4734 23714 4786 23726
rect 4734 23650 4786 23662
rect 5742 23714 5794 23726
rect 5742 23650 5794 23662
rect 25118 23714 25170 23726
rect 25118 23650 25170 23662
rect 26462 23714 26514 23726
rect 26462 23650 26514 23662
rect 26910 23714 26962 23726
rect 26910 23650 26962 23662
rect 28254 23714 28306 23726
rect 28254 23650 28306 23662
rect 1344 23546 28720 23580
rect 1344 23494 8018 23546
rect 8070 23494 8122 23546
rect 8174 23494 8226 23546
rect 8278 23494 14822 23546
rect 14874 23494 14926 23546
rect 14978 23494 15030 23546
rect 15082 23494 21626 23546
rect 21678 23494 21730 23546
rect 21782 23494 21834 23546
rect 21886 23494 28430 23546
rect 28482 23494 28534 23546
rect 28586 23494 28638 23546
rect 28690 23494 28720 23546
rect 1344 23460 28720 23494
rect 2046 23378 2098 23390
rect 2046 23314 2098 23326
rect 10558 23378 10610 23390
rect 10558 23314 10610 23326
rect 11230 23378 11282 23390
rect 11230 23314 11282 23326
rect 20974 23378 21026 23390
rect 20974 23314 21026 23326
rect 26462 23378 26514 23390
rect 26462 23314 26514 23326
rect 27134 23378 27186 23390
rect 27134 23314 27186 23326
rect 20638 23266 20690 23278
rect 20638 23202 20690 23214
rect 25790 23266 25842 23278
rect 25790 23202 25842 23214
rect 26126 23266 26178 23278
rect 26126 23202 26178 23214
rect 27470 23266 27522 23278
rect 27470 23202 27522 23214
rect 27806 23266 27858 23278
rect 27806 23202 27858 23214
rect 28142 23266 28194 23278
rect 28142 23202 28194 23214
rect 1710 23154 1762 23166
rect 10770 23102 10782 23154
rect 10834 23102 10846 23154
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 25554 23102 25566 23154
rect 25618 23102 25630 23154
rect 1710 23090 1762 23102
rect 2494 23042 2546 23054
rect 2494 22978 2546 22990
rect 1344 22762 28560 22796
rect 1344 22710 4616 22762
rect 4668 22710 4720 22762
rect 4772 22710 4824 22762
rect 4876 22710 11420 22762
rect 11472 22710 11524 22762
rect 11576 22710 11628 22762
rect 11680 22710 18224 22762
rect 18276 22710 18328 22762
rect 18380 22710 18432 22762
rect 18484 22710 25028 22762
rect 25080 22710 25132 22762
rect 25184 22710 25236 22762
rect 25288 22710 28560 22762
rect 1344 22676 28560 22710
rect 2942 22370 2994 22382
rect 28018 22318 28030 22370
rect 28082 22318 28094 22370
rect 2942 22306 2994 22318
rect 26462 22258 26514 22270
rect 26462 22194 26514 22206
rect 26798 22258 26850 22270
rect 26798 22194 26850 22206
rect 27134 22258 27186 22270
rect 27134 22194 27186 22206
rect 27470 22258 27522 22270
rect 27470 22194 27522 22206
rect 27806 22258 27858 22270
rect 27806 22194 27858 22206
rect 2158 22146 2210 22158
rect 2158 22082 2210 22094
rect 1344 21978 28720 22012
rect 1344 21926 8018 21978
rect 8070 21926 8122 21978
rect 8174 21926 8226 21978
rect 8278 21926 14822 21978
rect 14874 21926 14926 21978
rect 14978 21926 15030 21978
rect 15082 21926 21626 21978
rect 21678 21926 21730 21978
rect 21782 21926 21834 21978
rect 21886 21926 28430 21978
rect 28482 21926 28534 21978
rect 28586 21926 28638 21978
rect 28690 21926 28720 21978
rect 1344 21892 28720 21926
rect 2942 21810 2994 21822
rect 2942 21746 2994 21758
rect 27470 21810 27522 21822
rect 27470 21746 27522 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 22194 21646 22206 21698
rect 22258 21646 22270 21698
rect 28142 21586 28194 21598
rect 28142 21522 28194 21534
rect 27134 21474 27186 21486
rect 2258 21422 2270 21474
rect 2322 21422 2334 21474
rect 21186 21422 21198 21474
rect 21250 21422 21262 21474
rect 27134 21410 27186 21422
rect 1344 21194 28560 21228
rect 1344 21142 4616 21194
rect 4668 21142 4720 21194
rect 4772 21142 4824 21194
rect 4876 21142 11420 21194
rect 11472 21142 11524 21194
rect 11576 21142 11628 21194
rect 11680 21142 18224 21194
rect 18276 21142 18328 21194
rect 18380 21142 18432 21194
rect 18484 21142 25028 21194
rect 25080 21142 25132 21194
rect 25184 21142 25236 21194
rect 25288 21142 28560 21194
rect 1344 21108 28560 21142
rect 14466 20862 14478 20914
rect 14530 20862 14542 20914
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 2046 20690 2098 20702
rect 2046 20626 2098 20638
rect 2382 20690 2434 20702
rect 15474 20638 15486 20690
rect 15538 20638 15550 20690
rect 28018 20638 28030 20690
rect 28082 20638 28094 20690
rect 2382 20626 2434 20638
rect 19294 20578 19346 20590
rect 19294 20514 19346 20526
rect 1344 20410 28720 20444
rect 1344 20358 8018 20410
rect 8070 20358 8122 20410
rect 8174 20358 8226 20410
rect 8278 20358 14822 20410
rect 14874 20358 14926 20410
rect 14978 20358 15030 20410
rect 15082 20358 21626 20410
rect 21678 20358 21730 20410
rect 21782 20358 21834 20410
rect 21886 20358 28430 20410
rect 28482 20358 28534 20410
rect 28586 20358 28638 20410
rect 28690 20358 28720 20410
rect 1344 20324 28720 20358
rect 1822 20242 1874 20254
rect 1822 20178 1874 20190
rect 14366 20130 14418 20142
rect 19394 20078 19406 20130
rect 19458 20078 19470 20130
rect 22194 20078 22206 20130
rect 22258 20078 22270 20130
rect 14366 20066 14418 20078
rect 11454 20018 11506 20030
rect 12114 19966 12126 20018
rect 12178 19966 12190 20018
rect 16146 19966 16158 20018
rect 16210 19966 16222 20018
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 11454 19954 11506 19966
rect 18386 19854 18398 19906
rect 18450 19854 18462 19906
rect 21186 19854 21198 19906
rect 21250 19854 21262 19906
rect 28018 19854 28030 19906
rect 28082 19854 28094 19906
rect 15150 19794 15202 19806
rect 15150 19730 15202 19742
rect 16046 19794 16098 19806
rect 16046 19730 16098 19742
rect 1344 19626 28560 19660
rect 1344 19574 4616 19626
rect 4668 19574 4720 19626
rect 4772 19574 4824 19626
rect 4876 19574 11420 19626
rect 11472 19574 11524 19626
rect 11576 19574 11628 19626
rect 11680 19574 18224 19626
rect 18276 19574 18328 19626
rect 18380 19574 18432 19626
rect 18484 19574 25028 19626
rect 25080 19574 25132 19626
rect 25184 19574 25236 19626
rect 25288 19574 28560 19626
rect 1344 19540 28560 19574
rect 20638 19458 20690 19470
rect 20638 19394 20690 19406
rect 8642 19294 8654 19346
rect 8706 19294 8718 19346
rect 11442 19294 11454 19346
rect 11506 19294 11518 19346
rect 15250 19294 15262 19346
rect 15314 19294 15326 19346
rect 17166 19234 17218 19246
rect 23214 19234 23266 19246
rect 17602 19182 17614 19234
rect 17666 19182 17678 19234
rect 23874 19182 23886 19234
rect 23938 19182 23950 19234
rect 17166 19170 17218 19182
rect 23214 19170 23266 19182
rect 19854 19122 19906 19134
rect 9650 19070 9662 19122
rect 9714 19070 9726 19122
rect 12450 19070 12462 19122
rect 12514 19070 12526 19122
rect 16258 19070 16270 19122
rect 16322 19070 16334 19122
rect 19854 19058 19906 19070
rect 27470 19122 27522 19134
rect 27470 19058 27522 19070
rect 27806 19122 27858 19134
rect 27806 19058 27858 19070
rect 28142 19122 28194 19134
rect 28142 19058 28194 19070
rect 26910 19010 26962 19022
rect 26114 18958 26126 19010
rect 26178 18958 26190 19010
rect 26910 18946 26962 18958
rect 27134 19010 27186 19022
rect 27134 18946 27186 18958
rect 1344 18842 28720 18876
rect 1344 18790 8018 18842
rect 8070 18790 8122 18842
rect 8174 18790 8226 18842
rect 8278 18790 14822 18842
rect 14874 18790 14926 18842
rect 14978 18790 15030 18842
rect 15082 18790 21626 18842
rect 21678 18790 21730 18842
rect 21782 18790 21834 18842
rect 21886 18790 28430 18842
rect 28482 18790 28534 18842
rect 28586 18790 28638 18842
rect 28690 18790 28720 18842
rect 1344 18756 28720 18790
rect 8430 18674 8482 18686
rect 28254 18674 28306 18686
rect 12562 18622 12574 18674
rect 12626 18622 12638 18674
rect 16146 18622 16158 18674
rect 16210 18622 16222 18674
rect 8430 18610 8482 18622
rect 28254 18610 28306 18622
rect 7646 18562 7698 18574
rect 7646 18498 7698 18510
rect 21646 18562 21698 18574
rect 27234 18510 27246 18562
rect 27298 18510 27310 18562
rect 21646 18498 21698 18510
rect 4958 18450 5010 18462
rect 9438 18450 9490 18462
rect 13246 18450 13298 18462
rect 16942 18450 16994 18462
rect 18734 18450 18786 18462
rect 22430 18450 22482 18462
rect 5394 18398 5406 18450
rect 5458 18398 5470 18450
rect 10098 18398 10110 18450
rect 10162 18398 10174 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 18162 18398 18174 18450
rect 18226 18398 18238 18450
rect 19282 18398 19294 18450
rect 19346 18398 19358 18450
rect 23762 18398 23774 18450
rect 23826 18398 23838 18450
rect 4958 18386 5010 18398
rect 9438 18386 9490 18398
rect 13246 18386 13298 18398
rect 16942 18386 16994 18398
rect 18734 18386 18786 18398
rect 22430 18386 22482 18398
rect 13134 18338 13186 18350
rect 13134 18274 13186 18286
rect 23102 18338 23154 18350
rect 26226 18286 26238 18338
rect 26290 18286 26302 18338
rect 23102 18274 23154 18286
rect 18062 18226 18114 18238
rect 18062 18162 18114 18174
rect 23998 18226 24050 18238
rect 23998 18162 24050 18174
rect 1344 18058 28560 18092
rect 1344 18006 4616 18058
rect 4668 18006 4720 18058
rect 4772 18006 4824 18058
rect 4876 18006 11420 18058
rect 11472 18006 11524 18058
rect 11576 18006 11628 18058
rect 11680 18006 18224 18058
rect 18276 18006 18328 18058
rect 18380 18006 18432 18058
rect 18484 18006 25028 18058
rect 25080 18006 25132 18058
rect 25184 18006 25236 18058
rect 25288 18006 28560 18058
rect 1344 17972 28560 18006
rect 10782 17890 10834 17902
rect 6290 17838 6302 17890
rect 6354 17838 6366 17890
rect 10782 17826 10834 17838
rect 12574 17890 12626 17902
rect 12574 17826 12626 17838
rect 14142 17890 14194 17902
rect 14142 17826 14194 17838
rect 18958 17890 19010 17902
rect 18958 17826 19010 17838
rect 20066 17726 20078 17778
rect 20130 17726 20142 17778
rect 26114 17726 26126 17778
rect 26178 17726 26190 17778
rect 7086 17666 7138 17678
rect 15262 17666 15314 17678
rect 21198 17666 21250 17678
rect 4722 17614 4734 17666
rect 4786 17614 4798 17666
rect 6850 17614 6862 17666
rect 6914 17614 6926 17666
rect 7746 17614 7758 17666
rect 7810 17614 7822 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 14130 17614 14142 17666
rect 14194 17614 14206 17666
rect 15922 17614 15934 17666
rect 15986 17614 15998 17666
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 21858 17614 21870 17666
rect 21922 17614 21934 17666
rect 7086 17602 7138 17614
rect 15262 17602 15314 17614
rect 21198 17602 21250 17614
rect 18174 17554 18226 17566
rect 4834 17502 4846 17554
rect 4898 17502 4910 17554
rect 18174 17490 18226 17502
rect 24110 17554 24162 17566
rect 27122 17502 27134 17554
rect 27186 17502 27198 17554
rect 24110 17490 24162 17502
rect 24894 17442 24946 17454
rect 9986 17390 9998 17442
rect 10050 17390 10062 17442
rect 24894 17378 24946 17390
rect 1344 17274 28720 17308
rect 1344 17222 8018 17274
rect 8070 17222 8122 17274
rect 8174 17222 8226 17274
rect 8278 17222 14822 17274
rect 14874 17222 14926 17274
rect 14978 17222 15030 17274
rect 15082 17222 21626 17274
rect 21678 17222 21730 17274
rect 21782 17222 21834 17274
rect 21886 17222 28430 17274
rect 28482 17222 28534 17274
rect 28586 17222 28638 17274
rect 28690 17222 28720 17274
rect 1344 17188 28720 17222
rect 5842 17054 5854 17106
rect 5906 17054 5918 17106
rect 9762 16942 9774 16994
rect 9826 16942 9838 16994
rect 21410 16942 21422 16994
rect 21474 16942 21486 16994
rect 27234 16942 27246 16994
rect 27298 16942 27310 16994
rect 3166 16882 3218 16894
rect 3602 16830 3614 16882
rect 3666 16830 3678 16882
rect 7522 16830 7534 16882
rect 7586 16830 7598 16882
rect 14690 16830 14702 16882
rect 14754 16830 14766 16882
rect 19506 16830 19518 16882
rect 19570 16830 19582 16882
rect 3166 16818 3218 16830
rect 26226 16718 26238 16770
rect 26290 16718 26302 16770
rect 6638 16658 6690 16670
rect 6638 16594 6690 16606
rect 7310 16658 7362 16670
rect 7310 16594 7362 16606
rect 1344 16490 28560 16524
rect 1344 16438 4616 16490
rect 4668 16438 4720 16490
rect 4772 16438 4824 16490
rect 4876 16438 11420 16490
rect 11472 16438 11524 16490
rect 11576 16438 11628 16490
rect 11680 16438 18224 16490
rect 18276 16438 18328 16490
rect 18380 16438 18432 16490
rect 18484 16438 25028 16490
rect 25080 16438 25132 16490
rect 25184 16438 25236 16490
rect 25288 16438 28560 16490
rect 1344 16404 28560 16438
rect 3826 16158 3838 16210
rect 3890 16158 3902 16210
rect 6178 16158 6190 16210
rect 6242 16158 6254 16210
rect 9986 16158 9998 16210
rect 10050 16158 10062 16210
rect 26674 16158 26686 16210
rect 26738 16158 26750 16210
rect 19406 16098 19458 16110
rect 24670 16098 24722 16110
rect 12898 16046 12910 16098
rect 12962 16046 12974 16098
rect 13682 16046 13694 16098
rect 13746 16046 13758 16098
rect 19058 16046 19070 16098
rect 19122 16046 19134 16098
rect 19842 16046 19854 16098
rect 19906 16046 19918 16098
rect 24322 16046 24334 16098
rect 24386 16046 24398 16098
rect 19406 16034 19458 16046
rect 24670 16034 24722 16046
rect 2706 15934 2718 15986
rect 2770 15934 2782 15986
rect 7298 15934 7310 15986
rect 7362 15934 7374 15986
rect 11106 15934 11118 15986
rect 11170 15934 11182 15986
rect 27682 15934 27694 15986
rect 27746 15934 27758 15986
rect 13582 15874 13634 15886
rect 12338 15822 12350 15874
rect 12402 15822 12414 15874
rect 13582 15810 13634 15822
rect 15934 15874 15986 15886
rect 21198 15874 21250 15886
rect 25230 15874 25282 15886
rect 16706 15822 16718 15874
rect 16770 15822 16782 15874
rect 20402 15822 20414 15874
rect 20466 15822 20478 15874
rect 21970 15822 21982 15874
rect 22034 15822 22046 15874
rect 15934 15810 15986 15822
rect 21198 15810 21250 15822
rect 25230 15810 25282 15822
rect 1344 15706 28720 15740
rect 1344 15654 8018 15706
rect 8070 15654 8122 15706
rect 8174 15654 8226 15706
rect 8278 15654 14822 15706
rect 14874 15654 14926 15706
rect 14978 15654 15030 15706
rect 15082 15654 21626 15706
rect 21678 15654 21730 15706
rect 21782 15654 21834 15706
rect 21886 15654 28430 15706
rect 28482 15654 28534 15706
rect 28586 15654 28638 15706
rect 28690 15654 28720 15706
rect 1344 15620 28720 15654
rect 1934 15538 1986 15550
rect 1934 15474 1986 15486
rect 11118 15538 11170 15550
rect 16718 15538 16770 15550
rect 11890 15486 11902 15538
rect 11954 15486 11966 15538
rect 11118 15474 11170 15486
rect 16718 15474 16770 15486
rect 24558 15538 24610 15550
rect 24558 15474 24610 15486
rect 27694 15538 27746 15550
rect 27694 15474 27746 15486
rect 2718 15426 2770 15438
rect 7970 15374 7982 15426
rect 8034 15374 8046 15426
rect 9874 15374 9886 15426
rect 9938 15374 9950 15426
rect 17490 15374 17502 15426
rect 17554 15374 17566 15426
rect 22306 15374 22318 15426
rect 22370 15374 22382 15426
rect 2718 15362 2770 15374
rect 5406 15314 5458 15326
rect 14590 15314 14642 15326
rect 4946 15262 4958 15314
rect 5010 15262 5022 15314
rect 10210 15262 10222 15314
rect 10274 15262 10286 15314
rect 14130 15262 14142 15314
rect 14194 15262 14206 15314
rect 16482 15262 16494 15314
rect 16546 15262 16558 15314
rect 24322 15262 24334 15314
rect 24386 15262 24398 15314
rect 25666 15262 25678 15314
rect 25730 15262 25742 15314
rect 27010 15262 27022 15314
rect 27074 15262 27086 15314
rect 5406 15250 5458 15262
rect 14590 15250 14642 15262
rect 23550 15202 23602 15214
rect 6962 15150 6974 15202
rect 7026 15150 7038 15202
rect 18610 15150 18622 15202
rect 18674 15150 18686 15202
rect 21298 15150 21310 15202
rect 21362 15150 21374 15202
rect 25554 15150 25566 15202
rect 25618 15150 25630 15202
rect 23550 15138 23602 15150
rect 1344 14922 28560 14956
rect 1344 14870 4616 14922
rect 4668 14870 4720 14922
rect 4772 14870 4824 14922
rect 4876 14870 11420 14922
rect 11472 14870 11524 14922
rect 11576 14870 11628 14922
rect 11680 14870 18224 14922
rect 18276 14870 18328 14922
rect 18380 14870 18432 14922
rect 18484 14870 25028 14922
rect 25080 14870 25132 14922
rect 25184 14870 25236 14922
rect 25288 14870 28560 14922
rect 1344 14836 28560 14870
rect 3950 14754 4002 14766
rect 3950 14690 4002 14702
rect 26350 14754 26402 14766
rect 26350 14690 26402 14702
rect 14254 14642 14306 14654
rect 8082 14590 8094 14642
rect 8146 14590 8158 14642
rect 19506 14590 19518 14642
rect 19570 14590 19582 14642
rect 26898 14590 26910 14642
rect 26962 14590 26974 14642
rect 14254 14578 14306 14590
rect 9550 14530 9602 14542
rect 28142 14530 28194 14542
rect 4162 14478 4174 14530
rect 4226 14478 4238 14530
rect 9986 14478 9998 14530
rect 10050 14478 10062 14530
rect 14466 14478 14478 14530
rect 14530 14478 14542 14530
rect 22082 14478 22094 14530
rect 22146 14478 22158 14530
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 23314 14478 23326 14530
rect 23378 14478 23390 14530
rect 26562 14478 26574 14530
rect 26626 14478 26638 14530
rect 9550 14466 9602 14478
rect 28142 14466 28194 14478
rect 25566 14418 25618 14430
rect 6738 14366 6750 14418
rect 6802 14366 6814 14418
rect 25566 14354 25618 14366
rect 27806 14418 27858 14430
rect 27806 14354 27858 14366
rect 13022 14306 13074 14318
rect 12338 14254 12350 14306
rect 12402 14254 12414 14306
rect 13022 14242 13074 14254
rect 20750 14306 20802 14318
rect 20750 14242 20802 14254
rect 22318 14306 22370 14318
rect 22318 14242 22370 14254
rect 1344 14138 28720 14172
rect 1344 14086 8018 14138
rect 8070 14086 8122 14138
rect 8174 14086 8226 14138
rect 8278 14086 14822 14138
rect 14874 14086 14926 14138
rect 14978 14086 15030 14138
rect 15082 14086 21626 14138
rect 21678 14086 21730 14138
rect 21782 14086 21834 14138
rect 21886 14086 28430 14138
rect 28482 14086 28534 14138
rect 28586 14086 28638 14138
rect 28690 14086 28720 14138
rect 1344 14052 28720 14086
rect 5406 13970 5458 13982
rect 28254 13970 28306 13982
rect 6178 13918 6190 13970
rect 6242 13918 6254 13970
rect 20514 13918 20526 13970
rect 20578 13918 20590 13970
rect 5406 13906 5458 13918
rect 28254 13906 28306 13918
rect 2382 13858 2434 13870
rect 21310 13858 21362 13870
rect 11778 13806 11790 13858
rect 11842 13806 11854 13858
rect 13906 13806 13918 13858
rect 13970 13806 13982 13858
rect 22754 13806 22766 13858
rect 22818 13806 22830 13858
rect 2382 13794 2434 13806
rect 21310 13794 21362 13806
rect 17614 13746 17666 13758
rect 4722 13694 4734 13746
rect 4786 13694 4798 13746
rect 5170 13694 5182 13746
rect 5234 13694 5246 13746
rect 8418 13694 8430 13746
rect 8482 13694 8494 13746
rect 8978 13694 8990 13746
rect 9042 13694 9054 13746
rect 18274 13694 18286 13746
rect 18338 13694 18350 13746
rect 17614 13682 17666 13694
rect 25902 13634 25954 13646
rect 10770 13582 10782 13634
rect 10834 13582 10846 13634
rect 15026 13582 15038 13634
rect 15090 13582 15102 13634
rect 21970 13582 21982 13634
rect 22034 13582 22046 13634
rect 25902 13570 25954 13582
rect 26238 13634 26290 13646
rect 26238 13570 26290 13582
rect 1598 13522 1650 13534
rect 1598 13458 1650 13470
rect 1344 13354 28560 13388
rect 1344 13302 4616 13354
rect 4668 13302 4720 13354
rect 4772 13302 4824 13354
rect 4876 13302 11420 13354
rect 11472 13302 11524 13354
rect 11576 13302 11628 13354
rect 11680 13302 18224 13354
rect 18276 13302 18328 13354
rect 18380 13302 18432 13354
rect 18484 13302 25028 13354
rect 25080 13302 25132 13354
rect 25184 13302 25236 13354
rect 25288 13302 28560 13354
rect 1344 13268 28560 13302
rect 3278 13186 3330 13198
rect 3278 13122 3330 13134
rect 9214 13186 9266 13198
rect 9214 13122 9266 13134
rect 16382 13186 16434 13198
rect 16382 13122 16434 13134
rect 5518 12962 5570 12974
rect 12798 12962 12850 12974
rect 22206 12962 22258 12974
rect 3378 12910 3390 12962
rect 3442 12910 3454 12962
rect 4610 12910 4622 12962
rect 4674 12910 4686 12962
rect 6178 12910 6190 12962
rect 6242 12910 6254 12962
rect 12450 12910 12462 12962
rect 12514 12910 12526 12962
rect 18722 12910 18734 12962
rect 18786 12910 18798 12962
rect 22642 12910 22654 12962
rect 22706 12910 22718 12962
rect 25890 12910 25902 12962
rect 25954 12910 25966 12962
rect 5518 12898 5570 12910
rect 12798 12898 12850 12910
rect 22206 12898 22258 12910
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12738 2098 12750
rect 2046 12674 2098 12686
rect 2494 12738 2546 12750
rect 2494 12674 2546 12686
rect 4398 12738 4450 12750
rect 9326 12738 9378 12750
rect 21422 12738 21474 12750
rect 25678 12738 25730 12750
rect 8642 12686 8654 12738
rect 8706 12686 8718 12738
rect 10098 12686 10110 12738
rect 10162 12686 10174 12738
rect 25106 12686 25118 12738
rect 25170 12686 25182 12738
rect 4398 12674 4450 12686
rect 9326 12674 9378 12686
rect 21422 12674 21474 12686
rect 25678 12674 25730 12686
rect 26014 12738 26066 12750
rect 26014 12674 26066 12686
rect 1344 12570 28720 12604
rect 1344 12518 8018 12570
rect 8070 12518 8122 12570
rect 8174 12518 8226 12570
rect 8278 12518 14822 12570
rect 14874 12518 14926 12570
rect 14978 12518 15030 12570
rect 15082 12518 21626 12570
rect 21678 12518 21730 12570
rect 21782 12518 21834 12570
rect 21886 12518 28430 12570
rect 28482 12518 28534 12570
rect 28586 12518 28638 12570
rect 28690 12518 28720 12570
rect 1344 12484 28720 12518
rect 3502 12402 3554 12414
rect 4274 12350 4286 12402
rect 4338 12350 4350 12402
rect 3502 12338 3554 12350
rect 8642 12238 8654 12290
rect 8706 12238 8718 12290
rect 9762 12238 9774 12290
rect 9826 12238 9838 12290
rect 27234 12238 27246 12290
rect 27298 12238 27310 12290
rect 6974 12178 7026 12190
rect 2034 12126 2046 12178
rect 2098 12175 2110 12178
rect 2482 12175 2494 12178
rect 2098 12129 2494 12175
rect 2098 12126 2110 12129
rect 2482 12126 2494 12129
rect 2546 12126 2558 12178
rect 3266 12126 3278 12178
rect 3330 12126 3342 12178
rect 6626 12126 6638 12178
rect 6690 12126 6702 12178
rect 8530 12126 8542 12178
rect 8594 12126 8606 12178
rect 14802 12126 14814 12178
rect 14866 12126 14878 12178
rect 19506 12126 19518 12178
rect 19570 12126 19582 12178
rect 6974 12114 7026 12126
rect 18734 12066 18786 12078
rect 25566 12066 25618 12078
rect 19058 12014 19070 12066
rect 19122 12014 19134 12066
rect 24434 12014 24446 12066
rect 24498 12014 24510 12066
rect 26226 12014 26238 12066
rect 26290 12014 26302 12066
rect 18734 12002 18786 12014
rect 25566 12002 25618 12014
rect 3166 11954 3218 11966
rect 3166 11890 3218 11902
rect 1344 11786 28560 11820
rect 1344 11734 4616 11786
rect 4668 11734 4720 11786
rect 4772 11734 4824 11786
rect 4876 11734 11420 11786
rect 11472 11734 11524 11786
rect 11576 11734 11628 11786
rect 11680 11734 18224 11786
rect 18276 11734 18328 11786
rect 18380 11734 18432 11786
rect 18484 11734 25028 11786
rect 25080 11734 25132 11786
rect 25184 11734 25236 11786
rect 25288 11734 28560 11786
rect 1344 11700 28560 11734
rect 9102 11618 9154 11630
rect 9102 11554 9154 11566
rect 24894 11618 24946 11630
rect 24894 11554 24946 11566
rect 25230 11506 25282 11518
rect 3714 11454 3726 11506
rect 3778 11454 3790 11506
rect 16258 11454 16270 11506
rect 16322 11454 16334 11506
rect 19282 11454 19294 11506
rect 19346 11454 19358 11506
rect 26674 11454 26686 11506
rect 26738 11454 26750 11506
rect 25230 11442 25282 11454
rect 21422 11394 21474 11406
rect 5954 11342 5966 11394
rect 6018 11342 6030 11394
rect 12674 11342 12686 11394
rect 12738 11342 12750 11394
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 21422 11330 21474 11342
rect 24110 11282 24162 11294
rect 2594 11230 2606 11282
rect 2658 11230 2670 11282
rect 17266 11230 17278 11282
rect 17330 11230 17342 11282
rect 20290 11230 20302 11282
rect 20354 11230 20366 11282
rect 27682 11230 27694 11282
rect 27746 11230 27758 11282
rect 24110 11218 24162 11230
rect 5742 11170 5794 11182
rect 5742 11106 5794 11118
rect 1344 11002 28720 11036
rect 1344 10950 8018 11002
rect 8070 10950 8122 11002
rect 8174 10950 8226 11002
rect 8278 10950 14822 11002
rect 14874 10950 14926 11002
rect 14978 10950 15030 11002
rect 15082 10950 21626 11002
rect 21678 10950 21730 11002
rect 21782 10950 21834 11002
rect 21886 10950 28430 11002
rect 28482 10950 28534 11002
rect 28586 10950 28638 11002
rect 28690 10950 28720 11002
rect 1344 10916 28720 10950
rect 16270 10834 16322 10846
rect 25342 10834 25394 10846
rect 5506 10782 5518 10834
rect 5570 10782 5582 10834
rect 20178 10782 20190 10834
rect 20242 10782 20254 10834
rect 16270 10770 16322 10782
rect 25342 10770 25394 10782
rect 25790 10834 25842 10846
rect 25790 10770 25842 10782
rect 6078 10722 6130 10734
rect 15486 10722 15538 10734
rect 2034 10670 2046 10722
rect 2098 10670 2110 10722
rect 6402 10670 6414 10722
rect 6466 10670 6478 10722
rect 11778 10670 11790 10722
rect 11842 10670 11854 10722
rect 6078 10658 6130 10670
rect 15486 10658 15538 10670
rect 23998 10722 24050 10734
rect 27234 10670 27246 10722
rect 27298 10670 27310 10722
rect 23998 10658 24050 10670
rect 2382 10610 2434 10622
rect 12798 10610 12850 10622
rect 17278 10610 17330 10622
rect 21310 10610 21362 10622
rect 1810 10558 1822 10610
rect 1874 10558 1886 10610
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 13234 10558 13246 10610
rect 13298 10558 13310 10610
rect 17938 10558 17950 10610
rect 18002 10558 18014 10610
rect 21746 10558 21758 10610
rect 21810 10558 21822 10610
rect 2382 10546 2434 10558
rect 12798 10546 12850 10558
rect 17278 10546 17330 10558
rect 21310 10546 21362 10558
rect 16830 10498 16882 10510
rect 7522 10446 7534 10498
rect 7586 10446 7598 10498
rect 10770 10446 10782 10498
rect 10834 10446 10846 10498
rect 16482 10446 16494 10498
rect 16546 10446 16558 10498
rect 26226 10446 26238 10498
rect 26290 10446 26302 10498
rect 16830 10434 16882 10446
rect 20974 10386 21026 10398
rect 20974 10322 21026 10334
rect 24782 10386 24834 10398
rect 24782 10322 24834 10334
rect 1344 10218 28560 10252
rect 1344 10166 4616 10218
rect 4668 10166 4720 10218
rect 4772 10166 4824 10218
rect 4876 10166 11420 10218
rect 11472 10166 11524 10218
rect 11576 10166 11628 10218
rect 11680 10166 18224 10218
rect 18276 10166 18328 10218
rect 18380 10166 18432 10218
rect 18484 10166 25028 10218
rect 25080 10166 25132 10218
rect 25184 10166 25236 10218
rect 25288 10166 28560 10218
rect 1344 10132 28560 10166
rect 18958 10050 19010 10062
rect 18958 9986 19010 9998
rect 25566 10050 25618 10062
rect 25566 9986 25618 9998
rect 27694 10050 27746 10062
rect 27694 9986 27746 9998
rect 1822 9938 1874 9950
rect 19182 9938 19234 9950
rect 6626 9886 6638 9938
rect 6690 9886 6702 9938
rect 15026 9886 15038 9938
rect 15090 9886 15102 9938
rect 1822 9874 1874 9886
rect 19182 9874 19234 9886
rect 21422 9938 21474 9950
rect 21422 9874 21474 9886
rect 9550 9826 9602 9838
rect 14702 9826 14754 9838
rect 9986 9774 9998 9826
rect 10050 9774 10062 9826
rect 14130 9774 14142 9826
rect 14194 9774 14206 9826
rect 9550 9762 9602 9774
rect 14702 9762 14754 9774
rect 15486 9826 15538 9838
rect 19966 9826 20018 9838
rect 15922 9774 15934 9826
rect 15986 9774 15998 9826
rect 15486 9762 15538 9774
rect 19966 9762 20018 9774
rect 21870 9826 21922 9838
rect 26910 9826 26962 9838
rect 22530 9774 22542 9826
rect 22594 9774 22606 9826
rect 25778 9774 25790 9826
rect 25842 9774 25854 9826
rect 21870 9762 21922 9774
rect 26910 9762 26962 9774
rect 7634 9662 7646 9714
rect 7698 9662 7710 9714
rect 13906 9662 13918 9714
rect 13970 9662 13982 9714
rect 13022 9602 13074 9614
rect 19294 9602 19346 9614
rect 25902 9602 25954 9614
rect 12450 9550 12462 9602
rect 12514 9550 12526 9602
rect 18386 9550 18398 9602
rect 18450 9550 18462 9602
rect 24770 9550 24782 9602
rect 24834 9550 24846 9602
rect 13022 9538 13074 9550
rect 19294 9538 19346 9550
rect 25902 9538 25954 9550
rect 1344 9434 28720 9468
rect 1344 9382 8018 9434
rect 8070 9382 8122 9434
rect 8174 9382 8226 9434
rect 8278 9382 14822 9434
rect 14874 9382 14926 9434
rect 14978 9382 15030 9434
rect 15082 9382 21626 9434
rect 21678 9382 21730 9434
rect 21782 9382 21834 9434
rect 21886 9382 28430 9434
rect 28482 9382 28534 9434
rect 28586 9382 28638 9434
rect 28690 9382 28720 9434
rect 1344 9348 28720 9382
rect 5518 9266 5570 9278
rect 21646 9266 21698 9278
rect 4946 9214 4958 9266
rect 5010 9214 5022 9266
rect 16370 9214 16382 9266
rect 16434 9214 16446 9266
rect 5518 9202 5570 9214
rect 21646 9202 21698 9214
rect 23550 9266 23602 9278
rect 23550 9202 23602 9214
rect 24558 9266 24610 9278
rect 24558 9202 24610 9214
rect 25454 9266 25506 9278
rect 25454 9202 25506 9214
rect 12450 9102 12462 9154
rect 12514 9102 12526 9154
rect 27234 9102 27246 9154
rect 27298 9102 27310 9154
rect 2046 9042 2098 9054
rect 13246 9042 13298 9054
rect 2482 8990 2494 9042
rect 2546 8990 2558 9042
rect 9762 8990 9774 9042
rect 9826 8990 9838 9042
rect 12674 8990 12686 9042
rect 12738 8990 12750 9042
rect 13794 8990 13806 9042
rect 13858 8990 13870 9042
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 24322 8990 24334 9042
rect 24386 8990 24398 9042
rect 2046 8978 2098 8990
rect 13246 8978 13298 8990
rect 11902 8930 11954 8942
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 11902 8866 11954 8878
rect 16942 8818 16994 8830
rect 16942 8754 16994 8766
rect 1344 8650 28560 8684
rect 1344 8598 4616 8650
rect 4668 8598 4720 8650
rect 4772 8598 4824 8650
rect 4876 8598 11420 8650
rect 11472 8598 11524 8650
rect 11576 8598 11628 8650
rect 11680 8598 18224 8650
rect 18276 8598 18328 8650
rect 18380 8598 18432 8650
rect 18484 8598 25028 8650
rect 25080 8598 25132 8650
rect 25184 8598 25236 8650
rect 25288 8598 28560 8650
rect 1344 8564 28560 8598
rect 26574 8370 26626 8382
rect 14466 8318 14478 8370
rect 14530 8318 14542 8370
rect 17602 8318 17614 8370
rect 17666 8318 17678 8370
rect 27682 8318 27694 8370
rect 27746 8318 27758 8370
rect 26574 8306 26626 8318
rect 2930 8206 2942 8258
rect 2994 8206 3006 8258
rect 3378 8206 3390 8258
rect 3442 8206 3454 8258
rect 22978 8206 22990 8258
rect 23042 8206 23054 8258
rect 23538 8206 23550 8258
rect 23602 8206 23614 8258
rect 27010 8206 27022 8258
rect 27074 8206 27086 8258
rect 4062 8146 4114 8158
rect 2034 8094 2046 8146
rect 2098 8094 2110 8146
rect 15474 8094 15486 8146
rect 15538 8094 15550 8146
rect 18610 8094 18622 8146
rect 18674 8094 18686 8146
rect 4062 8082 4114 8094
rect 3614 8034 3666 8046
rect 25890 7982 25902 8034
rect 25954 7982 25966 8034
rect 3614 7970 3666 7982
rect 1344 7866 28720 7900
rect 1344 7814 8018 7866
rect 8070 7814 8122 7866
rect 8174 7814 8226 7866
rect 8278 7814 14822 7866
rect 14874 7814 14926 7866
rect 14978 7814 15030 7866
rect 15082 7814 21626 7866
rect 21678 7814 21730 7866
rect 21782 7814 21834 7866
rect 21886 7814 28430 7866
rect 28482 7814 28534 7866
rect 28586 7814 28638 7866
rect 28690 7814 28720 7866
rect 1344 7780 28720 7814
rect 23998 7698 24050 7710
rect 23998 7634 24050 7646
rect 22082 7534 22094 7586
rect 22146 7534 22158 7586
rect 25330 7534 25342 7586
rect 25394 7534 25406 7586
rect 2930 7422 2942 7474
rect 2994 7422 3006 7474
rect 23986 7422 23998 7474
rect 24050 7422 24062 7474
rect 23550 7362 23602 7374
rect 27134 7362 27186 7374
rect 1922 7310 1934 7362
rect 1986 7310 1998 7362
rect 20738 7310 20750 7362
rect 20802 7310 20814 7362
rect 26450 7310 26462 7362
rect 26514 7310 26526 7362
rect 23550 7298 23602 7310
rect 27134 7298 27186 7310
rect 27806 7362 27858 7374
rect 27806 7298 27858 7310
rect 27458 7198 27470 7250
rect 27522 7247 27534 7250
rect 27794 7247 27806 7250
rect 27522 7201 27806 7247
rect 27522 7198 27534 7201
rect 27794 7198 27806 7201
rect 27858 7198 27870 7250
rect 1344 7082 28560 7116
rect 1344 7030 4616 7082
rect 4668 7030 4720 7082
rect 4772 7030 4824 7082
rect 4876 7030 11420 7082
rect 11472 7030 11524 7082
rect 11576 7030 11628 7082
rect 11680 7030 18224 7082
rect 18276 7030 18328 7082
rect 18380 7030 18432 7082
rect 18484 7030 25028 7082
rect 25080 7030 25132 7082
rect 25184 7030 25236 7082
rect 25288 7030 28560 7082
rect 1344 6996 28560 7030
rect 23102 6914 23154 6926
rect 23102 6850 23154 6862
rect 22990 6690 23042 6702
rect 26798 6690 26850 6702
rect 3378 6638 3390 6690
rect 3442 6638 3454 6690
rect 4722 6638 4734 6690
rect 4786 6638 4798 6690
rect 26226 6638 26238 6690
rect 26290 6638 26302 6690
rect 22990 6626 23042 6638
rect 26798 6626 26850 6638
rect 28142 6690 28194 6702
rect 28142 6626 28194 6638
rect 1710 6578 1762 6590
rect 1710 6514 1762 6526
rect 2046 6578 2098 6590
rect 2046 6514 2098 6526
rect 3838 6578 3890 6590
rect 3838 6514 3890 6526
rect 4174 6578 4226 6590
rect 4174 6514 4226 6526
rect 27470 6578 27522 6590
rect 27470 6514 27522 6526
rect 27806 6578 27858 6590
rect 27806 6514 27858 6526
rect 2494 6466 2546 6478
rect 2494 6402 2546 6414
rect 3166 6466 3218 6478
rect 3166 6402 3218 6414
rect 4510 6466 4562 6478
rect 27134 6466 27186 6478
rect 23874 6414 23886 6466
rect 23938 6414 23950 6466
rect 4510 6402 4562 6414
rect 27134 6402 27186 6414
rect 1344 6298 28720 6332
rect 1344 6246 8018 6298
rect 8070 6246 8122 6298
rect 8174 6246 8226 6298
rect 8278 6246 14822 6298
rect 14874 6246 14926 6298
rect 14978 6246 15030 6298
rect 15082 6246 21626 6298
rect 21678 6246 21730 6298
rect 21782 6246 21834 6298
rect 21886 6246 28430 6298
rect 28482 6246 28534 6298
rect 28586 6246 28638 6298
rect 28690 6246 28720 6298
rect 1344 6212 28720 6246
rect 27694 6130 27746 6142
rect 25442 6078 25454 6130
rect 25506 6078 25518 6130
rect 27694 6066 27746 6078
rect 28254 6130 28306 6142
rect 28254 6066 28306 6078
rect 10334 6018 10386 6030
rect 10334 5954 10386 5966
rect 11118 6018 11170 6030
rect 11118 5954 11170 5966
rect 23998 6018 24050 6030
rect 23998 5954 24050 5966
rect 24670 6018 24722 6030
rect 24670 5954 24722 5966
rect 9998 5906 10050 5918
rect 24334 5906 24386 5918
rect 26910 5906 26962 5918
rect 2930 5854 2942 5906
rect 2994 5854 3006 5906
rect 10882 5854 10894 5906
rect 10946 5854 10958 5906
rect 25666 5854 25678 5906
rect 25730 5854 25742 5906
rect 9998 5842 10050 5854
rect 24334 5842 24386 5854
rect 26910 5842 26962 5854
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 1344 5514 28560 5548
rect 1344 5462 4616 5514
rect 4668 5462 4720 5514
rect 4772 5462 4824 5514
rect 4876 5462 11420 5514
rect 11472 5462 11524 5514
rect 11576 5462 11628 5514
rect 11680 5462 18224 5514
rect 18276 5462 18328 5514
rect 18380 5462 18432 5514
rect 18484 5462 25028 5514
rect 25080 5462 25132 5514
rect 25184 5462 25236 5514
rect 25288 5462 28560 5514
rect 1344 5428 28560 5462
rect 27570 5182 27582 5234
rect 27634 5182 27646 5234
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 2494 5122 2546 5134
rect 24334 5122 24386 5134
rect 9986 5070 9998 5122
rect 10050 5070 10062 5122
rect 2494 5058 2546 5070
rect 24334 5058 24386 5070
rect 24558 5122 24610 5134
rect 25902 5122 25954 5134
rect 25330 5070 25342 5122
rect 25394 5070 25406 5122
rect 24558 5058 24610 5070
rect 25902 5058 25954 5070
rect 26910 5122 26962 5134
rect 26910 5058 26962 5070
rect 2046 5010 2098 5022
rect 2046 4946 2098 4958
rect 20414 5010 20466 5022
rect 20414 4946 20466 4958
rect 10222 4898 10274 4910
rect 10222 4834 10274 4846
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 24894 4898 24946 4910
rect 24894 4834 24946 4846
rect 25566 4898 25618 4910
rect 25566 4834 25618 4846
rect 26238 4898 26290 4910
rect 26238 4834 26290 4846
rect 1344 4730 28720 4764
rect 1344 4678 8018 4730
rect 8070 4678 8122 4730
rect 8174 4678 8226 4730
rect 8278 4678 14822 4730
rect 14874 4678 14926 4730
rect 14978 4678 15030 4730
rect 15082 4678 21626 4730
rect 21678 4678 21730 4730
rect 21782 4678 21834 4730
rect 21886 4678 28430 4730
rect 28482 4678 28534 4730
rect 28586 4678 28638 4730
rect 28690 4678 28720 4730
rect 1344 4644 28720 4678
rect 10334 4562 10386 4574
rect 10334 4498 10386 4510
rect 11902 4562 11954 4574
rect 11902 4498 11954 4510
rect 23998 4562 24050 4574
rect 23998 4498 24050 4510
rect 26238 4562 26290 4574
rect 26238 4498 26290 4510
rect 26910 4562 26962 4574
rect 26910 4498 26962 4510
rect 27694 4562 27746 4574
rect 27694 4498 27746 4510
rect 24670 4450 24722 4462
rect 24670 4386 24722 4398
rect 25230 4450 25282 4462
rect 25230 4386 25282 4398
rect 25566 4450 25618 4462
rect 25566 4386 25618 4398
rect 25902 4450 25954 4462
rect 25902 4386 25954 4398
rect 24334 4338 24386 4350
rect 12114 4286 12126 4338
rect 12178 4286 12190 4338
rect 23762 4286 23774 4338
rect 23826 4286 23838 4338
rect 24334 4274 24386 4286
rect 8990 4226 9042 4238
rect 8990 4162 9042 4174
rect 9662 4226 9714 4238
rect 9662 4162 9714 4174
rect 11566 4226 11618 4238
rect 11566 4162 11618 4174
rect 20414 4226 20466 4238
rect 20414 4162 20466 4174
rect 23438 4226 23490 4238
rect 23438 4162 23490 4174
rect 11118 4114 11170 4126
rect 11118 4050 11170 4062
rect 1344 3946 28560 3980
rect 1344 3894 4616 3946
rect 4668 3894 4720 3946
rect 4772 3894 4824 3946
rect 4876 3894 11420 3946
rect 11472 3894 11524 3946
rect 11576 3894 11628 3946
rect 11680 3894 18224 3946
rect 18276 3894 18328 3946
rect 18380 3894 18432 3946
rect 18484 3894 25028 3946
rect 25080 3894 25132 3946
rect 25184 3894 25236 3946
rect 25288 3894 28560 3946
rect 1344 3860 28560 3894
rect 25454 3778 25506 3790
rect 25454 3714 25506 3726
rect 27358 3778 27410 3790
rect 27358 3714 27410 3726
rect 11442 3614 11454 3666
rect 11506 3614 11518 3666
rect 13570 3614 13582 3666
rect 13634 3614 13646 3666
rect 21522 3614 21534 3666
rect 21586 3614 21598 3666
rect 11006 3554 11058 3566
rect 8530 3502 8542 3554
rect 8594 3502 8606 3554
rect 11006 3490 11058 3502
rect 13134 3554 13186 3566
rect 21086 3554 21138 3566
rect 26574 3554 26626 3566
rect 19954 3502 19966 3554
rect 20018 3502 20030 3554
rect 23090 3502 23102 3554
rect 23154 3502 23166 3554
rect 23762 3502 23774 3554
rect 23826 3502 23838 3554
rect 26114 3502 26126 3554
rect 26178 3502 26190 3554
rect 13134 3490 13186 3502
rect 21086 3490 21138 3502
rect 26574 3490 26626 3502
rect 9662 3442 9714 3454
rect 9662 3378 9714 3390
rect 9998 3442 10050 3454
rect 9998 3378 10050 3390
rect 20190 3442 20242 3454
rect 20190 3378 20242 3390
rect 22766 3442 22818 3454
rect 22766 3378 22818 3390
rect 23326 3442 23378 3454
rect 23326 3378 23378 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 24894 3442 24946 3454
rect 24894 3378 24946 3390
rect 8766 3330 8818 3342
rect 8766 3266 8818 3278
rect 1344 3162 28720 3196
rect 1344 3110 8018 3162
rect 8070 3110 8122 3162
rect 8174 3110 8226 3162
rect 8278 3110 14822 3162
rect 14874 3110 14926 3162
rect 14978 3110 15030 3162
rect 15082 3110 21626 3162
rect 21678 3110 21730 3162
rect 21782 3110 21834 3162
rect 21886 3110 28430 3162
rect 28482 3110 28534 3162
rect 28586 3110 28638 3162
rect 28690 3110 28720 3162
rect 1344 3076 28720 3110
<< via1 >>
rect 8542 26798 8594 26850
rect 9438 26798 9490 26850
rect 10110 26798 10162 26850
rect 11118 26798 11170 26850
rect 16830 26798 16882 26850
rect 18286 26798 18338 26850
rect 22206 26798 22258 26850
rect 23214 26798 23266 26850
rect 23550 26798 23602 26850
rect 25006 26798 25058 26850
rect 8018 26630 8070 26682
rect 8122 26630 8174 26682
rect 8226 26630 8278 26682
rect 14822 26630 14874 26682
rect 14926 26630 14978 26682
rect 15030 26630 15082 26682
rect 21626 26630 21678 26682
rect 21730 26630 21782 26682
rect 21834 26630 21886 26682
rect 28430 26630 28482 26682
rect 28534 26630 28586 26682
rect 28638 26630 28690 26682
rect 3726 26462 3778 26514
rect 9438 26462 9490 26514
rect 15822 26462 15874 26514
rect 18286 26462 18338 26514
rect 20302 26462 20354 26514
rect 23214 26462 23266 26514
rect 6078 26350 6130 26402
rect 6750 26350 6802 26402
rect 7422 26350 7474 26402
rect 8094 26350 8146 26402
rect 8766 26350 8818 26402
rect 10670 26350 10722 26402
rect 12238 26350 12290 26402
rect 20750 26350 20802 26402
rect 21422 26350 21474 26402
rect 2942 26238 2994 26290
rect 4398 26238 4450 26290
rect 5854 26238 5906 26290
rect 6414 26238 6466 26290
rect 7198 26238 7250 26290
rect 7870 26238 7922 26290
rect 8542 26238 8594 26290
rect 9774 26238 9826 26290
rect 11342 26238 11394 26290
rect 13134 26238 13186 26290
rect 15038 26238 15090 26290
rect 17614 26238 17666 26290
rect 18622 26238 18674 26290
rect 20974 26238 21026 26290
rect 21646 26238 21698 26290
rect 22430 26238 22482 26290
rect 24558 26238 24610 26290
rect 26574 26238 26626 26290
rect 1934 26126 1986 26178
rect 3390 26126 3442 26178
rect 13582 26126 13634 26178
rect 19070 26126 19122 26178
rect 25006 26126 25058 26178
rect 27694 26126 27746 26178
rect 4616 25846 4668 25898
rect 4720 25846 4772 25898
rect 4824 25846 4876 25898
rect 11420 25846 11472 25898
rect 11524 25846 11576 25898
rect 11628 25846 11680 25898
rect 18224 25846 18276 25898
rect 18328 25846 18380 25898
rect 18432 25846 18484 25898
rect 25028 25846 25080 25898
rect 25132 25846 25184 25898
rect 25236 25846 25288 25898
rect 15038 25678 15090 25730
rect 15374 25678 15426 25730
rect 1822 25566 1874 25618
rect 5182 25566 5234 25618
rect 6414 25566 6466 25618
rect 6974 25566 7026 25618
rect 7646 25566 7698 25618
rect 8318 25566 8370 25618
rect 11118 25566 11170 25618
rect 12126 25566 12178 25618
rect 15038 25566 15090 25618
rect 15486 25566 15538 25618
rect 17502 25566 17554 25618
rect 18846 25566 18898 25618
rect 20414 25566 20466 25618
rect 20862 25566 20914 25618
rect 23550 25566 23602 25618
rect 25342 25566 25394 25618
rect 3278 25454 3330 25506
rect 3950 25454 4002 25506
rect 5630 25454 5682 25506
rect 15934 25454 15986 25506
rect 16382 25454 16434 25506
rect 17726 25454 17778 25506
rect 19070 25454 19122 25506
rect 21646 25454 21698 25506
rect 5966 25342 6018 25394
rect 13694 25342 13746 25394
rect 14366 25342 14418 25394
rect 21982 25342 22034 25394
rect 23102 25342 23154 25394
rect 26238 25342 26290 25394
rect 2158 25230 2210 25282
rect 2942 25230 2994 25282
rect 3614 25230 3666 25282
rect 4286 25230 4338 25282
rect 10558 25230 10610 25282
rect 11678 25230 11730 25282
rect 15710 25230 15762 25282
rect 16718 25230 16770 25282
rect 18062 25230 18114 25282
rect 19406 25230 19458 25282
rect 21310 25230 21362 25282
rect 24670 25230 24722 25282
rect 26574 25230 26626 25282
rect 26910 25230 26962 25282
rect 27694 25230 27746 25282
rect 28254 25230 28306 25282
rect 8018 25062 8070 25114
rect 8122 25062 8174 25114
rect 8226 25062 8278 25114
rect 14822 25062 14874 25114
rect 14926 25062 14978 25114
rect 15030 25062 15082 25114
rect 21626 25062 21678 25114
rect 21730 25062 21782 25114
rect 21834 25062 21886 25114
rect 28430 25062 28482 25114
rect 28534 25062 28586 25114
rect 28638 25062 28690 25114
rect 2158 24894 2210 24946
rect 3614 24894 3666 24946
rect 4622 24894 4674 24946
rect 10110 24894 10162 24946
rect 21198 24894 21250 24946
rect 24110 24894 24162 24946
rect 26126 24894 26178 24946
rect 28142 24894 28194 24946
rect 2942 24782 2994 24834
rect 4958 24782 5010 24834
rect 24670 24782 24722 24834
rect 3838 24670 3890 24722
rect 4286 24670 4338 24722
rect 5182 24670 5234 24722
rect 10894 24670 10946 24722
rect 20974 24670 21026 24722
rect 24446 24670 24498 24722
rect 25342 24670 25394 24722
rect 26910 24670 26962 24722
rect 27694 24670 27746 24722
rect 1822 24558 1874 24610
rect 4616 24278 4668 24330
rect 4720 24278 4772 24330
rect 4824 24278 4876 24330
rect 11420 24278 11472 24330
rect 11524 24278 11576 24330
rect 11628 24278 11680 24330
rect 18224 24278 18276 24330
rect 18328 24278 18380 24330
rect 18432 24278 18484 24330
rect 25028 24278 25080 24330
rect 25132 24278 25184 24330
rect 25236 24278 25288 24330
rect 3166 23998 3218 24050
rect 27582 23998 27634 24050
rect 2382 23886 2434 23938
rect 4174 23886 4226 23938
rect 4958 23886 5010 23938
rect 9326 23886 9378 23938
rect 10110 23886 10162 23938
rect 10670 23886 10722 23938
rect 11342 23886 11394 23938
rect 12126 23886 12178 23938
rect 17166 23886 17218 23938
rect 17950 23886 18002 23938
rect 20526 23886 20578 23938
rect 21422 23886 21474 23938
rect 24110 23886 24162 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 2718 23774 2770 23826
rect 3950 23774 4002 23826
rect 6078 23774 6130 23826
rect 9662 23774 9714 23826
rect 10334 23774 10386 23826
rect 11006 23774 11058 23826
rect 11678 23774 11730 23826
rect 12350 23774 12402 23826
rect 17502 23774 17554 23826
rect 18174 23774 18226 23826
rect 20750 23774 20802 23826
rect 21646 23774 21698 23826
rect 24334 23774 24386 23826
rect 24782 23774 24834 23826
rect 25454 23774 25506 23826
rect 25790 23774 25842 23826
rect 26126 23774 26178 23826
rect 4734 23662 4786 23714
rect 5742 23662 5794 23714
rect 25118 23662 25170 23714
rect 26462 23662 26514 23714
rect 26910 23662 26962 23714
rect 28254 23662 28306 23714
rect 8018 23494 8070 23546
rect 8122 23494 8174 23546
rect 8226 23494 8278 23546
rect 14822 23494 14874 23546
rect 14926 23494 14978 23546
rect 15030 23494 15082 23546
rect 21626 23494 21678 23546
rect 21730 23494 21782 23546
rect 21834 23494 21886 23546
rect 28430 23494 28482 23546
rect 28534 23494 28586 23546
rect 28638 23494 28690 23546
rect 2046 23326 2098 23378
rect 10558 23326 10610 23378
rect 11230 23326 11282 23378
rect 20974 23326 21026 23378
rect 26462 23326 26514 23378
rect 27134 23326 27186 23378
rect 20638 23214 20690 23266
rect 25790 23214 25842 23266
rect 26126 23214 26178 23266
rect 27470 23214 27522 23266
rect 27806 23214 27858 23266
rect 28142 23214 28194 23266
rect 1710 23102 1762 23154
rect 10782 23102 10834 23154
rect 11454 23102 11506 23154
rect 25566 23102 25618 23154
rect 2494 22990 2546 23042
rect 4616 22710 4668 22762
rect 4720 22710 4772 22762
rect 4824 22710 4876 22762
rect 11420 22710 11472 22762
rect 11524 22710 11576 22762
rect 11628 22710 11680 22762
rect 18224 22710 18276 22762
rect 18328 22710 18380 22762
rect 18432 22710 18484 22762
rect 25028 22710 25080 22762
rect 25132 22710 25184 22762
rect 25236 22710 25288 22762
rect 2942 22318 2994 22370
rect 28030 22318 28082 22370
rect 26462 22206 26514 22258
rect 26798 22206 26850 22258
rect 27134 22206 27186 22258
rect 27470 22206 27522 22258
rect 27806 22206 27858 22258
rect 2158 22094 2210 22146
rect 8018 21926 8070 21978
rect 8122 21926 8174 21978
rect 8226 21926 8278 21978
rect 14822 21926 14874 21978
rect 14926 21926 14978 21978
rect 15030 21926 15082 21978
rect 21626 21926 21678 21978
rect 21730 21926 21782 21978
rect 21834 21926 21886 21978
rect 28430 21926 28482 21978
rect 28534 21926 28586 21978
rect 28638 21926 28690 21978
rect 2942 21758 2994 21810
rect 27470 21758 27522 21810
rect 27806 21758 27858 21810
rect 22206 21646 22258 21698
rect 28142 21534 28194 21586
rect 2270 21422 2322 21474
rect 21198 21422 21250 21474
rect 27134 21422 27186 21474
rect 4616 21142 4668 21194
rect 4720 21142 4772 21194
rect 4824 21142 4876 21194
rect 11420 21142 11472 21194
rect 11524 21142 11576 21194
rect 11628 21142 11680 21194
rect 18224 21142 18276 21194
rect 18328 21142 18380 21194
rect 18432 21142 18484 21194
rect 25028 21142 25080 21194
rect 25132 21142 25184 21194
rect 25236 21142 25288 21194
rect 14478 20862 14530 20914
rect 1822 20750 1874 20802
rect 19070 20750 19122 20802
rect 26910 20750 26962 20802
rect 2046 20638 2098 20690
rect 2382 20638 2434 20690
rect 15486 20638 15538 20690
rect 28030 20638 28082 20690
rect 19294 20526 19346 20578
rect 8018 20358 8070 20410
rect 8122 20358 8174 20410
rect 8226 20358 8278 20410
rect 14822 20358 14874 20410
rect 14926 20358 14978 20410
rect 15030 20358 15082 20410
rect 21626 20358 21678 20410
rect 21730 20358 21782 20410
rect 21834 20358 21886 20410
rect 28430 20358 28482 20410
rect 28534 20358 28586 20410
rect 28638 20358 28690 20410
rect 1822 20190 1874 20242
rect 14366 20078 14418 20130
rect 19406 20078 19458 20130
rect 22206 20078 22258 20130
rect 11454 19966 11506 20018
rect 12126 19966 12178 20018
rect 16158 19966 16210 20018
rect 26910 19966 26962 20018
rect 18398 19854 18450 19906
rect 21198 19854 21250 19906
rect 28030 19854 28082 19906
rect 15150 19742 15202 19794
rect 16046 19742 16098 19794
rect 4616 19574 4668 19626
rect 4720 19574 4772 19626
rect 4824 19574 4876 19626
rect 11420 19574 11472 19626
rect 11524 19574 11576 19626
rect 11628 19574 11680 19626
rect 18224 19574 18276 19626
rect 18328 19574 18380 19626
rect 18432 19574 18484 19626
rect 25028 19574 25080 19626
rect 25132 19574 25184 19626
rect 25236 19574 25288 19626
rect 20638 19406 20690 19458
rect 8654 19294 8706 19346
rect 11454 19294 11506 19346
rect 15262 19294 15314 19346
rect 17166 19182 17218 19234
rect 17614 19182 17666 19234
rect 23214 19182 23266 19234
rect 23886 19182 23938 19234
rect 9662 19070 9714 19122
rect 12462 19070 12514 19122
rect 16270 19070 16322 19122
rect 19854 19070 19906 19122
rect 27470 19070 27522 19122
rect 27806 19070 27858 19122
rect 28142 19070 28194 19122
rect 26126 18958 26178 19010
rect 26910 18958 26962 19010
rect 27134 18958 27186 19010
rect 8018 18790 8070 18842
rect 8122 18790 8174 18842
rect 8226 18790 8278 18842
rect 14822 18790 14874 18842
rect 14926 18790 14978 18842
rect 15030 18790 15082 18842
rect 21626 18790 21678 18842
rect 21730 18790 21782 18842
rect 21834 18790 21886 18842
rect 28430 18790 28482 18842
rect 28534 18790 28586 18842
rect 28638 18790 28690 18842
rect 8430 18622 8482 18674
rect 12574 18622 12626 18674
rect 16158 18622 16210 18674
rect 28254 18622 28306 18674
rect 7646 18510 7698 18562
rect 21646 18510 21698 18562
rect 27246 18510 27298 18562
rect 4958 18398 5010 18450
rect 5406 18398 5458 18450
rect 9438 18398 9490 18450
rect 10110 18398 10162 18450
rect 13246 18398 13298 18450
rect 13918 18398 13970 18450
rect 16942 18398 16994 18450
rect 18174 18398 18226 18450
rect 18734 18398 18786 18450
rect 19294 18398 19346 18450
rect 22430 18398 22482 18450
rect 23774 18398 23826 18450
rect 13134 18286 13186 18338
rect 23102 18286 23154 18338
rect 26238 18286 26290 18338
rect 18062 18174 18114 18226
rect 23998 18174 24050 18226
rect 4616 18006 4668 18058
rect 4720 18006 4772 18058
rect 4824 18006 4876 18058
rect 11420 18006 11472 18058
rect 11524 18006 11576 18058
rect 11628 18006 11680 18058
rect 18224 18006 18276 18058
rect 18328 18006 18380 18058
rect 18432 18006 18484 18058
rect 25028 18006 25080 18058
rect 25132 18006 25184 18058
rect 25236 18006 25288 18058
rect 6302 17838 6354 17890
rect 10782 17838 10834 17890
rect 12574 17838 12626 17890
rect 14142 17838 14194 17890
rect 18958 17838 19010 17890
rect 20078 17726 20130 17778
rect 26126 17726 26178 17778
rect 4734 17614 4786 17666
rect 6862 17614 6914 17666
rect 7086 17614 7138 17666
rect 7758 17614 7810 17666
rect 12686 17614 12738 17666
rect 14142 17614 14194 17666
rect 15262 17614 15314 17666
rect 15934 17614 15986 17666
rect 19630 17614 19682 17666
rect 21198 17614 21250 17666
rect 21870 17614 21922 17666
rect 4846 17502 4898 17554
rect 18174 17502 18226 17554
rect 24110 17502 24162 17554
rect 27134 17502 27186 17554
rect 9998 17390 10050 17442
rect 24894 17390 24946 17442
rect 8018 17222 8070 17274
rect 8122 17222 8174 17274
rect 8226 17222 8278 17274
rect 14822 17222 14874 17274
rect 14926 17222 14978 17274
rect 15030 17222 15082 17274
rect 21626 17222 21678 17274
rect 21730 17222 21782 17274
rect 21834 17222 21886 17274
rect 28430 17222 28482 17274
rect 28534 17222 28586 17274
rect 28638 17222 28690 17274
rect 5854 17054 5906 17106
rect 9774 16942 9826 16994
rect 21422 16942 21474 16994
rect 27246 16942 27298 16994
rect 3166 16830 3218 16882
rect 3614 16830 3666 16882
rect 7534 16830 7586 16882
rect 14702 16830 14754 16882
rect 19518 16830 19570 16882
rect 26238 16718 26290 16770
rect 6638 16606 6690 16658
rect 7310 16606 7362 16658
rect 4616 16438 4668 16490
rect 4720 16438 4772 16490
rect 4824 16438 4876 16490
rect 11420 16438 11472 16490
rect 11524 16438 11576 16490
rect 11628 16438 11680 16490
rect 18224 16438 18276 16490
rect 18328 16438 18380 16490
rect 18432 16438 18484 16490
rect 25028 16438 25080 16490
rect 25132 16438 25184 16490
rect 25236 16438 25288 16490
rect 3838 16158 3890 16210
rect 6190 16158 6242 16210
rect 9998 16158 10050 16210
rect 26686 16158 26738 16210
rect 12910 16046 12962 16098
rect 13694 16046 13746 16098
rect 19070 16046 19122 16098
rect 19406 16046 19458 16098
rect 19854 16046 19906 16098
rect 24334 16046 24386 16098
rect 24670 16046 24722 16098
rect 2718 15934 2770 15986
rect 7310 15934 7362 15986
rect 11118 15934 11170 15986
rect 27694 15934 27746 15986
rect 12350 15822 12402 15874
rect 13582 15822 13634 15874
rect 15934 15822 15986 15874
rect 16718 15822 16770 15874
rect 20414 15822 20466 15874
rect 21198 15822 21250 15874
rect 21982 15822 22034 15874
rect 25230 15822 25282 15874
rect 8018 15654 8070 15706
rect 8122 15654 8174 15706
rect 8226 15654 8278 15706
rect 14822 15654 14874 15706
rect 14926 15654 14978 15706
rect 15030 15654 15082 15706
rect 21626 15654 21678 15706
rect 21730 15654 21782 15706
rect 21834 15654 21886 15706
rect 28430 15654 28482 15706
rect 28534 15654 28586 15706
rect 28638 15654 28690 15706
rect 1934 15486 1986 15538
rect 11118 15486 11170 15538
rect 11902 15486 11954 15538
rect 16718 15486 16770 15538
rect 24558 15486 24610 15538
rect 27694 15486 27746 15538
rect 2718 15374 2770 15426
rect 7982 15374 8034 15426
rect 9886 15374 9938 15426
rect 17502 15374 17554 15426
rect 22318 15374 22370 15426
rect 4958 15262 5010 15314
rect 5406 15262 5458 15314
rect 10222 15262 10274 15314
rect 14142 15262 14194 15314
rect 14590 15262 14642 15314
rect 16494 15262 16546 15314
rect 24334 15262 24386 15314
rect 25678 15262 25730 15314
rect 27022 15262 27074 15314
rect 6974 15150 7026 15202
rect 18622 15150 18674 15202
rect 21310 15150 21362 15202
rect 23550 15150 23602 15202
rect 25566 15150 25618 15202
rect 4616 14870 4668 14922
rect 4720 14870 4772 14922
rect 4824 14870 4876 14922
rect 11420 14870 11472 14922
rect 11524 14870 11576 14922
rect 11628 14870 11680 14922
rect 18224 14870 18276 14922
rect 18328 14870 18380 14922
rect 18432 14870 18484 14922
rect 25028 14870 25080 14922
rect 25132 14870 25184 14922
rect 25236 14870 25288 14922
rect 3950 14702 4002 14754
rect 26350 14702 26402 14754
rect 8094 14590 8146 14642
rect 14254 14590 14306 14642
rect 19518 14590 19570 14642
rect 26910 14590 26962 14642
rect 4174 14478 4226 14530
rect 9550 14478 9602 14530
rect 9998 14478 10050 14530
rect 14478 14478 14530 14530
rect 22094 14478 22146 14530
rect 22766 14478 22818 14530
rect 23326 14478 23378 14530
rect 26574 14478 26626 14530
rect 28142 14478 28194 14530
rect 6750 14366 6802 14418
rect 25566 14366 25618 14418
rect 27806 14366 27858 14418
rect 12350 14254 12402 14306
rect 13022 14254 13074 14306
rect 20750 14254 20802 14306
rect 22318 14254 22370 14306
rect 8018 14086 8070 14138
rect 8122 14086 8174 14138
rect 8226 14086 8278 14138
rect 14822 14086 14874 14138
rect 14926 14086 14978 14138
rect 15030 14086 15082 14138
rect 21626 14086 21678 14138
rect 21730 14086 21782 14138
rect 21834 14086 21886 14138
rect 28430 14086 28482 14138
rect 28534 14086 28586 14138
rect 28638 14086 28690 14138
rect 5406 13918 5458 13970
rect 6190 13918 6242 13970
rect 20526 13918 20578 13970
rect 28254 13918 28306 13970
rect 2382 13806 2434 13858
rect 11790 13806 11842 13858
rect 13918 13806 13970 13858
rect 21310 13806 21362 13858
rect 22766 13806 22818 13858
rect 4734 13694 4786 13746
rect 5182 13694 5234 13746
rect 8430 13694 8482 13746
rect 8990 13694 9042 13746
rect 17614 13694 17666 13746
rect 18286 13694 18338 13746
rect 10782 13582 10834 13634
rect 15038 13582 15090 13634
rect 21982 13582 22034 13634
rect 25902 13582 25954 13634
rect 26238 13582 26290 13634
rect 1598 13470 1650 13522
rect 4616 13302 4668 13354
rect 4720 13302 4772 13354
rect 4824 13302 4876 13354
rect 11420 13302 11472 13354
rect 11524 13302 11576 13354
rect 11628 13302 11680 13354
rect 18224 13302 18276 13354
rect 18328 13302 18380 13354
rect 18432 13302 18484 13354
rect 25028 13302 25080 13354
rect 25132 13302 25184 13354
rect 25236 13302 25288 13354
rect 3278 13134 3330 13186
rect 9214 13134 9266 13186
rect 16382 13134 16434 13186
rect 3390 12910 3442 12962
rect 4622 12910 4674 12962
rect 5518 12910 5570 12962
rect 6190 12910 6242 12962
rect 12462 12910 12514 12962
rect 12798 12910 12850 12962
rect 18734 12910 18786 12962
rect 22206 12910 22258 12962
rect 22654 12910 22706 12962
rect 25902 12910 25954 12962
rect 1710 12798 1762 12850
rect 2046 12686 2098 12738
rect 2494 12686 2546 12738
rect 4398 12686 4450 12738
rect 8654 12686 8706 12738
rect 9326 12686 9378 12738
rect 10110 12686 10162 12738
rect 21422 12686 21474 12738
rect 25118 12686 25170 12738
rect 25678 12686 25730 12738
rect 26014 12686 26066 12738
rect 8018 12518 8070 12570
rect 8122 12518 8174 12570
rect 8226 12518 8278 12570
rect 14822 12518 14874 12570
rect 14926 12518 14978 12570
rect 15030 12518 15082 12570
rect 21626 12518 21678 12570
rect 21730 12518 21782 12570
rect 21834 12518 21886 12570
rect 28430 12518 28482 12570
rect 28534 12518 28586 12570
rect 28638 12518 28690 12570
rect 3502 12350 3554 12402
rect 4286 12350 4338 12402
rect 8654 12238 8706 12290
rect 9774 12238 9826 12290
rect 27246 12238 27298 12290
rect 2046 12126 2098 12178
rect 2494 12126 2546 12178
rect 3278 12126 3330 12178
rect 6638 12126 6690 12178
rect 6974 12126 7026 12178
rect 8542 12126 8594 12178
rect 14814 12126 14866 12178
rect 19518 12126 19570 12178
rect 18734 12014 18786 12066
rect 19070 12014 19122 12066
rect 24446 12014 24498 12066
rect 25566 12014 25618 12066
rect 26238 12014 26290 12066
rect 3166 11902 3218 11954
rect 4616 11734 4668 11786
rect 4720 11734 4772 11786
rect 4824 11734 4876 11786
rect 11420 11734 11472 11786
rect 11524 11734 11576 11786
rect 11628 11734 11680 11786
rect 18224 11734 18276 11786
rect 18328 11734 18380 11786
rect 18432 11734 18484 11786
rect 25028 11734 25080 11786
rect 25132 11734 25184 11786
rect 25236 11734 25288 11786
rect 9102 11566 9154 11618
rect 24894 11566 24946 11618
rect 3726 11454 3778 11506
rect 16270 11454 16322 11506
rect 19294 11454 19346 11506
rect 25230 11454 25282 11506
rect 26686 11454 26738 11506
rect 5966 11342 6018 11394
rect 12686 11342 12738 11394
rect 21422 11342 21474 11394
rect 21870 11342 21922 11394
rect 2606 11230 2658 11282
rect 17278 11230 17330 11282
rect 20302 11230 20354 11282
rect 24110 11230 24162 11282
rect 27694 11230 27746 11282
rect 5742 11118 5794 11170
rect 8018 10950 8070 11002
rect 8122 10950 8174 11002
rect 8226 10950 8278 11002
rect 14822 10950 14874 11002
rect 14926 10950 14978 11002
rect 15030 10950 15082 11002
rect 21626 10950 21678 11002
rect 21730 10950 21782 11002
rect 21834 10950 21886 11002
rect 28430 10950 28482 11002
rect 28534 10950 28586 11002
rect 28638 10950 28690 11002
rect 5518 10782 5570 10834
rect 16270 10782 16322 10834
rect 20190 10782 20242 10834
rect 25342 10782 25394 10834
rect 25790 10782 25842 10834
rect 2046 10670 2098 10722
rect 6078 10670 6130 10722
rect 6414 10670 6466 10722
rect 11790 10670 11842 10722
rect 15486 10670 15538 10722
rect 23998 10670 24050 10722
rect 27246 10670 27298 10722
rect 1822 10558 1874 10610
rect 2382 10558 2434 10610
rect 3054 10558 3106 10610
rect 12798 10558 12850 10610
rect 13246 10558 13298 10610
rect 17278 10558 17330 10610
rect 17950 10558 18002 10610
rect 21310 10558 21362 10610
rect 21758 10558 21810 10610
rect 7534 10446 7586 10498
rect 10782 10446 10834 10498
rect 16494 10446 16546 10498
rect 16830 10446 16882 10498
rect 26238 10446 26290 10498
rect 20974 10334 21026 10386
rect 24782 10334 24834 10386
rect 4616 10166 4668 10218
rect 4720 10166 4772 10218
rect 4824 10166 4876 10218
rect 11420 10166 11472 10218
rect 11524 10166 11576 10218
rect 11628 10166 11680 10218
rect 18224 10166 18276 10218
rect 18328 10166 18380 10218
rect 18432 10166 18484 10218
rect 25028 10166 25080 10218
rect 25132 10166 25184 10218
rect 25236 10166 25288 10218
rect 18958 9998 19010 10050
rect 25566 9998 25618 10050
rect 27694 9998 27746 10050
rect 1822 9886 1874 9938
rect 6638 9886 6690 9938
rect 15038 9886 15090 9938
rect 19182 9886 19234 9938
rect 21422 9886 21474 9938
rect 9550 9774 9602 9826
rect 9998 9774 10050 9826
rect 14142 9774 14194 9826
rect 14702 9774 14754 9826
rect 15486 9774 15538 9826
rect 15934 9774 15986 9826
rect 19966 9774 20018 9826
rect 21870 9774 21922 9826
rect 22542 9774 22594 9826
rect 25790 9774 25842 9826
rect 26910 9774 26962 9826
rect 7646 9662 7698 9714
rect 13918 9662 13970 9714
rect 12462 9550 12514 9602
rect 13022 9550 13074 9602
rect 18398 9550 18450 9602
rect 19294 9550 19346 9602
rect 24782 9550 24834 9602
rect 25902 9550 25954 9602
rect 8018 9382 8070 9434
rect 8122 9382 8174 9434
rect 8226 9382 8278 9434
rect 14822 9382 14874 9434
rect 14926 9382 14978 9434
rect 15030 9382 15082 9434
rect 21626 9382 21678 9434
rect 21730 9382 21782 9434
rect 21834 9382 21886 9434
rect 28430 9382 28482 9434
rect 28534 9382 28586 9434
rect 28638 9382 28690 9434
rect 4958 9214 5010 9266
rect 5518 9214 5570 9266
rect 16382 9214 16434 9266
rect 21646 9214 21698 9266
rect 23550 9214 23602 9266
rect 24558 9214 24610 9266
rect 25454 9214 25506 9266
rect 12462 9102 12514 9154
rect 27246 9102 27298 9154
rect 2046 8990 2098 9042
rect 2494 8990 2546 9042
rect 9774 8990 9826 9042
rect 12686 8990 12738 9042
rect 13246 8990 13298 9042
rect 13806 8990 13858 9042
rect 17950 8990 18002 9042
rect 24334 8990 24386 9042
rect 11902 8878 11954 8930
rect 26238 8878 26290 8930
rect 16942 8766 16994 8818
rect 4616 8598 4668 8650
rect 4720 8598 4772 8650
rect 4824 8598 4876 8650
rect 11420 8598 11472 8650
rect 11524 8598 11576 8650
rect 11628 8598 11680 8650
rect 18224 8598 18276 8650
rect 18328 8598 18380 8650
rect 18432 8598 18484 8650
rect 25028 8598 25080 8650
rect 25132 8598 25184 8650
rect 25236 8598 25288 8650
rect 14478 8318 14530 8370
rect 17614 8318 17666 8370
rect 26574 8318 26626 8370
rect 27694 8318 27746 8370
rect 2942 8206 2994 8258
rect 3390 8206 3442 8258
rect 22990 8206 23042 8258
rect 23550 8206 23602 8258
rect 27022 8206 27074 8258
rect 2046 8094 2098 8146
rect 4062 8094 4114 8146
rect 15486 8094 15538 8146
rect 18622 8094 18674 8146
rect 3614 7982 3666 8034
rect 25902 7982 25954 8034
rect 8018 7814 8070 7866
rect 8122 7814 8174 7866
rect 8226 7814 8278 7866
rect 14822 7814 14874 7866
rect 14926 7814 14978 7866
rect 15030 7814 15082 7866
rect 21626 7814 21678 7866
rect 21730 7814 21782 7866
rect 21834 7814 21886 7866
rect 28430 7814 28482 7866
rect 28534 7814 28586 7866
rect 28638 7814 28690 7866
rect 23998 7646 24050 7698
rect 22094 7534 22146 7586
rect 25342 7534 25394 7586
rect 2942 7422 2994 7474
rect 23998 7422 24050 7474
rect 1934 7310 1986 7362
rect 20750 7310 20802 7362
rect 23550 7310 23602 7362
rect 26462 7310 26514 7362
rect 27134 7310 27186 7362
rect 27806 7310 27858 7362
rect 27470 7198 27522 7250
rect 27806 7198 27858 7250
rect 4616 7030 4668 7082
rect 4720 7030 4772 7082
rect 4824 7030 4876 7082
rect 11420 7030 11472 7082
rect 11524 7030 11576 7082
rect 11628 7030 11680 7082
rect 18224 7030 18276 7082
rect 18328 7030 18380 7082
rect 18432 7030 18484 7082
rect 25028 7030 25080 7082
rect 25132 7030 25184 7082
rect 25236 7030 25288 7082
rect 23102 6862 23154 6914
rect 3390 6638 3442 6690
rect 4734 6638 4786 6690
rect 22990 6638 23042 6690
rect 26238 6638 26290 6690
rect 26798 6638 26850 6690
rect 28142 6638 28194 6690
rect 1710 6526 1762 6578
rect 2046 6526 2098 6578
rect 3838 6526 3890 6578
rect 4174 6526 4226 6578
rect 27470 6526 27522 6578
rect 27806 6526 27858 6578
rect 2494 6414 2546 6466
rect 3166 6414 3218 6466
rect 4510 6414 4562 6466
rect 23886 6414 23938 6466
rect 27134 6414 27186 6466
rect 8018 6246 8070 6298
rect 8122 6246 8174 6298
rect 8226 6246 8278 6298
rect 14822 6246 14874 6298
rect 14926 6246 14978 6298
rect 15030 6246 15082 6298
rect 21626 6246 21678 6298
rect 21730 6246 21782 6298
rect 21834 6246 21886 6298
rect 28430 6246 28482 6298
rect 28534 6246 28586 6298
rect 28638 6246 28690 6298
rect 25454 6078 25506 6130
rect 27694 6078 27746 6130
rect 28254 6078 28306 6130
rect 10334 5966 10386 6018
rect 11118 5966 11170 6018
rect 23998 5966 24050 6018
rect 24670 5966 24722 6018
rect 2942 5854 2994 5906
rect 9998 5854 10050 5906
rect 10894 5854 10946 5906
rect 24334 5854 24386 5906
rect 25678 5854 25730 5906
rect 26910 5854 26962 5906
rect 1934 5742 1986 5794
rect 4616 5462 4668 5514
rect 4720 5462 4772 5514
rect 4824 5462 4876 5514
rect 11420 5462 11472 5514
rect 11524 5462 11576 5514
rect 11628 5462 11680 5514
rect 18224 5462 18276 5514
rect 18328 5462 18380 5514
rect 18432 5462 18484 5514
rect 25028 5462 25080 5514
rect 25132 5462 25184 5514
rect 25236 5462 25288 5514
rect 27582 5182 27634 5234
rect 1710 5070 1762 5122
rect 2494 5070 2546 5122
rect 9998 5070 10050 5122
rect 24334 5070 24386 5122
rect 24558 5070 24610 5122
rect 25342 5070 25394 5122
rect 25902 5070 25954 5122
rect 26910 5070 26962 5122
rect 2046 4958 2098 5010
rect 20414 4958 20466 5010
rect 10222 4846 10274 4898
rect 20750 4846 20802 4898
rect 24894 4846 24946 4898
rect 25566 4846 25618 4898
rect 26238 4846 26290 4898
rect 8018 4678 8070 4730
rect 8122 4678 8174 4730
rect 8226 4678 8278 4730
rect 14822 4678 14874 4730
rect 14926 4678 14978 4730
rect 15030 4678 15082 4730
rect 21626 4678 21678 4730
rect 21730 4678 21782 4730
rect 21834 4678 21886 4730
rect 28430 4678 28482 4730
rect 28534 4678 28586 4730
rect 28638 4678 28690 4730
rect 10334 4510 10386 4562
rect 11902 4510 11954 4562
rect 23998 4510 24050 4562
rect 26238 4510 26290 4562
rect 26910 4510 26962 4562
rect 27694 4510 27746 4562
rect 24670 4398 24722 4450
rect 25230 4398 25282 4450
rect 25566 4398 25618 4450
rect 25902 4398 25954 4450
rect 12126 4286 12178 4338
rect 23774 4286 23826 4338
rect 24334 4286 24386 4338
rect 8990 4174 9042 4226
rect 9662 4174 9714 4226
rect 11566 4174 11618 4226
rect 20414 4174 20466 4226
rect 23438 4174 23490 4226
rect 11118 4062 11170 4114
rect 4616 3894 4668 3946
rect 4720 3894 4772 3946
rect 4824 3894 4876 3946
rect 11420 3894 11472 3946
rect 11524 3894 11576 3946
rect 11628 3894 11680 3946
rect 18224 3894 18276 3946
rect 18328 3894 18380 3946
rect 18432 3894 18484 3946
rect 25028 3894 25080 3946
rect 25132 3894 25184 3946
rect 25236 3894 25288 3946
rect 25454 3726 25506 3778
rect 27358 3726 27410 3778
rect 11454 3614 11506 3666
rect 13582 3614 13634 3666
rect 21534 3614 21586 3666
rect 8542 3502 8594 3554
rect 11006 3502 11058 3554
rect 13134 3502 13186 3554
rect 19966 3502 20018 3554
rect 21086 3502 21138 3554
rect 23102 3502 23154 3554
rect 23774 3502 23826 3554
rect 26126 3502 26178 3554
rect 26574 3502 26626 3554
rect 9662 3390 9714 3442
rect 9998 3390 10050 3442
rect 20190 3390 20242 3442
rect 22766 3390 22818 3442
rect 23326 3390 23378 3442
rect 23998 3390 24050 3442
rect 24894 3390 24946 3442
rect 8766 3278 8818 3330
rect 8018 3110 8070 3162
rect 8122 3110 8174 3162
rect 8226 3110 8278 3162
rect 14822 3110 14874 3162
rect 14926 3110 14978 3162
rect 15030 3110 15082 3162
rect 21626 3110 21678 3162
rect 21730 3110 21782 3162
rect 21834 3110 21886 3162
rect 28430 3110 28482 3162
rect 28534 3110 28586 3162
rect 28638 3110 28690 3162
<< metal2 >>
rect 5376 29200 5488 30000
rect 6048 29200 6160 30000
rect 6720 29200 6832 30000
rect 7392 29200 7504 30000
rect 8064 29200 8176 30000
rect 8736 29200 8848 30000
rect 9408 29200 9520 30000
rect 10080 29200 10192 30000
rect 10752 29200 10864 30000
rect 11424 29200 11536 30000
rect 12096 29200 12208 30000
rect 12768 29200 12880 30000
rect 13440 29200 13552 30000
rect 14112 29200 14224 30000
rect 14784 29200 14896 30000
rect 15456 29200 15568 30000
rect 16128 29200 16240 30000
rect 16800 29200 16912 30000
rect 17472 29200 17584 30000
rect 18144 29200 18256 30000
rect 18816 29200 18928 30000
rect 19488 29204 19600 30000
rect 19740 29260 20020 29316
rect 19740 29204 19796 29260
rect 19488 29200 19796 29204
rect 1820 28308 1876 28318
rect 1820 25618 1876 28252
rect 3724 27636 3780 27646
rect 3388 26964 3444 26974
rect 2044 26292 2100 26302
rect 1820 25566 1822 25618
rect 1874 25566 1876 25618
rect 1820 25508 1876 25566
rect 1932 26178 1988 26190
rect 1932 26126 1934 26178
rect 1986 26126 1988 26178
rect 1932 25620 1988 26126
rect 1932 25554 1988 25564
rect 1820 25442 1876 25452
rect 2044 24948 2100 26236
rect 2940 26292 2996 26302
rect 2940 26198 2996 26236
rect 3388 26178 3444 26908
rect 3724 26514 3780 27580
rect 5404 26908 5460 29200
rect 6076 26964 6132 29200
rect 3724 26462 3726 26514
rect 3778 26462 3780 26514
rect 3724 26450 3780 26462
rect 5180 26852 5460 26908
rect 5852 26908 6468 26964
rect 6748 26908 6804 29200
rect 7420 26964 7476 29200
rect 8092 26964 8148 29200
rect 8764 27300 8820 29200
rect 7196 26908 7700 26964
rect 3948 26292 4004 26302
rect 4004 26236 4116 26292
rect 3948 26226 4004 26236
rect 3388 26126 3390 26178
rect 3442 26126 3444 26178
rect 3276 25508 3332 25518
rect 3388 25508 3444 26126
rect 3948 25508 4004 25518
rect 3388 25506 4004 25508
rect 3388 25454 3950 25506
rect 4002 25454 4004 25506
rect 3388 25452 4004 25454
rect 3276 25414 3332 25452
rect 3948 25442 4004 25452
rect 2156 25284 2212 25294
rect 2156 25190 2212 25228
rect 2940 25284 2996 25294
rect 2940 25190 2996 25228
rect 3500 25284 3556 25294
rect 2156 24948 2212 24958
rect 2044 24946 2212 24948
rect 2044 24894 2158 24946
rect 2210 24894 2212 24946
rect 2044 24892 2212 24894
rect 3500 24948 3556 25228
rect 3612 25284 3668 25294
rect 3612 25282 3892 25284
rect 3612 25230 3614 25282
rect 3666 25230 3892 25282
rect 3612 25228 3892 25230
rect 3612 25218 3668 25228
rect 3612 24948 3668 24958
rect 3500 24946 3668 24948
rect 3500 24894 3614 24946
rect 3666 24894 3668 24946
rect 3500 24892 3668 24894
rect 2156 24882 2212 24892
rect 3612 24882 3668 24892
rect 2940 24836 2996 24846
rect 2940 24742 2996 24780
rect 2716 24724 2772 24734
rect 1820 24610 1876 24622
rect 1820 24558 1822 24610
rect 1874 24558 1876 24610
rect 1708 23828 1764 23838
rect 1820 23828 1876 24558
rect 2380 24276 2436 24286
rect 2268 23940 2324 23950
rect 2156 23884 2268 23940
rect 1708 23826 1876 23828
rect 1708 23774 1710 23826
rect 1762 23774 1876 23826
rect 1708 23772 1876 23774
rect 2044 23828 2100 23838
rect 1708 23604 1764 23772
rect 2044 23734 2100 23772
rect 1708 23538 1764 23548
rect 2044 23380 2100 23390
rect 2156 23380 2212 23884
rect 2268 23874 2324 23884
rect 2380 23938 2436 24220
rect 2380 23886 2382 23938
rect 2434 23886 2436 23938
rect 2380 23874 2436 23886
rect 2716 23826 2772 24668
rect 3836 24722 3892 25228
rect 3836 24670 3838 24722
rect 3890 24670 3892 24722
rect 3836 24658 3892 24670
rect 3164 24276 3220 24286
rect 3164 24050 3220 24220
rect 3164 23998 3166 24050
rect 3218 23998 3220 24050
rect 3164 23986 3220 23998
rect 2716 23774 2718 23826
rect 2770 23774 2772 23826
rect 2716 23762 2772 23774
rect 3948 23828 4004 23838
rect 4060 23828 4116 26236
rect 4396 26290 4452 26302
rect 4396 26238 4398 26290
rect 4450 26238 4452 26290
rect 4284 25284 4340 25294
rect 4172 25282 4340 25284
rect 4172 25230 4286 25282
rect 4338 25230 4340 25282
rect 4172 25228 4340 25230
rect 4172 23938 4228 25228
rect 4284 25218 4340 25228
rect 4396 24948 4452 26238
rect 4614 25900 4878 25910
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4614 25834 4878 25844
rect 5180 25620 5236 26852
rect 5852 26290 5908 26908
rect 6412 26852 6580 26908
rect 6748 26852 7028 26908
rect 5852 26238 5854 26290
rect 5906 26238 5908 26290
rect 5852 26226 5908 26238
rect 6076 26402 6132 26414
rect 6076 26350 6078 26402
rect 6130 26350 6132 26402
rect 5180 25618 5684 25620
rect 5180 25566 5182 25618
rect 5234 25566 5684 25618
rect 5180 25564 5684 25566
rect 5180 25554 5236 25564
rect 5628 25506 5684 25564
rect 5628 25454 5630 25506
rect 5682 25454 5684 25506
rect 5628 25442 5684 25454
rect 6076 25508 6132 26350
rect 6412 26292 6468 26302
rect 6412 26198 6468 26236
rect 6412 25620 6468 25630
rect 6524 25620 6580 26852
rect 6412 25618 6580 25620
rect 6412 25566 6414 25618
rect 6466 25566 6580 25618
rect 6412 25564 6580 25566
rect 6748 26402 6804 26414
rect 6748 26350 6750 26402
rect 6802 26350 6804 26402
rect 6412 25554 6468 25564
rect 6076 25442 6132 25452
rect 5964 25396 6020 25406
rect 5964 25302 6020 25340
rect 6748 25284 6804 26350
rect 6972 26292 7028 26852
rect 6972 25618 7028 26236
rect 7196 26290 7252 26908
rect 7196 26238 7198 26290
rect 7250 26238 7252 26290
rect 7196 26226 7252 26238
rect 7420 26402 7476 26414
rect 7420 26350 7422 26402
rect 7474 26350 7476 26402
rect 6972 25566 6974 25618
rect 7026 25566 7028 25618
rect 6972 25554 7028 25566
rect 7420 25620 7476 26350
rect 7420 25554 7476 25564
rect 7644 25618 7700 26908
rect 7868 26908 8148 26964
rect 8540 27244 8820 27300
rect 7868 26292 7924 26908
rect 8540 26850 8596 27244
rect 9436 27076 9492 29200
rect 9436 27020 10052 27076
rect 8540 26798 8542 26850
rect 8594 26798 8596 26850
rect 8016 26684 8280 26694
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8016 26618 8280 26628
rect 8092 26404 8148 26414
rect 7868 26198 7924 26236
rect 7980 26402 8148 26404
rect 7980 26350 8094 26402
rect 8146 26350 8148 26402
rect 7980 26348 8148 26350
rect 7644 25566 7646 25618
rect 7698 25566 7700 25618
rect 7644 25554 7700 25566
rect 7980 25284 8036 26348
rect 8092 26338 8148 26348
rect 8316 26292 8372 26302
rect 8316 25618 8372 26236
rect 8540 26290 8596 26798
rect 9436 26850 9492 26862
rect 9436 26798 9438 26850
rect 9490 26798 9492 26850
rect 9436 26514 9492 26798
rect 9436 26462 9438 26514
rect 9490 26462 9492 26514
rect 9436 26450 9492 26462
rect 8764 26404 8820 26414
rect 8764 26310 8820 26348
rect 8540 26238 8542 26290
rect 8594 26238 8596 26290
rect 8540 26226 8596 26238
rect 9772 26290 9828 26302
rect 9772 26238 9774 26290
rect 9826 26238 9828 26290
rect 8316 25566 8318 25618
rect 8370 25566 8372 25618
rect 8316 25554 8372 25566
rect 6748 25218 6804 25228
rect 7868 25228 8036 25284
rect 9324 25284 9380 25294
rect 4620 24948 4676 24958
rect 4396 24946 4676 24948
rect 4396 24894 4622 24946
rect 4674 24894 4676 24946
rect 4396 24892 4676 24894
rect 4620 24882 4676 24892
rect 4956 24836 5012 24846
rect 4956 24742 5012 24780
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 5180 24722 5236 24734
rect 5180 24670 5182 24722
rect 5234 24670 5236 24722
rect 4614 24332 4878 24342
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4614 24266 4878 24276
rect 4172 23886 4174 23938
rect 4226 23886 4228 23938
rect 4172 23874 4228 23886
rect 4956 23940 5012 23950
rect 4956 23846 5012 23884
rect 3948 23826 4116 23828
rect 3948 23774 3950 23826
rect 4002 23774 4116 23826
rect 3948 23772 4116 23774
rect 5180 23828 5236 24670
rect 7868 23940 7924 25228
rect 8016 25116 8280 25126
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8016 25050 8280 25060
rect 7868 23874 7924 23884
rect 9324 23938 9380 25228
rect 9324 23886 9326 23938
rect 9378 23886 9380 23938
rect 9324 23874 9380 23886
rect 3948 23762 4004 23772
rect 5180 23762 5236 23772
rect 6076 23826 6132 23838
rect 6076 23774 6078 23826
rect 6130 23774 6132 23826
rect 2044 23378 2212 23380
rect 2044 23326 2046 23378
rect 2098 23326 2212 23378
rect 2044 23324 2212 23326
rect 2940 23716 2996 23726
rect 2044 23314 2100 23324
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 22932 1764 23102
rect 1708 22866 1764 22876
rect 2492 23042 2548 23054
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22932 2548 22990
rect 2492 22866 2548 22876
rect 2940 22370 2996 23660
rect 4732 23716 4788 23726
rect 4732 23622 4788 23660
rect 5740 23714 5796 23726
rect 5740 23662 5742 23714
rect 5794 23662 5796 23714
rect 4614 22764 4878 22774
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4614 22698 4878 22708
rect 2940 22318 2942 22370
rect 2994 22318 2996 22370
rect 2940 22306 2996 22318
rect 2268 22260 2324 22270
rect 2156 22146 2212 22158
rect 2156 22094 2158 22146
rect 2210 22094 2212 22146
rect 2156 21588 2212 22094
rect 2156 21522 2212 21532
rect 2268 21474 2324 22204
rect 2940 21812 2996 21822
rect 2940 21718 2996 21756
rect 5740 21812 5796 23662
rect 5740 21746 5796 21756
rect 2268 21422 2270 21474
rect 2322 21422 2324 21474
rect 2268 21410 2324 21422
rect 4614 21196 4878 21206
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4614 21130 4878 21140
rect 2380 20916 2436 20926
rect 1820 20802 1876 20814
rect 1820 20750 1822 20802
rect 1874 20750 1876 20802
rect 1820 20244 1876 20750
rect 2044 20692 2100 20702
rect 2044 20598 2100 20636
rect 2380 20690 2436 20860
rect 2380 20638 2382 20690
rect 2434 20638 2436 20690
rect 2380 20626 2436 20638
rect 6076 20692 6132 23774
rect 9660 23828 9716 23838
rect 9772 23828 9828 26238
rect 9996 24948 10052 27020
rect 10108 26850 10164 29200
rect 10780 26908 10836 29200
rect 10108 26798 10110 26850
rect 10162 26798 10164 26850
rect 10108 26786 10164 26798
rect 10668 26852 10836 26908
rect 10108 26404 10164 26414
rect 10164 26348 10276 26404
rect 10108 26338 10164 26348
rect 10108 24948 10164 24958
rect 9996 24946 10164 24948
rect 9996 24894 10110 24946
rect 10162 24894 10164 24946
rect 9996 24892 10164 24894
rect 10108 24882 10164 24892
rect 10108 23940 10164 23950
rect 10220 23940 10276 26348
rect 10668 26402 10724 26852
rect 10668 26350 10670 26402
rect 10722 26350 10724 26402
rect 10668 26338 10724 26350
rect 11116 26850 11172 26862
rect 11116 26798 11118 26850
rect 11170 26798 11172 26850
rect 11116 25618 11172 26798
rect 11340 26292 11396 26302
rect 11116 25566 11118 25618
rect 11170 25566 11172 25618
rect 11116 25554 11172 25566
rect 11228 26290 11396 26292
rect 11228 26238 11342 26290
rect 11394 26238 11396 26290
rect 11228 26236 11396 26238
rect 10668 25508 10724 25518
rect 10108 23938 10276 23940
rect 10108 23886 10110 23938
rect 10162 23886 10276 23938
rect 10108 23884 10276 23886
rect 10332 25284 10388 25294
rect 10108 23874 10164 23884
rect 9660 23826 9828 23828
rect 9660 23774 9662 23826
rect 9714 23774 9828 23826
rect 9660 23772 9828 23774
rect 10332 23826 10388 25228
rect 10332 23774 10334 23826
rect 10386 23774 10388 23826
rect 9660 23762 9716 23772
rect 10332 23762 10388 23774
rect 10556 25282 10612 25294
rect 10556 25230 10558 25282
rect 10610 25230 10612 25282
rect 8016 23548 8280 23558
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8016 23482 8280 23492
rect 10556 23378 10612 25230
rect 10668 23938 10724 25452
rect 10668 23886 10670 23938
rect 10722 23886 10724 23938
rect 10668 23874 10724 23886
rect 10780 25396 10836 25406
rect 10556 23326 10558 23378
rect 10610 23326 10612 23378
rect 10556 23314 10612 23326
rect 10780 23154 10836 25340
rect 11228 24948 11284 26236
rect 11340 26226 11396 26236
rect 11452 26068 11508 29200
rect 12124 26908 12180 29200
rect 12124 26852 12292 26908
rect 12236 26402 12292 26852
rect 12796 26516 12852 29200
rect 13468 26908 13524 29200
rect 14140 26908 14196 29200
rect 13468 26852 13748 26908
rect 14140 26852 14420 26908
rect 12796 26450 12852 26460
rect 13580 26516 13636 26526
rect 12236 26350 12238 26402
rect 12290 26350 12292 26402
rect 12236 26338 12292 26350
rect 13132 26292 13188 26302
rect 12348 26290 13188 26292
rect 12348 26238 13134 26290
rect 13186 26238 13188 26290
rect 12348 26236 13188 26238
rect 11452 26002 11508 26012
rect 12124 26068 12180 26078
rect 11418 25900 11682 25910
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11418 25834 11682 25844
rect 11004 24892 11284 24948
rect 11452 25620 11508 25630
rect 10892 24722 10948 24734
rect 10892 24670 10894 24722
rect 10946 24670 10948 24722
rect 10892 23492 10948 24670
rect 11004 23826 11060 24892
rect 11452 24500 11508 25564
rect 12124 25618 12180 26012
rect 12124 25566 12126 25618
rect 12178 25566 12180 25618
rect 12124 25554 12180 25566
rect 11676 25284 11732 25294
rect 11676 25190 11732 25228
rect 12124 25284 12180 25294
rect 11228 24444 11508 24500
rect 11228 24164 11284 24444
rect 11418 24332 11682 24342
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11418 24266 11682 24276
rect 11228 24108 11508 24164
rect 11340 23940 11396 23950
rect 11340 23846 11396 23884
rect 11004 23774 11006 23826
rect 11058 23774 11060 23826
rect 11004 23762 11060 23774
rect 10892 23436 11060 23492
rect 11004 23380 11060 23436
rect 11228 23380 11284 23390
rect 11004 23378 11284 23380
rect 11004 23326 11230 23378
rect 11282 23326 11284 23378
rect 11004 23324 11284 23326
rect 11228 23314 11284 23324
rect 10780 23102 10782 23154
rect 10834 23102 10836 23154
rect 10780 23090 10836 23102
rect 11452 23154 11508 24108
rect 12124 23938 12180 25228
rect 12124 23886 12126 23938
rect 12178 23886 12180 23938
rect 12124 23874 12180 23886
rect 11676 23828 11732 23838
rect 11676 23734 11732 23772
rect 12348 23826 12404 26236
rect 13132 26226 13188 26236
rect 13580 26178 13636 26460
rect 13580 26126 13582 26178
rect 13634 26126 13636 26178
rect 13580 26114 13636 26126
rect 13692 25394 13748 26852
rect 13692 25342 13694 25394
rect 13746 25342 13748 25394
rect 13692 25330 13748 25342
rect 14364 25394 14420 26852
rect 14812 26852 14868 29200
rect 14812 26786 14868 26796
rect 14820 26684 15084 26694
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 14820 26618 15084 26628
rect 15036 26292 15092 26302
rect 15036 26290 15316 26292
rect 15036 26238 15038 26290
rect 15090 26238 15316 26290
rect 15036 26236 15316 26238
rect 15036 26226 15092 26236
rect 15036 25730 15092 25742
rect 15036 25678 15038 25730
rect 15090 25678 15092 25730
rect 15036 25618 15092 25678
rect 15036 25566 15038 25618
rect 15090 25566 15092 25618
rect 15036 25554 15092 25566
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 14364 25330 14420 25342
rect 14820 25116 15084 25126
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 14820 25050 15084 25060
rect 12348 23774 12350 23826
rect 12402 23774 12404 23826
rect 12348 23762 12404 23774
rect 15260 23828 15316 26236
rect 15484 25844 15540 29200
rect 15820 26852 15876 26862
rect 15820 26514 15876 26796
rect 15820 26462 15822 26514
rect 15874 26462 15876 26514
rect 15820 26450 15876 26462
rect 15372 25788 15540 25844
rect 15372 25730 15428 25788
rect 16156 25732 16212 29200
rect 16828 26850 16884 29200
rect 16828 26798 16830 26850
rect 16882 26798 16884 26850
rect 16828 26786 16884 26798
rect 15372 25678 15374 25730
rect 15426 25678 15428 25730
rect 15372 25508 15428 25678
rect 15484 25676 16212 25732
rect 15484 25618 15540 25676
rect 15484 25566 15486 25618
rect 15538 25566 15540 25618
rect 15484 25554 15540 25566
rect 15372 25442 15428 25452
rect 15932 25508 15988 25518
rect 16156 25508 16212 25676
rect 17500 26516 17556 29200
rect 18172 26516 18228 29200
rect 17500 26460 17780 26516
rect 17500 25618 17556 26460
rect 17500 25566 17502 25618
rect 17554 25566 17556 25618
rect 17500 25554 17556 25566
rect 17612 26290 17668 26302
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 16380 25508 16436 25518
rect 16156 25506 16436 25508
rect 16156 25454 16382 25506
rect 16434 25454 16436 25506
rect 16156 25452 16436 25454
rect 15932 25414 15988 25452
rect 16380 25442 16436 25452
rect 15708 25284 15764 25294
rect 15708 25190 15764 25228
rect 16716 25284 16772 25294
rect 16716 25282 17220 25284
rect 16716 25230 16718 25282
rect 16770 25230 17220 25282
rect 16716 25228 17220 25230
rect 16716 25218 16772 25228
rect 17164 23938 17220 25228
rect 17164 23886 17166 23938
rect 17218 23886 17220 23938
rect 17164 23874 17220 23886
rect 15260 23762 15316 23772
rect 17500 23828 17556 23838
rect 17612 23828 17668 26238
rect 17724 25506 17780 26460
rect 18172 26450 18228 26460
rect 18284 26850 18340 26862
rect 18284 26798 18286 26850
rect 18338 26798 18340 26850
rect 18284 26514 18340 26798
rect 18284 26462 18286 26514
rect 18338 26462 18340 26514
rect 18284 26450 18340 26462
rect 18620 26290 18676 26302
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18222 25900 18486 25910
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18222 25834 18486 25844
rect 17724 25454 17726 25506
rect 17778 25454 17780 25506
rect 17724 25442 17780 25454
rect 18060 25284 18116 25294
rect 18620 25284 18676 26238
rect 18844 25620 18900 29200
rect 19516 29148 19796 29200
rect 19964 26852 20020 29260
rect 20160 29200 20272 30000
rect 20832 29200 20944 30000
rect 21504 29200 21616 30000
rect 22176 29200 22288 30000
rect 22848 29200 22960 30000
rect 23520 29200 23632 30000
rect 24192 29200 24304 30000
rect 20188 27076 20244 29200
rect 20188 27020 20468 27076
rect 19964 26796 20356 26852
rect 19068 26516 19124 26526
rect 19068 26178 19124 26460
rect 20300 26514 20356 26796
rect 20300 26462 20302 26514
rect 20354 26462 20356 26514
rect 20300 26292 20356 26462
rect 20300 26226 20356 26236
rect 20412 26404 20468 27020
rect 20748 26404 20804 26414
rect 19068 26126 19070 26178
rect 19122 26126 19124 26178
rect 19068 26114 19124 26126
rect 18844 25618 19124 25620
rect 18844 25566 18846 25618
rect 18898 25566 19124 25618
rect 18844 25564 19124 25566
rect 18844 25554 18900 25564
rect 19068 25506 19124 25564
rect 20412 25618 20468 26348
rect 20412 25566 20414 25618
rect 20466 25566 20468 25618
rect 20412 25554 20468 25566
rect 20524 26402 20804 26404
rect 20524 26350 20750 26402
rect 20802 26350 20804 26402
rect 20524 26348 20804 26350
rect 19068 25454 19070 25506
rect 19122 25454 19124 25506
rect 19068 25442 19124 25454
rect 17948 25282 18116 25284
rect 17948 25230 18062 25282
rect 18114 25230 18116 25282
rect 17948 25228 18116 25230
rect 17948 23938 18004 25228
rect 18060 25218 18116 25228
rect 18284 25228 18676 25284
rect 19404 25284 19460 25294
rect 18284 24500 18340 25228
rect 19404 25190 19460 25228
rect 17948 23886 17950 23938
rect 18002 23886 18004 23938
rect 17948 23874 18004 23886
rect 18060 24444 18340 24500
rect 17500 23826 17668 23828
rect 17500 23774 17502 23826
rect 17554 23774 17668 23826
rect 17500 23772 17668 23774
rect 18060 23828 18116 24444
rect 18222 24332 18486 24342
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18222 24266 18486 24276
rect 20524 23938 20580 26348
rect 20748 26338 20804 26348
rect 20860 25618 20916 29200
rect 21532 26852 21588 29200
rect 21532 26796 22036 26852
rect 21624 26684 21888 26694
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21624 26618 21888 26628
rect 21420 26402 21476 26414
rect 21420 26350 21422 26402
rect 21474 26350 21476 26402
rect 20972 26292 21028 26302
rect 20972 26198 21028 26236
rect 20860 25566 20862 25618
rect 20914 25566 20916 25618
rect 20860 25508 20916 25566
rect 20860 25442 20916 25452
rect 20748 25396 20804 25406
rect 20524 23886 20526 23938
rect 20578 23886 20580 23938
rect 20524 23874 20580 23886
rect 20636 25284 20692 25294
rect 18172 23828 18228 23838
rect 18060 23826 18228 23828
rect 18060 23774 18174 23826
rect 18226 23774 18228 23826
rect 18060 23772 18228 23774
rect 17500 23762 17556 23772
rect 18172 23762 18228 23772
rect 14820 23548 15084 23558
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 14820 23482 15084 23492
rect 20636 23266 20692 25228
rect 20748 23826 20804 25340
rect 21308 25284 21364 25294
rect 20972 25282 21364 25284
rect 20972 25230 21310 25282
rect 21362 25230 21364 25282
rect 20972 25228 21364 25230
rect 20972 24722 21028 25228
rect 21308 25218 21364 25228
rect 21196 25060 21252 25070
rect 21196 24946 21252 25004
rect 21196 24894 21198 24946
rect 21250 24894 21252 24946
rect 21196 24882 21252 24894
rect 20972 24670 20974 24722
rect 21026 24670 21028 24722
rect 20972 24658 21028 24670
rect 20748 23774 20750 23826
rect 20802 23774 20804 23826
rect 20748 23762 20804 23774
rect 20972 24500 21028 24510
rect 20972 23378 21028 24444
rect 21420 23938 21476 26350
rect 21532 26404 21588 26414
rect 21588 26348 21700 26404
rect 21532 26338 21588 26348
rect 21644 26290 21700 26348
rect 21644 26238 21646 26290
rect 21698 26238 21700 26290
rect 21644 26226 21700 26238
rect 21644 25508 21700 25518
rect 21644 25414 21700 25452
rect 21980 25394 22036 26796
rect 22204 26850 22260 29200
rect 22204 26798 22206 26850
rect 22258 26798 22260 26850
rect 22204 26786 22260 26798
rect 21980 25342 21982 25394
rect 22034 25342 22036 25394
rect 21980 25330 22036 25342
rect 22428 26290 22484 26302
rect 22428 26238 22430 26290
rect 22482 26238 22484 26290
rect 21624 25116 21888 25126
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21624 25050 21888 25060
rect 22428 24500 22484 26238
rect 22876 25732 22932 29200
rect 23212 26850 23268 26862
rect 23212 26798 23214 26850
rect 23266 26798 23268 26850
rect 23212 26514 23268 26798
rect 23548 26850 23604 29200
rect 23548 26798 23550 26850
rect 23602 26798 23604 26850
rect 23548 26786 23604 26798
rect 23212 26462 23214 26514
rect 23266 26462 23268 26514
rect 23212 26450 23268 26462
rect 22876 25666 22932 25676
rect 23548 25732 23604 25742
rect 23548 25618 23604 25676
rect 24220 25732 24276 29200
rect 24220 25666 24276 25676
rect 24444 28980 24500 28990
rect 23548 25566 23550 25618
rect 23602 25566 23604 25618
rect 23548 25554 23604 25566
rect 23100 25396 23156 25406
rect 23100 25302 23156 25340
rect 24108 24948 24164 24958
rect 24444 24948 24500 28924
rect 27804 28308 27860 28318
rect 26124 26964 26180 26974
rect 25004 26850 25060 26862
rect 25004 26798 25006 26850
rect 25058 26798 25060 26850
rect 24108 24946 24500 24948
rect 24108 24894 24110 24946
rect 24162 24894 24500 24946
rect 24108 24892 24500 24894
rect 24108 24882 24164 24892
rect 24444 24722 24500 24892
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24444 24658 24500 24670
rect 24556 26290 24612 26302
rect 24556 26238 24558 26290
rect 24610 26238 24612 26290
rect 22428 24434 22484 24444
rect 24332 24500 24388 24510
rect 21420 23886 21422 23938
rect 21474 23886 21476 23938
rect 21420 23874 21476 23886
rect 24108 23938 24164 23950
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 21644 23828 21700 23838
rect 21644 23734 21700 23772
rect 21624 23548 21888 23558
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21624 23482 21888 23492
rect 20972 23326 20974 23378
rect 21026 23326 21028 23378
rect 20972 23314 21028 23326
rect 20636 23214 20638 23266
rect 20690 23214 20692 23266
rect 20636 23202 20692 23214
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11452 23090 11508 23102
rect 24108 23156 24164 23886
rect 24332 23826 24388 24444
rect 24332 23774 24334 23826
rect 24386 23774 24388 23826
rect 24332 23762 24388 23774
rect 24556 23828 24612 26238
rect 25004 26178 25060 26798
rect 25004 26126 25006 26178
rect 25058 26126 25060 26178
rect 25004 26114 25060 26126
rect 25026 25900 25290 25910
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25026 25834 25290 25844
rect 25340 25732 25396 25742
rect 25340 25618 25396 25676
rect 25340 25566 25342 25618
rect 25394 25566 25396 25618
rect 25340 25554 25396 25566
rect 24668 25284 24724 25294
rect 24668 25190 24724 25228
rect 26124 24946 26180 26908
rect 26572 26292 26628 26302
rect 26348 26290 26628 26292
rect 26348 26238 26574 26290
rect 26626 26238 26628 26290
rect 26348 26236 26628 26238
rect 26124 24894 26126 24946
rect 26178 24894 26180 24946
rect 26124 24882 26180 24894
rect 26236 25394 26292 25406
rect 26236 25342 26238 25394
rect 26290 25342 26292 25394
rect 24556 23762 24612 23772
rect 24668 24834 24724 24846
rect 24668 24782 24670 24834
rect 24722 24782 24724 24834
rect 24668 23268 24724 24782
rect 25340 24722 25396 24734
rect 25340 24670 25342 24722
rect 25394 24670 25396 24722
rect 25340 24500 25396 24670
rect 25340 24434 25396 24444
rect 25788 24724 25844 24734
rect 25026 24332 25290 24342
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25026 24266 25290 24276
rect 24668 23202 24724 23212
rect 24780 23826 24836 23838
rect 24780 23774 24782 23826
rect 24834 23774 24836 23826
rect 24108 23090 24164 23100
rect 11418 22764 11682 22774
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11418 22698 11682 22708
rect 18222 22764 18486 22774
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18222 22698 18486 22708
rect 8016 21980 8280 21990
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8016 21914 8280 21924
rect 14820 21980 15084 21990
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 14820 21914 15084 21924
rect 21624 21980 21888 21990
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21624 21914 21888 21924
rect 20636 21700 20692 21710
rect 11418 21196 11682 21206
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11418 21130 11682 21140
rect 18222 21196 18486 21206
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18222 21130 18486 21140
rect 6076 20626 6132 20636
rect 12124 20916 12180 20926
rect 8016 20412 8280 20422
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8016 20346 8280 20356
rect 1820 20178 1876 20188
rect 11452 20020 11508 20030
rect 11228 20018 11508 20020
rect 11228 19966 11454 20018
rect 11506 19966 11508 20018
rect 11228 19964 11508 19966
rect 4614 19628 4878 19638
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4614 19562 4878 19572
rect 7756 19348 7812 19358
rect 6300 18564 6356 18574
rect 4956 18450 5012 18462
rect 4956 18398 4958 18450
rect 5010 18398 5012 18450
rect 4614 18060 4878 18070
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4614 17994 4878 18004
rect 4732 17666 4788 17678
rect 4732 17614 4734 17666
rect 4786 17614 4788 17666
rect 4732 16996 4788 17614
rect 4844 17556 4900 17566
rect 4844 17462 4900 17500
rect 4844 16996 4900 17006
rect 4732 16940 4844 16996
rect 4844 16930 4900 16940
rect 3164 16884 3220 16894
rect 3164 16790 3220 16828
rect 3612 16882 3668 16894
rect 3612 16830 3614 16882
rect 3666 16830 3668 16882
rect 3612 16212 3668 16830
rect 4956 16884 5012 18398
rect 5404 18452 5460 18462
rect 5404 18450 5572 18452
rect 5404 18398 5406 18450
rect 5458 18398 5572 18450
rect 5404 18396 5572 18398
rect 5404 18386 5460 18396
rect 4956 16818 5012 16828
rect 5404 16884 5460 16894
rect 4614 16492 4878 16502
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4614 16426 4878 16436
rect 3836 16212 3892 16222
rect 3612 16210 3892 16212
rect 3612 16158 3838 16210
rect 3890 16158 3892 16210
rect 3612 16156 3892 16158
rect 3836 16146 3892 16156
rect 4956 16212 5012 16222
rect 2716 15988 2772 15998
rect 1932 15986 2772 15988
rect 1932 15934 2718 15986
rect 2770 15934 2772 15986
rect 1932 15932 2772 15934
rect 1932 15538 1988 15932
rect 2716 15922 2772 15932
rect 1932 15486 1934 15538
rect 1986 15486 1988 15538
rect 1932 15474 1988 15486
rect 2716 15426 2772 15438
rect 2716 15374 2718 15426
rect 2770 15374 2772 15426
rect 2716 14756 2772 15374
rect 4956 15314 5012 16156
rect 4956 15262 4958 15314
rect 5010 15262 5012 15314
rect 4956 15250 5012 15262
rect 5404 15314 5460 16828
rect 5516 16212 5572 18396
rect 6300 17890 6356 18508
rect 7644 18564 7700 18574
rect 7644 18470 7700 18508
rect 6300 17838 6302 17890
rect 6354 17838 6356 17890
rect 6300 17826 6356 17838
rect 6860 17666 6916 17678
rect 6860 17614 6862 17666
rect 6914 17614 6916 17666
rect 5852 17556 5908 17566
rect 5852 17106 5908 17500
rect 5852 17054 5854 17106
rect 5906 17054 5908 17106
rect 5852 17042 5908 17054
rect 6860 16996 6916 17614
rect 6860 16930 6916 16940
rect 7084 17668 7140 17678
rect 7084 16884 7140 17612
rect 7756 17666 7812 19292
rect 8652 19348 8708 19358
rect 10444 19348 10500 19358
rect 8652 19254 8708 19292
rect 10108 19292 10444 19348
rect 9660 19124 9716 19134
rect 8428 19122 9716 19124
rect 8428 19070 9662 19122
rect 9714 19070 9716 19122
rect 8428 19068 9716 19070
rect 8016 18844 8280 18854
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8016 18778 8280 18788
rect 8428 18674 8484 19068
rect 9660 19058 9716 19068
rect 8428 18622 8430 18674
rect 8482 18622 8484 18674
rect 8428 18610 8484 18622
rect 7756 17614 7758 17666
rect 7810 17614 7812 17666
rect 7756 17602 7812 17614
rect 9436 18452 9492 18462
rect 9436 17668 9492 18396
rect 10108 18450 10164 19292
rect 10444 19282 10500 19292
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18386 10164 18398
rect 10780 19124 10836 19134
rect 10780 17890 10836 19068
rect 11228 18452 11284 19964
rect 11452 19954 11508 19964
rect 12124 20018 12180 20860
rect 14476 20916 14532 20926
rect 14476 20822 14532 20860
rect 19068 20802 19124 20814
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 15484 20690 15540 20702
rect 15484 20638 15486 20690
rect 15538 20638 15540 20690
rect 14820 20412 15084 20422
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 14820 20346 15084 20356
rect 14364 20132 14420 20142
rect 12124 19966 12126 20018
rect 12178 19966 12180 20018
rect 12124 19954 12180 19966
rect 14140 20130 14420 20132
rect 14140 20078 14366 20130
rect 14418 20078 14420 20130
rect 14140 20076 14420 20078
rect 11418 19628 11682 19638
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11418 19562 11682 19572
rect 11452 19348 11508 19358
rect 11452 19254 11508 19292
rect 13916 19348 13972 19358
rect 12460 19124 12516 19134
rect 12460 19030 12516 19068
rect 11228 18386 11284 18396
rect 12572 18674 12628 18686
rect 12572 18622 12574 18674
rect 12626 18622 12628 18674
rect 11418 18060 11682 18070
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11418 17994 11682 18004
rect 10780 17838 10782 17890
rect 10834 17838 10836 17890
rect 10780 17826 10836 17838
rect 12572 17890 12628 18622
rect 13244 18452 13300 18462
rect 13244 18358 13300 18396
rect 13916 18450 13972 19292
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13916 18386 13972 18398
rect 13132 18340 13188 18350
rect 13132 18246 13188 18284
rect 12572 17838 12574 17890
rect 12626 17838 12628 17890
rect 12572 17826 12628 17838
rect 14140 17890 14196 20076
rect 14364 20066 14420 20076
rect 15148 19794 15204 19806
rect 15148 19742 15150 19794
rect 15202 19742 15204 19794
rect 15148 19684 15204 19742
rect 15372 19684 15428 19694
rect 15148 19628 15372 19684
rect 15372 19618 15428 19628
rect 15260 19348 15316 19358
rect 15260 19254 15316 19292
rect 14140 17838 14142 17890
rect 14194 17838 14196 17890
rect 14140 17826 14196 17838
rect 14252 19012 14308 19022
rect 9492 17612 9828 17668
rect 9436 17602 9492 17612
rect 8016 17276 8280 17286
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8016 17210 8280 17220
rect 9772 16996 9828 17612
rect 12684 17666 12740 17678
rect 12684 17614 12686 17666
rect 12738 17614 12740 17666
rect 9996 17444 10052 17454
rect 9660 16994 9828 16996
rect 9660 16942 9774 16994
rect 9826 16942 9828 16994
rect 9660 16940 9828 16942
rect 7084 16818 7140 16828
rect 7532 16884 7588 16894
rect 7532 16790 7588 16828
rect 6300 16660 6356 16670
rect 6188 16212 6244 16222
rect 5516 16210 6244 16212
rect 5516 16158 6190 16210
rect 6242 16158 6244 16210
rect 5516 16156 6244 16158
rect 6188 16146 6244 16156
rect 5404 15262 5406 15314
rect 5458 15262 5460 15314
rect 5404 15250 5460 15262
rect 5516 15428 5572 15438
rect 5516 15148 5572 15372
rect 5404 15092 5572 15148
rect 4614 14924 4878 14934
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4614 14858 4878 14868
rect 2716 14690 2772 14700
rect 3948 14756 4004 14766
rect 3948 14662 4004 14700
rect 4172 14530 4228 14542
rect 4172 14478 4174 14530
rect 4226 14478 4228 14530
rect 3500 14420 3556 14430
rect 2380 13858 2436 13870
rect 2380 13806 2382 13858
rect 2434 13806 2436 13858
rect 1596 13522 1652 13534
rect 1596 13470 1598 13522
rect 1650 13470 1652 13522
rect 1596 12404 1652 13470
rect 2380 13188 2436 13806
rect 2380 13122 2436 13132
rect 3276 13188 3332 13198
rect 3276 13094 3332 13132
rect 2380 12964 2436 12974
rect 1596 12338 1652 12348
rect 1708 12850 1764 12862
rect 1708 12798 1710 12850
rect 1762 12798 1764 12850
rect 1708 12740 1764 12798
rect 1708 12180 1764 12684
rect 1708 12114 1764 12124
rect 2044 12738 2100 12750
rect 2044 12686 2046 12738
rect 2098 12686 2100 12738
rect 2044 12178 2100 12686
rect 2044 12126 2046 12178
rect 2098 12126 2100 12178
rect 2044 12114 2100 12126
rect 2044 10722 2100 10734
rect 2044 10670 2046 10722
rect 2098 10670 2100 10722
rect 1820 10610 1876 10622
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 10164 1876 10558
rect 2044 10388 2100 10670
rect 2380 10612 2436 12908
rect 3388 12962 3444 12974
rect 3388 12910 3390 12962
rect 3442 12910 3444 12962
rect 3388 12852 3444 12910
rect 2492 12740 2548 12750
rect 2492 12646 2548 12684
rect 2604 12404 2660 12414
rect 2044 10322 2100 10332
rect 2268 10610 2436 10612
rect 2268 10558 2382 10610
rect 2434 10558 2436 10610
rect 2268 10556 2436 10558
rect 1820 9938 1876 10108
rect 1820 9886 1822 9938
rect 1874 9886 1876 9938
rect 1820 9874 1876 9886
rect 2044 9044 2100 9054
rect 2268 9044 2324 10556
rect 2380 10546 2436 10556
rect 2492 12178 2548 12190
rect 2492 12126 2494 12178
rect 2546 12126 2548 12178
rect 2044 9042 2324 9044
rect 2044 8990 2046 9042
rect 2098 8990 2324 9042
rect 2044 8988 2324 8990
rect 2492 9042 2548 12126
rect 2604 11282 2660 12348
rect 3276 12180 3332 12190
rect 3388 12180 3444 12796
rect 3500 12402 3556 14364
rect 4172 12852 4228 14478
rect 5404 13970 5460 15092
rect 5404 13918 5406 13970
rect 5458 13918 5460 13970
rect 5404 13906 5460 13918
rect 6188 13972 6244 13982
rect 6300 13972 6356 16604
rect 6636 16658 6692 16670
rect 6636 16606 6638 16658
rect 6690 16606 6692 16658
rect 6636 15988 6692 16606
rect 7308 16660 7364 16670
rect 7308 16566 7364 16604
rect 6636 15922 6692 15932
rect 7308 15988 7364 15998
rect 7308 15894 7364 15932
rect 8016 15708 8280 15718
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8016 15642 8280 15652
rect 7980 15428 8036 15438
rect 7980 15334 8036 15372
rect 6972 15202 7028 15214
rect 6972 15150 6974 15202
rect 7026 15150 7028 15202
rect 6748 14420 6804 14430
rect 6748 14326 6804 14364
rect 6188 13970 6356 13972
rect 6188 13918 6190 13970
rect 6242 13918 6356 13970
rect 6188 13916 6356 13918
rect 6188 13906 6244 13916
rect 4732 13746 4788 13758
rect 4732 13694 4734 13746
rect 4786 13694 4788 13746
rect 4732 13524 4788 13694
rect 4732 13458 4788 13468
rect 5180 13746 5236 13758
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 4614 13356 4878 13366
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4614 13290 4878 13300
rect 4172 12786 4228 12796
rect 4620 12962 4676 12974
rect 4620 12910 4622 12962
rect 4674 12910 4676 12962
rect 4620 12852 4676 12910
rect 5180 12964 5236 13694
rect 6524 13524 6580 13534
rect 6188 13412 6244 13422
rect 5180 12898 5236 12908
rect 5516 12964 5572 12974
rect 5516 12870 5572 12908
rect 6188 12962 6244 13356
rect 6188 12910 6190 12962
rect 6242 12910 6244 12962
rect 6188 12898 6244 12910
rect 4396 12738 4452 12750
rect 4396 12686 4398 12738
rect 4450 12686 4452 12738
rect 3500 12350 3502 12402
rect 3554 12350 3556 12402
rect 3500 12338 3556 12350
rect 4284 12404 4340 12414
rect 4396 12404 4452 12686
rect 4284 12402 4452 12404
rect 4284 12350 4286 12402
rect 4338 12350 4452 12402
rect 4284 12348 4452 12350
rect 4284 12338 4340 12348
rect 3276 12178 3444 12180
rect 3276 12126 3278 12178
rect 3330 12126 3444 12178
rect 3276 12124 3444 12126
rect 3276 12114 3332 12124
rect 2604 11230 2606 11282
rect 2658 11230 2660 11282
rect 2604 11218 2660 11230
rect 3164 11954 3220 11966
rect 3164 11902 3166 11954
rect 3218 11902 3220 11954
rect 3164 11060 3220 11902
rect 4620 11956 4676 12796
rect 4620 11890 4676 11900
rect 4614 11788 4878 11798
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4614 11722 4878 11732
rect 5964 11732 6020 11742
rect 3164 10994 3220 11004
rect 3724 11506 3780 11518
rect 3724 11454 3726 11506
rect 3778 11454 3780 11506
rect 3052 10612 3108 10622
rect 3052 10518 3108 10556
rect 3724 10612 3780 11454
rect 5964 11394 6020 11676
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 11330 6020 11342
rect 5740 11172 5796 11182
rect 5516 11170 5796 11172
rect 5516 11118 5742 11170
rect 5794 11118 5796 11170
rect 5516 11116 5796 11118
rect 4844 11060 4900 11070
rect 4900 11004 5012 11060
rect 4844 10994 4900 11004
rect 3724 10546 3780 10556
rect 4614 10220 4878 10230
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4614 10154 4878 10164
rect 4956 9266 5012 11004
rect 5516 10834 5572 11116
rect 5740 11106 5796 11116
rect 5516 10782 5518 10834
rect 5570 10782 5572 10834
rect 5516 10770 5572 10782
rect 6076 10724 6132 10734
rect 6412 10724 6468 10734
rect 6076 10722 6468 10724
rect 6076 10670 6078 10722
rect 6130 10670 6414 10722
rect 6466 10670 6468 10722
rect 6076 10668 6468 10670
rect 6076 10658 6132 10668
rect 6412 10658 6468 10668
rect 6524 9940 6580 13468
rect 6972 13412 7028 15150
rect 8092 14642 8148 14654
rect 8092 14590 8094 14642
rect 8146 14590 8148 14642
rect 8092 14308 8148 14590
rect 9548 14532 9604 14542
rect 9660 14532 9716 16940
rect 9772 16930 9828 16940
rect 9884 17442 10052 17444
rect 9884 17390 9998 17442
rect 10050 17390 10052 17442
rect 9884 17388 10052 17390
rect 9884 15426 9940 17388
rect 9996 17378 10052 17388
rect 10220 16884 10276 16894
rect 9996 16212 10052 16222
rect 9996 16118 10052 16156
rect 9884 15374 9886 15426
rect 9938 15374 9940 15426
rect 9884 15362 9940 15374
rect 10220 15314 10276 16828
rect 11418 16492 11682 16502
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11418 16426 11682 16436
rect 12684 16100 12740 17614
rect 14140 17666 14196 17678
rect 14140 17614 14142 17666
rect 14194 17614 14196 17666
rect 13692 16772 13748 16782
rect 12908 16100 12964 16110
rect 12684 16044 12908 16100
rect 12908 16006 12964 16044
rect 13692 16100 13748 16716
rect 14140 16772 14196 17614
rect 14140 16706 14196 16716
rect 13692 16006 13748 16044
rect 11116 15986 11172 15998
rect 11116 15934 11118 15986
rect 11170 15934 11172 15986
rect 11116 15538 11172 15934
rect 11116 15486 11118 15538
rect 11170 15486 11172 15538
rect 11116 15474 11172 15486
rect 11900 15876 11956 15886
rect 11900 15538 11956 15820
rect 11900 15486 11902 15538
rect 11954 15486 11956 15538
rect 11900 15474 11956 15486
rect 12348 15874 12404 15886
rect 12348 15822 12350 15874
rect 12402 15822 12404 15874
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 9548 14530 9716 14532
rect 9548 14478 9550 14530
rect 9602 14478 9716 14530
rect 9548 14476 9716 14478
rect 9996 14530 10052 14542
rect 9996 14478 9998 14530
rect 10050 14478 10052 14530
rect 9548 14466 9604 14476
rect 8092 14252 8484 14308
rect 8016 14140 8280 14150
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8016 14074 8280 14084
rect 8428 13746 8484 14252
rect 9212 13860 9268 13870
rect 8428 13694 8430 13746
rect 8482 13694 8484 13746
rect 8428 13682 8484 13694
rect 8988 13746 9044 13758
rect 8988 13694 8990 13746
rect 9042 13694 9044 13746
rect 6972 13346 7028 13356
rect 6972 12964 7028 12974
rect 6636 12178 6692 12190
rect 6636 12126 6638 12178
rect 6690 12126 6692 12178
rect 6636 10500 6692 12126
rect 6972 12178 7028 12908
rect 6972 12126 6974 12178
rect 7026 12126 7028 12178
rect 6972 12114 7028 12126
rect 7868 12964 7924 12974
rect 6636 10434 6692 10444
rect 7532 10500 7588 10510
rect 7532 10406 7588 10444
rect 6636 9940 6692 9950
rect 6524 9938 6692 9940
rect 6524 9886 6638 9938
rect 6690 9886 6692 9938
rect 6524 9884 6692 9886
rect 6636 9874 6692 9884
rect 7868 9940 7924 12908
rect 8988 12964 9044 13694
rect 9212 13186 9268 13804
rect 9996 13636 10052 14478
rect 9996 13570 10052 13580
rect 9212 13134 9214 13186
rect 9266 13134 9268 13186
rect 9212 13122 9268 13134
rect 8652 12738 8708 12750
rect 8652 12686 8654 12738
rect 8706 12686 8708 12738
rect 8016 12572 8280 12582
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8016 12506 8280 12516
rect 8652 12290 8708 12686
rect 8652 12238 8654 12290
rect 8706 12238 8708 12290
rect 8652 12226 8708 12238
rect 8988 12292 9044 12908
rect 8988 12226 9044 12236
rect 9324 12738 9380 12750
rect 9324 12686 9326 12738
rect 9378 12686 9380 12738
rect 8540 12178 8596 12190
rect 8540 12126 8542 12178
rect 8594 12126 8596 12178
rect 8540 11732 8596 12126
rect 8540 11666 8596 11676
rect 9100 11732 9156 11742
rect 9100 11618 9156 11676
rect 9100 11566 9102 11618
rect 9154 11566 9156 11618
rect 9100 11554 9156 11566
rect 8016 11004 8280 11014
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8016 10938 8280 10948
rect 9324 10724 9380 12686
rect 10108 12738 10164 12750
rect 10108 12686 10110 12738
rect 10162 12686 10164 12738
rect 9772 12292 9828 12302
rect 9772 12198 9828 12236
rect 10108 10836 10164 12686
rect 10220 11732 10276 15262
rect 11418 14924 11682 14934
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11418 14858 11682 14868
rect 12348 14306 12404 15822
rect 13580 15876 13636 15886
rect 13580 15782 13636 15820
rect 14140 15314 14196 15326
rect 14140 15262 14142 15314
rect 14194 15262 14196 15314
rect 12348 14254 12350 14306
rect 12402 14254 12404 14306
rect 12348 14242 12404 14254
rect 13020 14308 13076 14318
rect 13020 14214 13076 14252
rect 13916 14308 13972 14318
rect 11788 13860 11844 13870
rect 11788 13766 11844 13804
rect 13916 13858 13972 14252
rect 13916 13806 13918 13858
rect 13970 13806 13972 13858
rect 13916 13794 13972 13806
rect 10780 13636 10836 13646
rect 14140 13636 14196 15262
rect 14252 14644 14308 18956
rect 14820 18844 15084 18854
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 14820 18778 15084 18788
rect 15484 18340 15540 20638
rect 16156 20020 16212 20030
rect 16156 20018 16436 20020
rect 16156 19966 16158 20018
rect 16210 19966 16436 20018
rect 16156 19964 16436 19966
rect 16156 19954 16212 19964
rect 15484 18274 15540 18284
rect 15932 19796 15988 19806
rect 14588 17668 14644 17678
rect 14588 15314 14644 17612
rect 15260 17668 15316 17678
rect 15260 17574 15316 17612
rect 15932 17666 15988 19740
rect 16044 19796 16100 19806
rect 16044 19794 16212 19796
rect 16044 19742 16046 19794
rect 16098 19742 16212 19794
rect 16044 19740 16212 19742
rect 16044 19730 16100 19740
rect 16156 18674 16212 19740
rect 16268 19684 16324 19694
rect 16268 19122 16324 19628
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 16268 19058 16324 19070
rect 16156 18622 16158 18674
rect 16210 18622 16212 18674
rect 16156 18610 16212 18622
rect 15932 17614 15934 17666
rect 15986 17614 15988 17666
rect 15932 17602 15988 17614
rect 16380 18340 16436 19964
rect 17612 19908 17668 19918
rect 17164 19234 17220 19246
rect 17164 19182 17166 19234
rect 17218 19182 17220 19234
rect 16940 18676 16996 18686
rect 16940 18450 16996 18620
rect 16940 18398 16942 18450
rect 16994 18398 16996 18450
rect 16940 18386 16996 18398
rect 17164 18452 17220 19182
rect 17612 19234 17668 19852
rect 18396 19906 18452 19918
rect 18396 19854 18398 19906
rect 18450 19854 18452 19906
rect 18396 19796 18452 19854
rect 18396 19730 18452 19740
rect 18222 19628 18486 19638
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18222 19562 18486 19572
rect 17612 19182 17614 19234
rect 17666 19182 17668 19234
rect 17612 19170 17668 19182
rect 18956 19012 19012 19022
rect 14820 17276 15084 17286
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 14820 17210 15084 17220
rect 14588 15262 14590 15314
rect 14642 15262 14644 15314
rect 14588 15250 14644 15262
rect 14700 16882 14756 16894
rect 14700 16830 14702 16882
rect 14754 16830 14756 16882
rect 14252 14642 14532 14644
rect 14252 14590 14254 14642
rect 14306 14590 14532 14642
rect 14252 14588 14532 14590
rect 14252 14578 14308 14588
rect 14476 14530 14532 14588
rect 14476 14478 14478 14530
rect 14530 14478 14532 14530
rect 14476 14466 14532 14478
rect 14252 13636 14308 13646
rect 14140 13580 14252 13636
rect 10780 13542 10836 13580
rect 14252 13570 14308 13580
rect 11418 13356 11682 13366
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11418 13290 11682 13300
rect 12460 12964 12516 12974
rect 12460 12870 12516 12908
rect 12796 12962 12852 12974
rect 12796 12910 12798 12962
rect 12850 12910 12852 12962
rect 11418 11788 11682 11798
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11418 11722 11682 11732
rect 10220 11666 10276 11676
rect 12684 11394 12740 11406
rect 12684 11342 12686 11394
rect 12738 11342 12740 11394
rect 10108 10770 10164 10780
rect 12348 10836 12404 10846
rect 9324 10658 9380 10668
rect 11788 10724 11844 10734
rect 11788 10630 11844 10668
rect 9996 10500 10052 10510
rect 7868 9874 7924 9884
rect 9772 10388 9828 10398
rect 9548 9828 9604 9838
rect 9548 9734 9604 9772
rect 4956 9214 4958 9266
rect 5010 9214 5012 9266
rect 4956 9202 5012 9214
rect 5516 9716 5572 9726
rect 5516 9266 5572 9660
rect 7644 9716 7700 9726
rect 7644 9622 7700 9660
rect 8016 9436 8280 9446
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8016 9370 8280 9380
rect 5516 9214 5518 9266
rect 5570 9214 5572 9266
rect 5516 9202 5572 9214
rect 2492 8990 2494 9042
rect 2546 8990 2548 9042
rect 2044 8978 2100 8988
rect 2492 8978 2548 8990
rect 9772 9042 9828 10332
rect 9996 9826 10052 10444
rect 10780 10500 10836 10510
rect 10780 10406 10836 10444
rect 11418 10220 11682 10230
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11418 10154 11682 10164
rect 9996 9774 9998 9826
rect 10050 9774 10052 9826
rect 9996 9762 10052 9774
rect 12348 9156 12404 10780
rect 12460 9716 12516 9726
rect 12460 9602 12516 9660
rect 12460 9550 12462 9602
rect 12514 9550 12516 9602
rect 12460 9538 12516 9550
rect 12460 9156 12516 9166
rect 12348 9154 12516 9156
rect 12348 9102 12462 9154
rect 12514 9102 12516 9154
rect 12348 9100 12516 9102
rect 12460 9090 12516 9100
rect 9772 8990 9774 9042
rect 9826 8990 9828 9042
rect 9772 8978 9828 8990
rect 12684 9042 12740 11342
rect 12796 10612 12852 12910
rect 14700 12180 14756 16830
rect 16380 16772 16436 18284
rect 17164 17668 17220 18396
rect 18172 18450 18228 18462
rect 18172 18398 18174 18450
rect 18226 18398 18228 18450
rect 18172 18340 18228 18398
rect 18732 18452 18788 18462
rect 18732 18358 18788 18396
rect 18172 18274 18228 18284
rect 17164 17602 17220 17612
rect 18060 18226 18116 18238
rect 18060 18174 18062 18226
rect 18114 18174 18116 18226
rect 18060 17556 18116 18174
rect 18222 18060 18486 18070
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18222 17994 18486 18004
rect 18956 17890 19012 18956
rect 19068 18340 19124 20750
rect 19292 20580 19348 20590
rect 19292 20578 19908 20580
rect 19292 20526 19294 20578
rect 19346 20526 19908 20578
rect 19292 20524 19908 20526
rect 19292 20514 19348 20524
rect 19292 20132 19348 20142
rect 19292 18450 19348 20076
rect 19404 20130 19460 20142
rect 19404 20078 19406 20130
rect 19458 20078 19460 20130
rect 19404 18676 19460 20078
rect 19852 19122 19908 20524
rect 20636 19458 20692 21644
rect 22204 21700 22260 21710
rect 22204 21606 22260 21644
rect 21196 21474 21252 21486
rect 21196 21422 21198 21474
rect 21250 21422 21252 21474
rect 21196 20132 21252 21422
rect 21624 20412 21888 20422
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21624 20346 21888 20356
rect 21196 20066 21252 20076
rect 22204 20130 22260 20142
rect 22204 20078 22206 20130
rect 22258 20078 22260 20130
rect 21196 19908 21252 19918
rect 21196 19814 21252 19852
rect 20636 19406 20638 19458
rect 20690 19406 20692 19458
rect 20636 19394 20692 19406
rect 19852 19070 19854 19122
rect 19906 19070 19908 19122
rect 19852 19058 19908 19070
rect 22204 19012 22260 20078
rect 22204 18946 22260 18956
rect 23212 19234 23268 19246
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 21624 18844 21888 18854
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21624 18778 21888 18788
rect 19404 18610 19460 18620
rect 20076 18564 20132 18574
rect 19292 18398 19294 18450
rect 19346 18398 19348 18450
rect 19292 18386 19348 18398
rect 19404 18452 19460 18462
rect 19068 18274 19124 18284
rect 18956 17838 18958 17890
rect 19010 17838 19012 17890
rect 18956 17826 19012 17838
rect 19404 17668 19460 18396
rect 18172 17556 18228 17566
rect 18060 17554 18228 17556
rect 18060 17502 18174 17554
rect 18226 17502 18228 17554
rect 18060 17500 18228 17502
rect 18172 17490 18228 17500
rect 15932 15876 15988 15886
rect 15932 15782 15988 15820
rect 14820 15708 15084 15718
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 14820 15642 15084 15652
rect 16380 15316 16436 16716
rect 18222 16492 18486 16502
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18222 16426 18486 16436
rect 19068 16098 19124 16110
rect 19068 16046 19070 16098
rect 19122 16046 19124 16098
rect 16716 15874 16772 15886
rect 16716 15822 16718 15874
rect 16770 15822 16772 15874
rect 16716 15538 16772 15822
rect 16716 15486 16718 15538
rect 16770 15486 16772 15538
rect 16716 15474 16772 15486
rect 17500 15876 17556 15886
rect 17500 15426 17556 15820
rect 17500 15374 17502 15426
rect 17554 15374 17556 15426
rect 17500 15362 17556 15374
rect 16492 15316 16548 15326
rect 16380 15314 16548 15316
rect 16380 15262 16494 15314
rect 16546 15262 16548 15314
rect 16380 15260 16548 15262
rect 14820 14140 15084 14150
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 14820 14074 15084 14084
rect 15036 13636 15092 13646
rect 15036 13542 15092 13580
rect 16380 13186 16436 15260
rect 16492 15250 16548 15260
rect 18620 15202 18676 15214
rect 18620 15150 18622 15202
rect 18674 15150 18676 15202
rect 18222 14924 18486 14934
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18222 14858 18486 14868
rect 18620 14756 18676 15150
rect 19068 15204 19124 16046
rect 19404 16098 19460 17612
rect 19628 18340 19684 18350
rect 19628 17668 19684 18284
rect 20076 17778 20132 18508
rect 21644 18564 21700 18574
rect 21644 18470 21700 18508
rect 22428 18452 22484 18462
rect 22428 18358 22484 18396
rect 20076 17726 20078 17778
rect 20130 17726 20132 17778
rect 20076 17714 20132 17726
rect 21868 18340 21924 18350
rect 21196 17668 21252 17678
rect 19628 17666 19908 17668
rect 19628 17614 19630 17666
rect 19682 17614 19908 17666
rect 19628 17612 19908 17614
rect 19628 17602 19684 17612
rect 19404 16046 19406 16098
rect 19458 16046 19460 16098
rect 19404 16034 19460 16046
rect 19516 16882 19572 16894
rect 19516 16830 19518 16882
rect 19570 16830 19572 16882
rect 19068 15138 19124 15148
rect 18284 14700 18676 14756
rect 16380 13134 16382 13186
rect 16434 13134 16436 13186
rect 16380 13122 16436 13134
rect 17612 13746 17668 13758
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 14820 12572 15084 12582
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 14820 12506 15084 12516
rect 14812 12180 14868 12190
rect 14700 12124 14812 12180
rect 14812 12086 14868 12124
rect 13916 11508 13972 11518
rect 13804 11452 13916 11508
rect 13244 10612 13300 10622
rect 12796 10610 12964 10612
rect 12796 10558 12798 10610
rect 12850 10558 12964 10610
rect 12796 10556 12964 10558
rect 12796 10546 12852 10556
rect 12684 8990 12686 9042
rect 12738 8990 12740 9042
rect 11900 8932 11956 8942
rect 11900 8838 11956 8876
rect 12684 8932 12740 8990
rect 12908 9828 12964 10556
rect 13244 10518 13300 10556
rect 12908 9044 12964 9772
rect 13020 9604 13076 9614
rect 13020 9602 13412 9604
rect 13020 9550 13022 9602
rect 13074 9550 13412 9602
rect 13020 9548 13412 9550
rect 13020 9538 13076 9548
rect 13244 9044 13300 9054
rect 12908 9042 13300 9044
rect 12908 8990 13246 9042
rect 13298 8990 13300 9042
rect 12908 8988 13300 8990
rect 13244 8978 13300 8988
rect 12684 8866 12740 8876
rect 4614 8652 4878 8662
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4614 8586 4878 8596
rect 11418 8652 11682 8662
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11418 8586 11682 8596
rect 2940 8258 2996 8270
rect 2940 8206 2942 8258
rect 2994 8206 2996 8258
rect 2044 8146 2100 8158
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 7476 2100 8094
rect 2940 7700 2996 8206
rect 3388 8258 3444 8270
rect 3388 8206 3390 8258
rect 3442 8206 3444 8258
rect 3388 8148 3444 8206
rect 3388 8082 3444 8092
rect 4060 8148 4116 8158
rect 4060 8054 4116 8092
rect 13356 8148 13412 9548
rect 13804 9042 13860 11452
rect 13916 11442 13972 11452
rect 16268 11508 16324 11546
rect 16268 11442 16324 11452
rect 16268 11284 16324 11294
rect 14820 11004 15084 11014
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 14820 10938 15084 10948
rect 16268 10834 16324 11228
rect 17276 11284 17332 11294
rect 17276 11190 17332 11228
rect 16268 10782 16270 10834
rect 16322 10782 16324 10834
rect 16268 10770 16324 10782
rect 15484 10724 15540 10734
rect 15036 10722 15540 10724
rect 15036 10670 15486 10722
rect 15538 10670 15540 10722
rect 15036 10668 15540 10670
rect 14476 10612 14532 10622
rect 14140 9828 14196 9838
rect 13916 9716 13972 9726
rect 13916 9622 13972 9660
rect 13804 8990 13806 9042
rect 13858 8990 13860 9042
rect 13804 8978 13860 8990
rect 14140 8932 14196 9772
rect 14140 8866 14196 8876
rect 14476 8370 14532 10556
rect 15036 9938 15092 10668
rect 15484 10658 15540 10668
rect 17276 10612 17332 10622
rect 17612 10612 17668 13694
rect 18284 13746 18340 14700
rect 18284 13694 18286 13746
rect 18338 13694 18340 13746
rect 18284 13682 18340 13694
rect 19516 14642 19572 16830
rect 19852 16098 19908 17612
rect 21252 17612 21476 17668
rect 21196 17574 21252 17612
rect 21420 16994 21476 17612
rect 21868 17666 21924 18284
rect 23100 18338 23156 18350
rect 23100 18286 23102 18338
rect 23154 18286 23156 18338
rect 23100 18228 23156 18286
rect 23100 18162 23156 18172
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17602 21924 17614
rect 23212 17668 23268 19182
rect 23884 19234 23940 19246
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 21624 17276 21888 17286
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21624 17210 21888 17220
rect 21420 16942 21422 16994
rect 21474 16942 21476 16994
rect 21420 16930 21476 16942
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19852 16034 19908 16046
rect 22764 16100 22820 16110
rect 20412 15876 20468 15886
rect 21196 15876 21252 15886
rect 20412 15874 20580 15876
rect 20412 15822 20414 15874
rect 20466 15822 20580 15874
rect 20412 15820 20580 15822
rect 20412 15810 20468 15820
rect 19516 14590 19518 14642
rect 19570 14590 19572 14642
rect 18222 13356 18486 13366
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18222 13290 18486 13300
rect 18732 12962 18788 12974
rect 18732 12910 18734 12962
rect 18786 12910 18788 12962
rect 18732 12066 18788 12910
rect 19516 12180 19572 14590
rect 20524 13970 20580 15820
rect 21196 15782 21252 15820
rect 21980 15874 22036 15886
rect 21980 15822 21982 15874
rect 22034 15822 22036 15874
rect 21624 15708 21888 15718
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21624 15642 21888 15652
rect 21308 15204 21364 15214
rect 21308 15110 21364 15148
rect 21980 15204 22036 15822
rect 22316 15876 22372 15886
rect 22316 15426 22372 15820
rect 22316 15374 22318 15426
rect 22370 15374 22372 15426
rect 22316 15362 22372 15374
rect 21980 15138 22036 15148
rect 22092 14530 22148 14542
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 20748 14308 20804 14318
rect 20860 14308 20916 14318
rect 20748 14306 20860 14308
rect 20748 14254 20750 14306
rect 20802 14254 20860 14306
rect 20748 14252 20860 14254
rect 20748 14242 20804 14252
rect 20524 13918 20526 13970
rect 20578 13918 20580 13970
rect 20524 13906 20580 13918
rect 19516 12086 19572 12124
rect 20748 12964 20804 12974
rect 18732 12014 18734 12066
rect 18786 12014 18788 12066
rect 18222 11788 18486 11798
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18222 11722 18486 11732
rect 17276 10610 17668 10612
rect 17276 10558 17278 10610
rect 17330 10558 17668 10610
rect 17276 10556 17668 10558
rect 17948 11508 18004 11518
rect 17948 10610 18004 11452
rect 17948 10558 17950 10610
rect 18002 10558 18004 10610
rect 16492 10500 16548 10510
rect 15036 9886 15038 9938
rect 15090 9886 15092 9938
rect 15036 9874 15092 9886
rect 16380 10498 16548 10500
rect 16380 10446 16494 10498
rect 16546 10446 16548 10498
rect 16380 10444 16548 10446
rect 14700 9828 14756 9838
rect 14700 9734 14756 9772
rect 15484 9828 15540 9838
rect 15484 9734 15540 9772
rect 15932 9826 15988 9838
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 14820 9436 15084 9446
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 14820 9370 15084 9380
rect 14476 8318 14478 8370
rect 14530 8318 14532 8370
rect 14476 8306 14532 8318
rect 15932 8372 15988 9774
rect 16380 9266 16436 10444
rect 16492 10434 16548 10444
rect 16828 10498 16884 10510
rect 16828 10446 16830 10498
rect 16882 10446 16884 10498
rect 16828 9940 16884 10446
rect 16828 9874 16884 9884
rect 17276 9828 17332 10556
rect 17948 10546 18004 10558
rect 18222 10220 18486 10230
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18222 10154 18486 10164
rect 17276 9762 17332 9772
rect 17948 9940 18004 9950
rect 16380 9214 16382 9266
rect 16434 9214 16436 9266
rect 16380 9202 16436 9214
rect 17948 9042 18004 9884
rect 18732 9940 18788 12014
rect 19068 12066 19124 12078
rect 19068 12014 19070 12066
rect 19122 12014 19124 12066
rect 18956 11284 19012 11294
rect 18956 10050 19012 11228
rect 19068 10836 19124 12014
rect 19292 11508 19348 11518
rect 19292 11414 19348 11452
rect 20300 11284 20356 11294
rect 20300 11190 20356 11228
rect 19068 10770 19124 10780
rect 20188 10836 20244 10846
rect 20188 10742 20244 10780
rect 18956 9998 18958 10050
rect 19010 9998 19012 10050
rect 18956 9986 19012 9998
rect 18732 9874 18788 9884
rect 19180 9940 19236 9950
rect 19180 9846 19236 9884
rect 19964 9828 20020 9838
rect 19964 9734 20020 9772
rect 18396 9604 18452 9614
rect 18396 9510 18452 9548
rect 19292 9604 19348 9614
rect 19292 9510 19348 9548
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 8978 18004 8990
rect 15932 8306 15988 8316
rect 16940 8818 16996 8830
rect 16940 8766 16942 8818
rect 16994 8766 16996 8818
rect 13356 8082 13412 8092
rect 15484 8148 15540 8158
rect 15484 8054 15540 8092
rect 16940 8148 16996 8766
rect 18222 8652 18486 8662
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18222 8586 18486 8596
rect 17612 8372 17668 8382
rect 17612 8278 17668 8316
rect 16940 8082 16996 8092
rect 18620 8148 18676 8158
rect 18620 8054 18676 8092
rect 3612 8036 3668 8046
rect 3612 8034 4004 8036
rect 3612 7982 3614 8034
rect 3666 7982 4004 8034
rect 3612 7980 4004 7982
rect 3612 7970 3668 7980
rect 2940 7634 2996 7644
rect 3836 7700 3892 7710
rect 2044 7410 2100 7420
rect 2940 7474 2996 7486
rect 2940 7422 2942 7474
rect 2994 7422 2996 7474
rect 1932 7362 1988 7374
rect 1932 7310 1934 7362
rect 1986 7310 1988 7362
rect 1932 6804 1988 7310
rect 1932 6738 1988 6748
rect 2940 6804 2996 7422
rect 2940 6738 2996 6748
rect 3388 6690 3444 6702
rect 3388 6638 3390 6690
rect 3442 6638 3444 6690
rect 1708 6578 1764 6590
rect 1708 6526 1710 6578
rect 1762 6526 1764 6578
rect 1708 6132 1764 6526
rect 2044 6580 2100 6590
rect 2044 6486 2100 6524
rect 1708 6066 1764 6076
rect 2492 6466 2548 6478
rect 3164 6468 3220 6478
rect 2492 6414 2494 6466
rect 2546 6414 2548 6466
rect 2492 6132 2548 6414
rect 2492 6066 2548 6076
rect 2940 6466 3220 6468
rect 2940 6414 3166 6466
rect 3218 6414 3220 6466
rect 2940 6412 3220 6414
rect 2940 5906 2996 6412
rect 3164 6402 3220 6412
rect 2940 5854 2942 5906
rect 2994 5854 2996 5906
rect 2940 5842 2996 5854
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5460 1988 5742
rect 1932 5394 1988 5404
rect 2044 5684 2100 5694
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 4788 1764 5070
rect 2044 5010 2100 5628
rect 3388 5684 3444 6638
rect 3836 6578 3892 7644
rect 3948 7028 4004 7980
rect 8016 7868 8280 7878
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8016 7802 8280 7812
rect 14820 7868 15084 7878
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 14820 7802 15084 7812
rect 20748 7362 20804 12908
rect 20860 9268 20916 14252
rect 22092 14308 22148 14478
rect 22764 14530 22820 16044
rect 23212 16100 23268 17612
rect 23772 18450 23828 18462
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 23772 18228 23828 18398
rect 23212 16034 23268 16044
rect 23324 16772 23380 16782
rect 22764 14478 22766 14530
rect 22818 14478 22820 14530
rect 22764 14466 22820 14478
rect 23324 14530 23380 16716
rect 23548 15316 23604 15326
rect 23772 15316 23828 18172
rect 23884 17668 23940 19182
rect 24780 19124 24836 23774
rect 25452 23826 25508 23838
rect 25452 23774 25454 23826
rect 25506 23774 25508 23826
rect 25116 23716 25172 23726
rect 24892 23714 25172 23716
rect 24892 23662 25118 23714
rect 25170 23662 25172 23714
rect 24892 23660 25172 23662
rect 24892 20020 24948 23660
rect 25116 23650 25172 23660
rect 25026 22764 25290 22774
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25026 22698 25290 22708
rect 25452 21812 25508 23774
rect 25788 23826 25844 24668
rect 25788 23774 25790 23826
rect 25842 23774 25844 23826
rect 25788 23762 25844 23774
rect 26124 23826 26180 23838
rect 26124 23774 26126 23826
rect 26178 23774 26180 23826
rect 26124 23492 26180 23774
rect 26124 23426 26180 23436
rect 26236 23380 26292 25342
rect 26348 23380 26404 26236
rect 26572 26226 26628 26236
rect 27580 26292 27636 26302
rect 26572 25284 26628 25294
rect 26908 25284 26964 25294
rect 26572 25282 26964 25284
rect 26572 25230 26574 25282
rect 26626 25230 26910 25282
rect 26962 25230 26964 25282
rect 26572 25228 26964 25230
rect 26572 25218 26628 25228
rect 26908 25218 26964 25228
rect 27468 24836 27524 24846
rect 26908 24724 26964 24734
rect 26908 24630 26964 24668
rect 26460 23716 26516 23726
rect 26908 23716 26964 23726
rect 26460 23714 26964 23716
rect 26460 23662 26462 23714
rect 26514 23662 26910 23714
rect 26962 23662 26964 23714
rect 26460 23660 26964 23662
rect 26460 23650 26516 23660
rect 26908 23650 26964 23660
rect 26908 23492 26964 23502
rect 26964 23436 27076 23492
rect 26908 23426 26964 23436
rect 26460 23380 26516 23390
rect 26348 23378 26516 23380
rect 26348 23326 26462 23378
rect 26514 23326 26516 23378
rect 26348 23324 26516 23326
rect 26236 23314 26292 23324
rect 26460 23314 26516 23324
rect 25788 23266 25844 23278
rect 25788 23214 25790 23266
rect 25842 23214 25844 23266
rect 25564 23154 25620 23166
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25564 22596 25620 23102
rect 25564 22530 25620 22540
rect 25452 21746 25508 21756
rect 25026 21196 25290 21206
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25026 21130 25290 21140
rect 25788 20804 25844 23214
rect 26124 23268 26180 23278
rect 26124 23174 26180 23212
rect 26796 22932 26852 22942
rect 26460 22260 26516 22270
rect 26460 22166 26516 22204
rect 26796 22258 26852 22876
rect 26796 22206 26798 22258
rect 26850 22206 26852 22258
rect 26796 22194 26852 22206
rect 27020 22260 27076 23436
rect 27132 23380 27188 23390
rect 27132 23286 27188 23324
rect 27468 23266 27524 24780
rect 27580 24050 27636 26236
rect 27692 26178 27748 26190
rect 27692 26126 27694 26178
rect 27746 26126 27748 26178
rect 27692 25620 27748 26126
rect 27692 25554 27748 25564
rect 27692 25282 27748 25294
rect 27692 25230 27694 25282
rect 27746 25230 27748 25282
rect 27692 24948 27748 25230
rect 27692 24882 27748 24892
rect 27692 24724 27748 24734
rect 27804 24724 27860 28252
rect 28140 27636 28196 27646
rect 28140 24946 28196 27580
rect 28428 26684 28692 26694
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28428 26618 28692 26628
rect 28140 24894 28142 24946
rect 28194 24894 28196 24946
rect 28140 24836 28196 24894
rect 28140 24770 28196 24780
rect 28252 25282 28308 25294
rect 28252 25230 28254 25282
rect 28306 25230 28308 25282
rect 27692 24722 27860 24724
rect 27692 24670 27694 24722
rect 27746 24670 27860 24722
rect 27692 24668 27860 24670
rect 27692 24658 27748 24668
rect 28252 24276 28308 25230
rect 28428 25116 28692 25126
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28428 25050 28692 25060
rect 27580 23998 27582 24050
rect 27634 23998 27636 24050
rect 27580 23986 27636 23998
rect 28140 24220 28252 24276
rect 27468 23214 27470 23266
rect 27522 23214 27524 23266
rect 27468 23202 27524 23214
rect 27580 23716 27636 23726
rect 27132 22260 27188 22270
rect 27020 22258 27188 22260
rect 27020 22206 27134 22258
rect 27186 22206 27188 22258
rect 27020 22204 27188 22206
rect 27132 22194 27188 22204
rect 27468 22260 27524 22270
rect 27468 22166 27524 22204
rect 27468 21812 27524 21822
rect 27580 21812 27636 23660
rect 27804 23266 27860 23278
rect 27804 23214 27806 23266
rect 27858 23214 27860 23266
rect 27804 23156 27860 23214
rect 28140 23266 28196 24220
rect 28252 24210 28308 24220
rect 28140 23214 28142 23266
rect 28194 23214 28196 23266
rect 28140 23202 28196 23214
rect 28252 23714 28308 23726
rect 28252 23662 28254 23714
rect 28306 23662 28308 23714
rect 27804 23090 27860 23100
rect 27804 22596 27860 22606
rect 27804 22258 27860 22540
rect 27804 22206 27806 22258
rect 27858 22206 27860 22258
rect 27804 22194 27860 22206
rect 28028 22372 28084 22382
rect 28252 22372 28308 23662
rect 28428 23548 28692 23558
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28428 23482 28692 23492
rect 28028 22370 28308 22372
rect 28028 22318 28030 22370
rect 28082 22318 28308 22370
rect 28028 22316 28308 22318
rect 27468 21810 27636 21812
rect 27468 21758 27470 21810
rect 27522 21758 27636 21810
rect 27468 21756 27636 21758
rect 27804 21812 27860 21822
rect 27468 21746 27524 21756
rect 27804 21718 27860 21756
rect 28028 21588 28084 22316
rect 28428 21980 28692 21990
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28428 21914 28692 21924
rect 28028 21522 28084 21532
rect 28140 21586 28196 21598
rect 28140 21534 28142 21586
rect 28194 21534 28196 21586
rect 27132 21476 27188 21486
rect 27132 21382 27188 21420
rect 28140 21476 28196 21534
rect 28140 20916 28196 21420
rect 28140 20850 28196 20860
rect 25788 20738 25844 20748
rect 26908 20804 26964 20814
rect 26908 20710 26964 20748
rect 28028 20690 28084 20702
rect 28028 20638 28030 20690
rect 28082 20638 28084 20690
rect 28028 20244 28084 20638
rect 28428 20412 28692 20422
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28428 20346 28692 20356
rect 28028 20178 28084 20188
rect 24892 19954 24948 19964
rect 26908 20020 26964 20030
rect 26908 19926 26964 19964
rect 28028 19906 28084 19918
rect 28028 19854 28030 19906
rect 28082 19854 28084 19906
rect 25026 19628 25290 19638
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25026 19562 25290 19572
rect 28028 19572 28084 19854
rect 28028 19506 28084 19516
rect 24780 19058 24836 19068
rect 27468 19124 27524 19134
rect 27804 19124 27860 19134
rect 27468 19122 27636 19124
rect 27468 19070 27470 19122
rect 27522 19070 27636 19122
rect 27468 19068 27636 19070
rect 27468 19058 27524 19068
rect 26124 19010 26180 19022
rect 26124 18958 26126 19010
rect 26178 18958 26180 19010
rect 23996 18228 24052 18238
rect 24556 18228 24612 18238
rect 23996 18226 24164 18228
rect 23996 18174 23998 18226
rect 24050 18174 24164 18226
rect 23996 18172 24164 18174
rect 23996 18162 24052 18172
rect 23884 17602 23940 17612
rect 24108 17554 24164 18172
rect 24108 17502 24110 17554
rect 24162 17502 24164 17554
rect 24108 17490 24164 17502
rect 24332 17780 24388 17790
rect 24332 16098 24388 17724
rect 24332 16046 24334 16098
rect 24386 16046 24388 16098
rect 24332 16034 24388 16046
rect 24556 15538 24612 18172
rect 26124 18228 26180 18958
rect 26908 19012 26964 19022
rect 27132 19012 27188 19022
rect 26908 19010 27076 19012
rect 26908 18958 26910 19010
rect 26962 18958 27076 19010
rect 26908 18956 27076 18958
rect 26908 18946 26964 18956
rect 26236 18340 26292 18350
rect 26236 18246 26292 18284
rect 27020 18228 27076 18956
rect 27132 19010 27412 19012
rect 27132 18958 27134 19010
rect 27186 18958 27412 19010
rect 27132 18956 27412 18958
rect 27132 18946 27188 18956
rect 27244 18562 27300 18574
rect 27244 18510 27246 18562
rect 27298 18510 27300 18562
rect 27244 18452 27300 18510
rect 27244 18386 27300 18396
rect 27020 18172 27188 18228
rect 26124 18162 26180 18172
rect 25026 18060 25290 18070
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25026 17994 25290 18004
rect 26124 17780 26180 17790
rect 26124 17686 26180 17724
rect 26684 17668 26740 17678
rect 24892 17444 24948 17454
rect 24892 17350 24948 17388
rect 26236 16772 26292 16782
rect 26236 16678 26292 16716
rect 25026 16492 25290 16502
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25026 16426 25290 16436
rect 26684 16210 26740 17612
rect 27132 17554 27188 18172
rect 27132 17502 27134 17554
rect 27186 17502 27188 17554
rect 27132 17490 27188 17502
rect 27244 17444 27300 17454
rect 27244 16994 27300 17388
rect 27244 16942 27246 16994
rect 27298 16942 27300 16994
rect 27244 16930 27300 16942
rect 27356 16772 27412 18956
rect 26684 16158 26686 16210
rect 26738 16158 26740 16210
rect 26684 16146 26740 16158
rect 27020 16716 27412 16772
rect 24668 16100 24724 16110
rect 24668 16006 24724 16044
rect 26348 15988 26404 15998
rect 24556 15486 24558 15538
rect 24610 15486 24612 15538
rect 24556 15474 24612 15486
rect 25228 15874 25284 15886
rect 25228 15822 25230 15874
rect 25282 15822 25284 15874
rect 23604 15260 23828 15316
rect 24332 15316 24388 15326
rect 23548 15204 23604 15260
rect 24332 15222 24388 15260
rect 25228 15316 25284 15822
rect 25228 15250 25284 15260
rect 25676 15316 25732 15326
rect 25676 15222 25732 15260
rect 23324 14478 23326 14530
rect 23378 14478 23380 14530
rect 23324 14466 23380 14478
rect 23436 15202 23604 15204
rect 23436 15150 23550 15202
rect 23602 15150 23604 15202
rect 23436 15148 23604 15150
rect 22092 14242 22148 14252
rect 22316 14306 22372 14318
rect 22316 14254 22318 14306
rect 22370 14254 22372 14306
rect 21624 14140 21888 14150
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21624 14074 21888 14084
rect 21308 13860 21364 13870
rect 21308 13766 21364 13804
rect 21980 13634 22036 13646
rect 21980 13582 21982 13634
rect 22034 13582 22036 13634
rect 21420 12738 21476 12750
rect 21420 12686 21422 12738
rect 21474 12686 21476 12738
rect 21420 12068 21476 12686
rect 21624 12572 21888 12582
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21624 12506 21888 12516
rect 21420 11396 21476 12012
rect 21308 11394 21476 11396
rect 21308 11342 21422 11394
rect 21474 11342 21476 11394
rect 21308 11340 21476 11342
rect 21308 10610 21364 11340
rect 21420 11330 21476 11340
rect 21868 11396 21924 11406
rect 21980 11396 22036 13582
rect 22204 12962 22260 12974
rect 22204 12910 22206 12962
rect 22258 12910 22260 12962
rect 22204 12068 22260 12910
rect 22316 12740 22372 14254
rect 23436 14308 23492 15148
rect 23548 15138 23604 15148
rect 25564 15202 25620 15214
rect 25564 15150 25566 15202
rect 25618 15150 25620 15202
rect 25026 14924 25290 14934
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25026 14858 25290 14868
rect 25564 14418 25620 15150
rect 26348 14754 26404 15932
rect 27020 15314 27076 16716
rect 27020 15262 27022 15314
rect 27074 15262 27076 15314
rect 27020 15250 27076 15262
rect 27580 15316 27636 19068
rect 27804 19030 27860 19068
rect 28140 19124 28196 19134
rect 28140 19122 28308 19124
rect 28140 19070 28142 19122
rect 28194 19070 28308 19122
rect 28140 19068 28308 19070
rect 28140 19058 28196 19068
rect 28252 18676 28308 19068
rect 28428 18844 28692 18854
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28428 18778 28692 18788
rect 28252 18582 28308 18620
rect 27804 17556 27860 17566
rect 27692 15988 27748 15998
rect 27692 15894 27748 15932
rect 27692 15540 27748 15550
rect 27804 15540 27860 17500
rect 28428 17276 28692 17286
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28428 17210 28692 17220
rect 27692 15538 27860 15540
rect 27692 15486 27694 15538
rect 27746 15486 27860 15538
rect 27692 15484 27860 15486
rect 28140 16884 28196 16894
rect 27692 15474 27748 15484
rect 27580 15260 27860 15316
rect 26348 14702 26350 14754
rect 26402 14702 26404 14754
rect 26348 14690 26404 14702
rect 26908 15204 26964 15214
rect 26908 14642 26964 15148
rect 26908 14590 26910 14642
rect 26962 14590 26964 14642
rect 26908 14578 26964 14590
rect 25564 14366 25566 14418
rect 25618 14366 25620 14418
rect 25564 14354 25620 14366
rect 26572 14530 26628 14542
rect 26572 14478 26574 14530
rect 26626 14478 26628 14530
rect 23436 14242 23492 14252
rect 22764 13860 22820 13870
rect 22764 13766 22820 13804
rect 25900 13636 25956 13646
rect 25452 13634 25956 13636
rect 25452 13582 25902 13634
rect 25954 13582 25956 13634
rect 25452 13580 25956 13582
rect 25026 13356 25290 13366
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25026 13290 25290 13300
rect 22316 12674 22372 12684
rect 22652 12962 22708 12974
rect 22652 12910 22654 12962
rect 22706 12910 22708 12962
rect 22652 12516 22708 12910
rect 22652 12450 22708 12460
rect 24108 12740 24164 12750
rect 22204 12002 22260 12012
rect 21868 11394 22036 11396
rect 21868 11342 21870 11394
rect 21922 11342 22036 11394
rect 21868 11340 22036 11342
rect 21868 11330 21924 11340
rect 24108 11282 24164 12684
rect 25116 12740 25172 12750
rect 25116 12646 25172 12684
rect 24444 12068 24500 12078
rect 25452 12068 25508 13580
rect 25900 13570 25956 13580
rect 26236 13636 26292 13646
rect 26572 13636 26628 14478
rect 27804 14418 27860 15260
rect 27804 14366 27806 14418
rect 27858 14366 27860 14418
rect 27804 14354 27860 14366
rect 28140 14530 28196 16828
rect 28428 15708 28692 15718
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28428 15642 28692 15652
rect 28140 14478 28142 14530
rect 28194 14478 28196 14530
rect 28140 13972 28196 14478
rect 28428 14140 28692 14150
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28428 14074 28692 14084
rect 28252 13972 28308 13982
rect 28140 13970 28308 13972
rect 28140 13918 28254 13970
rect 28306 13918 28308 13970
rect 28140 13916 28308 13918
rect 28252 13906 28308 13916
rect 26236 13634 26628 13636
rect 26236 13582 26238 13634
rect 26290 13582 26628 13634
rect 26236 13580 26628 13582
rect 25900 12964 25956 12974
rect 26236 12964 26292 13580
rect 25900 12962 26292 12964
rect 25900 12910 25902 12962
rect 25954 12910 26292 12962
rect 25900 12908 26292 12910
rect 25676 12738 25732 12750
rect 25676 12686 25678 12738
rect 25730 12686 25732 12738
rect 24500 12012 25508 12068
rect 24444 11974 24500 12012
rect 24892 11844 24948 11854
rect 24892 11618 24948 11788
rect 25026 11788 25290 11798
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25026 11722 25290 11732
rect 25452 11620 25508 12012
rect 24892 11566 24894 11618
rect 24946 11566 24948 11618
rect 24892 11554 24948 11566
rect 25228 11564 25508 11620
rect 25564 12066 25620 12078
rect 25564 12014 25566 12066
rect 25618 12014 25620 12066
rect 25228 11506 25284 11564
rect 25228 11454 25230 11506
rect 25282 11454 25284 11506
rect 25228 11442 25284 11454
rect 24108 11230 24110 11282
rect 24162 11230 24164 11282
rect 24108 11218 24164 11230
rect 21624 11004 21888 11014
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21624 10938 21888 10948
rect 25340 10836 25396 11564
rect 25564 11060 25620 12014
rect 25676 11284 25732 12686
rect 25676 11218 25732 11228
rect 25900 11060 25956 12908
rect 26012 12740 26068 12750
rect 26012 12646 26068 12684
rect 28428 12572 28692 12582
rect 26236 12516 26292 12526
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28428 12506 28692 12516
rect 26236 12066 26292 12460
rect 26236 12014 26238 12066
rect 26290 12014 26292 12066
rect 26236 12002 26292 12014
rect 27244 12290 27300 12302
rect 27244 12238 27246 12290
rect 27298 12238 27300 12290
rect 27244 11956 27300 12238
rect 27244 11890 27300 11900
rect 25564 11004 25956 11060
rect 25788 10836 25844 10846
rect 25340 10834 25844 10836
rect 25340 10782 25342 10834
rect 25394 10782 25790 10834
rect 25842 10782 25844 10834
rect 25340 10780 25844 10782
rect 25340 10770 25396 10780
rect 25788 10770 25844 10780
rect 23996 10722 24052 10734
rect 23996 10670 23998 10722
rect 24050 10670 24052 10722
rect 21308 10558 21310 10610
rect 21362 10558 21364 10610
rect 20972 10388 21028 10398
rect 20972 10294 21028 10332
rect 21308 9940 21364 10558
rect 21756 10610 21812 10622
rect 21756 10558 21758 10610
rect 21810 10558 21812 10610
rect 21756 10500 21812 10558
rect 21756 10434 21812 10444
rect 23772 10052 23828 10062
rect 23660 9996 23772 10052
rect 21420 9940 21476 9950
rect 21364 9938 21924 9940
rect 21364 9886 21422 9938
rect 21474 9886 21924 9938
rect 21364 9884 21924 9886
rect 21308 9846 21364 9884
rect 21420 9874 21476 9884
rect 21868 9828 21924 9884
rect 21868 9734 21924 9772
rect 22540 9826 22596 9838
rect 22540 9774 22542 9826
rect 22594 9774 22596 9826
rect 21624 9436 21888 9446
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21624 9370 21888 9380
rect 20860 9202 20916 9212
rect 21644 9268 21700 9278
rect 21644 9174 21700 9212
rect 22540 8932 22596 9774
rect 22540 8866 22596 8876
rect 22988 9828 23044 9838
rect 22988 8258 23044 9772
rect 23548 9268 23604 9278
rect 23548 9174 23604 9212
rect 23660 8428 23716 9996
rect 23772 9986 23828 9996
rect 22988 8206 22990 8258
rect 23042 8206 23044 8258
rect 21624 7868 21888 7878
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21624 7802 21888 7812
rect 22092 7588 22148 7598
rect 22092 7494 22148 7532
rect 20748 7310 20750 7362
rect 20802 7310 20804 7362
rect 20748 7298 20804 7310
rect 4614 7084 4878 7094
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 3948 6972 4452 7028
rect 4614 7018 4878 7028
rect 11418 7084 11682 7094
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11418 7018 11682 7028
rect 18222 7084 18486 7094
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18222 7018 18486 7028
rect 4172 6804 4228 6814
rect 4228 6748 4340 6804
rect 4172 6738 4228 6748
rect 3836 6526 3838 6578
rect 3890 6526 3892 6578
rect 3836 6514 3892 6526
rect 4172 6580 4228 6590
rect 4284 6580 4340 6748
rect 4396 6692 4452 6972
rect 4732 6692 4788 6702
rect 4396 6690 4788 6692
rect 4396 6638 4734 6690
rect 4786 6638 4788 6690
rect 4396 6636 4788 6638
rect 4732 6626 4788 6636
rect 22988 6692 23044 8206
rect 23548 8372 23716 8428
rect 23772 9268 23828 9278
rect 23548 8258 23604 8372
rect 23548 8206 23550 8258
rect 23602 8206 23604 8258
rect 23548 8194 23604 8206
rect 23100 7588 23156 7598
rect 23100 6914 23156 7532
rect 23548 7364 23604 7374
rect 23772 7364 23828 9212
rect 23996 7698 24052 10670
rect 24780 10388 24836 10398
rect 24780 10386 24948 10388
rect 24780 10334 24782 10386
rect 24834 10334 24948 10386
rect 24780 10332 24948 10334
rect 24780 10322 24836 10332
rect 24780 9604 24836 9614
rect 24556 9602 24836 9604
rect 24556 9550 24782 9602
rect 24834 9550 24836 9602
rect 24556 9548 24836 9550
rect 24332 9268 24388 9278
rect 24332 9042 24388 9212
rect 24556 9266 24612 9548
rect 24780 9538 24836 9548
rect 24556 9214 24558 9266
rect 24610 9214 24612 9266
rect 24556 9202 24612 9214
rect 24332 8990 24334 9042
rect 24386 8990 24388 9042
rect 24332 8978 24388 8990
rect 24892 8428 24948 10332
rect 25026 10220 25290 10230
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25026 10154 25290 10164
rect 25564 10164 25620 10174
rect 25564 10050 25620 10108
rect 25564 9998 25566 10050
rect 25618 9998 25620 10050
rect 25564 9986 25620 9998
rect 25788 9828 25844 9838
rect 25900 9828 25956 11004
rect 26684 11506 26740 11518
rect 26684 11454 26686 11506
rect 26738 11454 26740 11506
rect 26236 10500 26292 10510
rect 26236 10406 26292 10444
rect 26684 10052 26740 11454
rect 27692 11284 27748 11294
rect 27692 11190 27748 11228
rect 28428 11004 28692 11014
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28428 10938 28692 10948
rect 27244 10722 27300 10734
rect 27244 10670 27246 10722
rect 27298 10670 27300 10722
rect 26684 9986 26740 9996
rect 26908 10388 26964 10398
rect 25788 9826 25956 9828
rect 25788 9774 25790 9826
rect 25842 9774 25956 9826
rect 25788 9772 25956 9774
rect 26908 9826 26964 10332
rect 27244 10164 27300 10670
rect 27244 10098 27300 10108
rect 27692 10052 27748 10062
rect 27692 9958 27748 9996
rect 26908 9774 26910 9826
rect 26962 9774 26964 9826
rect 25452 9268 25508 9278
rect 25788 9268 25844 9772
rect 26908 9762 26964 9774
rect 25508 9212 25844 9268
rect 25900 9602 25956 9614
rect 25900 9550 25902 9602
rect 25954 9550 25956 9602
rect 25452 9174 25508 9212
rect 25026 8652 25290 8662
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25026 8586 25290 8596
rect 24892 8372 25396 8428
rect 23996 7646 23998 7698
rect 24050 7646 24052 7698
rect 23996 7634 24052 7646
rect 25340 7586 25396 8372
rect 25900 8034 25956 9550
rect 28428 9436 28692 9446
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28428 9370 28692 9380
rect 27244 9154 27300 9166
rect 27244 9102 27246 9154
rect 27298 9102 27300 9154
rect 26236 8932 26292 8942
rect 26236 8838 26292 8876
rect 27244 8428 27300 9102
rect 26572 8372 27300 8428
rect 27692 8372 27748 8382
rect 26572 8370 26628 8372
rect 26572 8318 26574 8370
rect 26626 8318 26628 8370
rect 26572 8306 26628 8318
rect 27692 8278 27748 8316
rect 27020 8260 27076 8270
rect 27020 8258 27412 8260
rect 27020 8206 27022 8258
rect 27074 8206 27412 8258
rect 27020 8204 27412 8206
rect 27020 8194 27076 8204
rect 25900 7982 25902 8034
rect 25954 7982 25956 8034
rect 25900 7970 25956 7982
rect 25340 7534 25342 7586
rect 25394 7534 25396 7586
rect 25340 7522 25396 7534
rect 23996 7474 24052 7486
rect 23996 7422 23998 7474
rect 24050 7422 24052 7474
rect 23996 7364 24052 7422
rect 26460 7364 26516 7374
rect 23548 7362 24052 7364
rect 23548 7310 23550 7362
rect 23602 7310 24052 7362
rect 23548 7308 24052 7310
rect 23548 7298 23604 7308
rect 23100 6862 23102 6914
rect 23154 6862 23156 6914
rect 23100 6850 23156 6862
rect 23772 6916 23828 6926
rect 22988 6598 23044 6636
rect 4284 6524 4564 6580
rect 4172 6486 4228 6524
rect 4508 6466 4564 6524
rect 4508 6414 4510 6466
rect 4562 6414 4564 6466
rect 4508 6402 4564 6414
rect 8016 6300 8280 6310
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8016 6234 8280 6244
rect 14820 6300 15084 6310
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 14820 6234 15084 6244
rect 21624 6300 21888 6310
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21624 6234 21888 6244
rect 10332 6020 10388 6030
rect 10332 6018 10836 6020
rect 10332 5966 10334 6018
rect 10386 5966 10836 6018
rect 10332 5964 10836 5966
rect 10332 5954 10388 5964
rect 9212 5908 9268 5918
rect 3388 5618 3444 5628
rect 9100 5852 9212 5908
rect 4614 5516 4878 5526
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4614 5450 4878 5460
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 1708 4722 1764 4732
rect 2492 4788 2548 5070
rect 2492 4722 2548 4732
rect 8016 4732 8280 4742
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8016 4666 8280 4676
rect 8988 4226 9044 4238
rect 8988 4174 8990 4226
rect 9042 4174 9044 4226
rect 4614 3948 4878 3958
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4614 3882 4878 3892
rect 8540 3556 8596 3566
rect 8988 3556 9044 4174
rect 8540 3554 9044 3556
rect 8540 3502 8542 3554
rect 8594 3502 9044 3554
rect 8540 3500 9044 3502
rect 8016 3164 8280 3174
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8016 3098 8280 3108
rect 8540 2548 8596 3500
rect 9100 3444 9156 5852
rect 9212 5842 9268 5852
rect 9996 5908 10052 5918
rect 9996 5814 10052 5852
rect 9996 5122 10052 5134
rect 9996 5070 9998 5122
rect 10050 5070 10052 5122
rect 9660 4226 9716 4238
rect 9660 4174 9662 4226
rect 9714 4174 9716 4226
rect 9660 3444 9716 4174
rect 8764 3388 9156 3444
rect 9436 3442 9716 3444
rect 9436 3390 9662 3442
rect 9714 3390 9716 3442
rect 9436 3388 9716 3390
rect 8764 3330 8820 3388
rect 8764 3278 8766 3330
rect 8818 3278 8820 3330
rect 8764 3266 8820 3278
rect 8540 2492 8820 2548
rect 8764 800 8820 2492
rect 9436 800 9492 3388
rect 9660 3378 9716 3388
rect 9996 3442 10052 5070
rect 10220 4898 10276 4910
rect 10220 4846 10222 4898
rect 10274 4846 10276 4898
rect 10220 4564 10276 4846
rect 10332 4564 10388 4574
rect 10220 4562 10388 4564
rect 10220 4510 10334 4562
rect 10386 4510 10388 4562
rect 10220 4508 10388 4510
rect 10332 4498 10388 4508
rect 10780 4340 10836 5964
rect 11116 6018 11172 6030
rect 11116 5966 11118 6018
rect 11170 5966 11172 6018
rect 10892 5906 10948 5918
rect 10892 5854 10894 5906
rect 10946 5854 10948 5906
rect 10892 4564 10948 5854
rect 11116 4676 11172 5966
rect 23324 5908 23380 5918
rect 11418 5516 11682 5526
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11418 5450 11682 5460
rect 18222 5516 18486 5526
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18222 5450 18486 5460
rect 20412 5012 20468 5022
rect 20188 5010 20468 5012
rect 20188 4958 20414 5010
rect 20466 4958 20468 5010
rect 20188 4956 20468 4958
rect 14820 4732 15084 4742
rect 11116 4610 11172 4620
rect 13132 4676 13188 4686
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 14820 4666 15084 4676
rect 10892 4498 10948 4508
rect 11900 4564 11956 4574
rect 11900 4470 11956 4508
rect 10780 4284 11060 4340
rect 11004 3554 11060 4284
rect 12124 4338 12180 4350
rect 12124 4286 12126 4338
rect 12178 4286 12180 4338
rect 11564 4228 11620 4238
rect 12124 4228 12180 4286
rect 11564 4226 12180 4228
rect 11564 4174 11566 4226
rect 11618 4174 12180 4226
rect 11564 4172 12180 4174
rect 11564 4162 11620 4172
rect 11004 3502 11006 3554
rect 11058 3502 11060 3554
rect 11004 3490 11060 3502
rect 11116 4114 11172 4126
rect 11116 4062 11118 4114
rect 11170 4062 11172 4114
rect 9996 3390 9998 3442
rect 10050 3390 10052 3442
rect 9996 3378 10052 3390
rect 11116 2212 11172 4062
rect 11418 3948 11682 3958
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11418 3882 11682 3892
rect 11788 3780 11844 4172
rect 11676 3724 11844 3780
rect 11452 3668 11508 3678
rect 10332 2156 11172 2212
rect 11228 3666 11508 3668
rect 11228 3614 11454 3666
rect 11506 3614 11508 3666
rect 11228 3612 11508 3614
rect 10332 980 10388 2156
rect 11228 980 11284 3612
rect 11452 3602 11508 3612
rect 11676 2884 11732 3724
rect 10108 924 10388 980
rect 10780 924 11284 980
rect 11452 2828 11732 2884
rect 12124 3668 12180 3678
rect 10108 800 10164 924
rect 10780 800 10836 924
rect 11452 800 11508 2828
rect 12124 800 12180 3612
rect 13132 3554 13188 4620
rect 18222 3948 18486 3958
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18222 3882 18486 3892
rect 13580 3668 13636 3678
rect 13580 3574 13636 3612
rect 13132 3502 13134 3554
rect 13186 3502 13188 3554
rect 13132 3490 13188 3502
rect 19964 3556 20020 3566
rect 19964 3554 20132 3556
rect 19964 3502 19966 3554
rect 20018 3502 20132 3554
rect 19964 3500 20132 3502
rect 19964 3490 20020 3500
rect 20076 3220 20132 3500
rect 20188 3442 20244 4956
rect 20412 4946 20468 4956
rect 20748 4900 20804 4910
rect 20748 4898 21140 4900
rect 20748 4846 20750 4898
rect 20802 4846 21140 4898
rect 20748 4844 21140 4846
rect 20748 4834 20804 4844
rect 20188 3390 20190 3442
rect 20242 3390 20244 3442
rect 20188 3378 20244 3390
rect 20412 4226 20468 4238
rect 20412 4174 20414 4226
rect 20466 4174 20468 4226
rect 20412 3220 20468 4174
rect 21084 3554 21140 4844
rect 21624 4732 21888 4742
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21624 4666 21888 4676
rect 21532 3668 21588 3678
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 21420 3666 21588 3668
rect 21420 3614 21534 3666
rect 21586 3614 21588 3666
rect 21420 3612 21588 3614
rect 14820 3164 15084 3174
rect 20076 3164 20468 3220
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 14820 3098 15084 3108
rect 20188 800 20244 3164
rect 20860 924 21140 980
rect 20860 800 20916 924
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21084 756 21140 924
rect 21420 756 21476 3612
rect 21532 3602 21588 3612
rect 23100 3554 23156 3566
rect 23100 3502 23102 3554
rect 23154 3502 23156 3554
rect 22764 3444 22820 3454
rect 23100 3444 23156 3502
rect 22764 3442 23156 3444
rect 22764 3390 22766 3442
rect 22818 3390 23156 3442
rect 22764 3388 23156 3390
rect 22764 3378 22820 3388
rect 21624 3164 21888 3174
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21624 3098 21888 3108
rect 23100 2772 23156 3388
rect 23324 3442 23380 5852
rect 23772 4338 23828 6860
rect 23884 6466 23940 6478
rect 23884 6414 23886 6466
rect 23938 6414 23940 6466
rect 23884 6132 23940 6414
rect 23884 6066 23940 6076
rect 23996 6020 24052 7308
rect 26236 7362 26516 7364
rect 26236 7310 26462 7362
rect 26514 7310 26516 7362
rect 26236 7308 26516 7310
rect 25026 7084 25290 7094
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25026 7018 25290 7028
rect 25676 6804 25732 6814
rect 25564 6748 25676 6804
rect 25452 6132 25508 6142
rect 25452 6038 25508 6076
rect 23996 5926 24052 5964
rect 24668 6018 24724 6030
rect 24668 5966 24670 6018
rect 24722 5966 24724 6018
rect 24332 5908 24388 5918
rect 24332 5814 24388 5852
rect 24108 5236 24164 5246
rect 23996 5012 24052 5022
rect 23996 4562 24052 4956
rect 23996 4510 23998 4562
rect 24050 4510 24052 4562
rect 23996 4498 24052 4510
rect 23772 4286 23774 4338
rect 23826 4286 23828 4338
rect 23772 4274 23828 4286
rect 23436 4226 23492 4238
rect 23436 4174 23438 4226
rect 23490 4174 23492 4226
rect 23436 3556 23492 4174
rect 23772 3556 23828 3566
rect 23436 3554 23828 3556
rect 23436 3502 23774 3554
rect 23826 3502 23828 3554
rect 23436 3500 23828 3502
rect 23324 3390 23326 3442
rect 23378 3390 23380 3442
rect 23324 3378 23380 3390
rect 23100 2706 23156 2716
rect 23772 1428 23828 3500
rect 23996 3444 24052 3454
rect 24108 3444 24164 5180
rect 24332 5124 24388 5134
rect 24556 5124 24612 5134
rect 24332 5122 24612 5124
rect 24332 5070 24334 5122
rect 24386 5070 24558 5122
rect 24610 5070 24612 5122
rect 24332 5068 24612 5070
rect 24332 5058 24388 5068
rect 23996 3442 24164 3444
rect 23996 3390 23998 3442
rect 24050 3390 24164 3442
rect 23996 3388 24164 3390
rect 24332 4338 24388 4350
rect 24332 4286 24334 4338
rect 24386 4286 24388 4338
rect 24332 3444 24388 4286
rect 23996 3378 24052 3388
rect 24332 3378 24388 3388
rect 24556 2100 24612 5068
rect 24668 5124 24724 5966
rect 25026 5516 25290 5526
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25026 5450 25290 5460
rect 24668 5058 24724 5068
rect 25340 5124 25396 5134
rect 25564 5124 25620 6748
rect 25676 6738 25732 6748
rect 26236 6690 26292 7308
rect 26460 7298 26516 7308
rect 27132 7362 27188 7374
rect 27132 7310 27134 7362
rect 27186 7310 27188 7362
rect 26236 6638 26238 6690
rect 26290 6638 26292 6690
rect 26236 6626 26292 6638
rect 26796 6692 26852 6702
rect 27132 6692 27188 7310
rect 26852 6636 27188 6692
rect 27244 6804 27300 6814
rect 26796 6598 26852 6636
rect 27132 6468 27188 6478
rect 27244 6468 27300 6748
rect 27132 6466 27300 6468
rect 27132 6414 27134 6466
rect 27186 6414 27300 6466
rect 27132 6412 27300 6414
rect 27132 6402 27188 6412
rect 25676 6020 25732 6030
rect 25676 5906 25732 5964
rect 26908 5908 26964 5918
rect 25676 5854 25678 5906
rect 25730 5854 25732 5906
rect 25676 5842 25732 5854
rect 26348 5906 26964 5908
rect 26348 5854 26910 5906
rect 26962 5854 26964 5906
rect 26348 5852 26964 5854
rect 25340 5122 25620 5124
rect 25340 5070 25342 5122
rect 25394 5070 25620 5122
rect 25340 5068 25620 5070
rect 25900 5236 25956 5246
rect 25900 5122 25956 5180
rect 25900 5070 25902 5122
rect 25954 5070 25956 5122
rect 25340 5058 25396 5068
rect 25900 5058 25956 5070
rect 24892 4898 24948 4910
rect 24892 4846 24894 4898
rect 24946 4846 24948 4898
rect 24892 4676 24948 4846
rect 24892 4610 24948 4620
rect 25452 4900 25508 4910
rect 24668 4452 24724 4462
rect 25228 4452 25284 4462
rect 24668 4450 25284 4452
rect 24668 4398 24670 4450
rect 24722 4398 25230 4450
rect 25282 4398 25284 4450
rect 24668 4396 25284 4398
rect 24668 4386 24724 4396
rect 25228 4386 25284 4396
rect 25026 3948 25290 3958
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25026 3882 25290 3892
rect 25452 3778 25508 4844
rect 25564 4900 25620 4910
rect 26236 4900 26292 4910
rect 25564 4898 25732 4900
rect 25564 4846 25566 4898
rect 25618 4846 25732 4898
rect 25564 4844 25732 4846
rect 25564 4834 25620 4844
rect 25676 4564 25732 4844
rect 26124 4898 26292 4900
rect 26124 4846 26238 4898
rect 26290 4846 26292 4898
rect 26124 4844 26292 4846
rect 25900 4676 25956 4686
rect 25788 4564 25844 4574
rect 25676 4508 25788 4564
rect 25788 4498 25844 4508
rect 25564 4452 25620 4462
rect 25564 4358 25620 4396
rect 25900 4450 25956 4620
rect 25900 4398 25902 4450
rect 25954 4398 25956 4450
rect 25900 4386 25956 4398
rect 25452 3726 25454 3778
rect 25506 3726 25508 3778
rect 25452 3714 25508 3726
rect 26124 3554 26180 4844
rect 26236 4834 26292 4844
rect 26236 4564 26292 4574
rect 26348 4564 26404 5852
rect 26908 5842 26964 5852
rect 27356 5684 27412 8204
rect 28140 8148 28196 8158
rect 27692 7476 27748 7486
rect 27244 5628 27412 5684
rect 27468 7250 27524 7262
rect 27468 7198 27470 7250
rect 27522 7198 27524 7250
rect 27468 6578 27524 7198
rect 27468 6526 27470 6578
rect 27522 6526 27524 6578
rect 26908 5124 26964 5134
rect 26908 5030 26964 5068
rect 27244 5012 27300 5628
rect 27244 4946 27300 4956
rect 27356 5460 27412 5470
rect 26236 4562 26404 4564
rect 26236 4510 26238 4562
rect 26290 4510 26404 4562
rect 26236 4508 26404 4510
rect 26908 4564 26964 4574
rect 26236 4498 26292 4508
rect 26908 4470 26964 4508
rect 26460 4452 26516 4462
rect 26516 4396 26628 4452
rect 26460 4386 26516 4396
rect 26124 3502 26126 3554
rect 26178 3502 26180 3554
rect 26124 3490 26180 3502
rect 26572 3554 26628 4396
rect 27356 3778 27412 5404
rect 27468 4116 27524 6526
rect 27580 6804 27636 6814
rect 27580 5234 27636 6748
rect 27692 6130 27748 7420
rect 27804 7362 27860 7374
rect 27804 7310 27806 7362
rect 27858 7310 27860 7362
rect 27804 7250 27860 7310
rect 27804 7198 27806 7250
rect 27858 7198 27860 7250
rect 27804 7186 27860 7198
rect 27804 6916 27860 6926
rect 27804 6578 27860 6860
rect 28140 6692 28196 8092
rect 28428 7868 28692 7878
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28428 7802 28692 7812
rect 28140 6690 28308 6692
rect 28140 6638 28142 6690
rect 28194 6638 28308 6690
rect 28140 6636 28308 6638
rect 28140 6626 28196 6636
rect 27804 6526 27806 6578
rect 27858 6526 27860 6578
rect 27804 6514 27860 6526
rect 27692 6078 27694 6130
rect 27746 6078 27748 6130
rect 27692 6066 27748 6078
rect 28252 6130 28308 6636
rect 28428 6300 28692 6310
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28428 6234 28692 6244
rect 28252 6078 28254 6130
rect 28306 6078 28308 6130
rect 28252 6066 28308 6078
rect 27580 5182 27582 5234
rect 27634 5182 27636 5234
rect 27580 5170 27636 5182
rect 27692 5908 27748 5918
rect 27692 4562 27748 5852
rect 28428 4732 28692 4742
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28428 4666 28692 4676
rect 27692 4510 27694 4562
rect 27746 4510 27748 4562
rect 27692 4498 27748 4510
rect 27468 4050 27524 4060
rect 27356 3726 27358 3778
rect 27410 3726 27412 3778
rect 27356 3714 27412 3726
rect 26572 3502 26574 3554
rect 26626 3502 26628 3554
rect 26572 3490 26628 3502
rect 24892 3444 24948 3454
rect 24892 3350 24948 3388
rect 28428 3164 28692 3174
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28428 3098 28692 3108
rect 24668 2100 24724 2110
rect 24556 2044 24668 2100
rect 24668 2034 24724 2044
rect 23772 1362 23828 1372
rect 21084 700 21476 756
<< via2 >>
rect 1820 28252 1876 28308
rect 3724 27580 3780 27636
rect 3388 26908 3444 26964
rect 2044 26236 2100 26292
rect 1932 25564 1988 25620
rect 1820 25452 1876 25508
rect 2940 26290 2996 26292
rect 2940 26238 2942 26290
rect 2942 26238 2994 26290
rect 2994 26238 2996 26290
rect 2940 26236 2996 26238
rect 3948 26236 4004 26292
rect 3276 25506 3332 25508
rect 3276 25454 3278 25506
rect 3278 25454 3330 25506
rect 3330 25454 3332 25506
rect 3276 25452 3332 25454
rect 2156 25282 2212 25284
rect 2156 25230 2158 25282
rect 2158 25230 2210 25282
rect 2210 25230 2212 25282
rect 2156 25228 2212 25230
rect 2940 25282 2996 25284
rect 2940 25230 2942 25282
rect 2942 25230 2994 25282
rect 2994 25230 2996 25282
rect 2940 25228 2996 25230
rect 3500 25228 3556 25284
rect 2940 24834 2996 24836
rect 2940 24782 2942 24834
rect 2942 24782 2994 24834
rect 2994 24782 2996 24834
rect 2940 24780 2996 24782
rect 2716 24668 2772 24724
rect 2380 24220 2436 24276
rect 2268 23884 2324 23940
rect 2044 23826 2100 23828
rect 2044 23774 2046 23826
rect 2046 23774 2098 23826
rect 2098 23774 2100 23826
rect 2044 23772 2100 23774
rect 1708 23548 1764 23604
rect 3164 24220 3220 24276
rect 4614 25898 4670 25900
rect 4614 25846 4616 25898
rect 4616 25846 4668 25898
rect 4668 25846 4670 25898
rect 4614 25844 4670 25846
rect 4718 25898 4774 25900
rect 4718 25846 4720 25898
rect 4720 25846 4772 25898
rect 4772 25846 4774 25898
rect 4718 25844 4774 25846
rect 4822 25898 4878 25900
rect 4822 25846 4824 25898
rect 4824 25846 4876 25898
rect 4876 25846 4878 25898
rect 4822 25844 4878 25846
rect 6412 26290 6468 26292
rect 6412 26238 6414 26290
rect 6414 26238 6466 26290
rect 6466 26238 6468 26290
rect 6412 26236 6468 26238
rect 6076 25452 6132 25508
rect 5964 25394 6020 25396
rect 5964 25342 5966 25394
rect 5966 25342 6018 25394
rect 6018 25342 6020 25394
rect 5964 25340 6020 25342
rect 6972 26236 7028 26292
rect 7420 25564 7476 25620
rect 8016 26682 8072 26684
rect 8016 26630 8018 26682
rect 8018 26630 8070 26682
rect 8070 26630 8072 26682
rect 8016 26628 8072 26630
rect 8120 26682 8176 26684
rect 8120 26630 8122 26682
rect 8122 26630 8174 26682
rect 8174 26630 8176 26682
rect 8120 26628 8176 26630
rect 8224 26682 8280 26684
rect 8224 26630 8226 26682
rect 8226 26630 8278 26682
rect 8278 26630 8280 26682
rect 8224 26628 8280 26630
rect 7868 26290 7924 26292
rect 7868 26238 7870 26290
rect 7870 26238 7922 26290
rect 7922 26238 7924 26290
rect 7868 26236 7924 26238
rect 8316 26236 8372 26292
rect 8764 26402 8820 26404
rect 8764 26350 8766 26402
rect 8766 26350 8818 26402
rect 8818 26350 8820 26402
rect 8764 26348 8820 26350
rect 6748 25228 6804 25284
rect 9324 25228 9380 25284
rect 4956 24834 5012 24836
rect 4956 24782 4958 24834
rect 4958 24782 5010 24834
rect 5010 24782 5012 24834
rect 4956 24780 5012 24782
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 4614 24330 4670 24332
rect 4614 24278 4616 24330
rect 4616 24278 4668 24330
rect 4668 24278 4670 24330
rect 4614 24276 4670 24278
rect 4718 24330 4774 24332
rect 4718 24278 4720 24330
rect 4720 24278 4772 24330
rect 4772 24278 4774 24330
rect 4718 24276 4774 24278
rect 4822 24330 4878 24332
rect 4822 24278 4824 24330
rect 4824 24278 4876 24330
rect 4876 24278 4878 24330
rect 4822 24276 4878 24278
rect 4956 23938 5012 23940
rect 4956 23886 4958 23938
rect 4958 23886 5010 23938
rect 5010 23886 5012 23938
rect 4956 23884 5012 23886
rect 8016 25114 8072 25116
rect 8016 25062 8018 25114
rect 8018 25062 8070 25114
rect 8070 25062 8072 25114
rect 8016 25060 8072 25062
rect 8120 25114 8176 25116
rect 8120 25062 8122 25114
rect 8122 25062 8174 25114
rect 8174 25062 8176 25114
rect 8120 25060 8176 25062
rect 8224 25114 8280 25116
rect 8224 25062 8226 25114
rect 8226 25062 8278 25114
rect 8278 25062 8280 25114
rect 8224 25060 8280 25062
rect 7868 23884 7924 23940
rect 5180 23772 5236 23828
rect 2940 23660 2996 23716
rect 1708 22876 1764 22932
rect 2492 22876 2548 22932
rect 4732 23714 4788 23716
rect 4732 23662 4734 23714
rect 4734 23662 4786 23714
rect 4786 23662 4788 23714
rect 4732 23660 4788 23662
rect 4614 22762 4670 22764
rect 4614 22710 4616 22762
rect 4616 22710 4668 22762
rect 4668 22710 4670 22762
rect 4614 22708 4670 22710
rect 4718 22762 4774 22764
rect 4718 22710 4720 22762
rect 4720 22710 4772 22762
rect 4772 22710 4774 22762
rect 4718 22708 4774 22710
rect 4822 22762 4878 22764
rect 4822 22710 4824 22762
rect 4824 22710 4876 22762
rect 4876 22710 4878 22762
rect 4822 22708 4878 22710
rect 2268 22204 2324 22260
rect 2156 21532 2212 21588
rect 2940 21810 2996 21812
rect 2940 21758 2942 21810
rect 2942 21758 2994 21810
rect 2994 21758 2996 21810
rect 2940 21756 2996 21758
rect 5740 21756 5796 21812
rect 4614 21194 4670 21196
rect 4614 21142 4616 21194
rect 4616 21142 4668 21194
rect 4668 21142 4670 21194
rect 4614 21140 4670 21142
rect 4718 21194 4774 21196
rect 4718 21142 4720 21194
rect 4720 21142 4772 21194
rect 4772 21142 4774 21194
rect 4718 21140 4774 21142
rect 4822 21194 4878 21196
rect 4822 21142 4824 21194
rect 4824 21142 4876 21194
rect 4876 21142 4878 21194
rect 4822 21140 4878 21142
rect 2380 20860 2436 20916
rect 2044 20690 2100 20692
rect 2044 20638 2046 20690
rect 2046 20638 2098 20690
rect 2098 20638 2100 20690
rect 2044 20636 2100 20638
rect 10108 26348 10164 26404
rect 10668 25452 10724 25508
rect 10332 25228 10388 25284
rect 8016 23546 8072 23548
rect 8016 23494 8018 23546
rect 8018 23494 8070 23546
rect 8070 23494 8072 23546
rect 8016 23492 8072 23494
rect 8120 23546 8176 23548
rect 8120 23494 8122 23546
rect 8122 23494 8174 23546
rect 8174 23494 8176 23546
rect 8120 23492 8176 23494
rect 8224 23546 8280 23548
rect 8224 23494 8226 23546
rect 8226 23494 8278 23546
rect 8278 23494 8280 23546
rect 8224 23492 8280 23494
rect 10780 25340 10836 25396
rect 12796 26460 12852 26516
rect 13580 26460 13636 26516
rect 11452 26012 11508 26068
rect 12124 26012 12180 26068
rect 11418 25898 11474 25900
rect 11418 25846 11420 25898
rect 11420 25846 11472 25898
rect 11472 25846 11474 25898
rect 11418 25844 11474 25846
rect 11522 25898 11578 25900
rect 11522 25846 11524 25898
rect 11524 25846 11576 25898
rect 11576 25846 11578 25898
rect 11522 25844 11578 25846
rect 11626 25898 11682 25900
rect 11626 25846 11628 25898
rect 11628 25846 11680 25898
rect 11680 25846 11682 25898
rect 11626 25844 11682 25846
rect 11452 25564 11508 25620
rect 11676 25282 11732 25284
rect 11676 25230 11678 25282
rect 11678 25230 11730 25282
rect 11730 25230 11732 25282
rect 11676 25228 11732 25230
rect 12124 25228 12180 25284
rect 11418 24330 11474 24332
rect 11418 24278 11420 24330
rect 11420 24278 11472 24330
rect 11472 24278 11474 24330
rect 11418 24276 11474 24278
rect 11522 24330 11578 24332
rect 11522 24278 11524 24330
rect 11524 24278 11576 24330
rect 11576 24278 11578 24330
rect 11522 24276 11578 24278
rect 11626 24330 11682 24332
rect 11626 24278 11628 24330
rect 11628 24278 11680 24330
rect 11680 24278 11682 24330
rect 11626 24276 11682 24278
rect 11340 23938 11396 23940
rect 11340 23886 11342 23938
rect 11342 23886 11394 23938
rect 11394 23886 11396 23938
rect 11340 23884 11396 23886
rect 11676 23826 11732 23828
rect 11676 23774 11678 23826
rect 11678 23774 11730 23826
rect 11730 23774 11732 23826
rect 11676 23772 11732 23774
rect 14812 26796 14868 26852
rect 14820 26682 14876 26684
rect 14820 26630 14822 26682
rect 14822 26630 14874 26682
rect 14874 26630 14876 26682
rect 14820 26628 14876 26630
rect 14924 26682 14980 26684
rect 14924 26630 14926 26682
rect 14926 26630 14978 26682
rect 14978 26630 14980 26682
rect 14924 26628 14980 26630
rect 15028 26682 15084 26684
rect 15028 26630 15030 26682
rect 15030 26630 15082 26682
rect 15082 26630 15084 26682
rect 15028 26628 15084 26630
rect 14820 25114 14876 25116
rect 14820 25062 14822 25114
rect 14822 25062 14874 25114
rect 14874 25062 14876 25114
rect 14820 25060 14876 25062
rect 14924 25114 14980 25116
rect 14924 25062 14926 25114
rect 14926 25062 14978 25114
rect 14978 25062 14980 25114
rect 14924 25060 14980 25062
rect 15028 25114 15084 25116
rect 15028 25062 15030 25114
rect 15030 25062 15082 25114
rect 15082 25062 15084 25114
rect 15028 25060 15084 25062
rect 15820 26796 15876 26852
rect 15372 25452 15428 25508
rect 15932 25506 15988 25508
rect 15932 25454 15934 25506
rect 15934 25454 15986 25506
rect 15986 25454 15988 25506
rect 15932 25452 15988 25454
rect 15708 25282 15764 25284
rect 15708 25230 15710 25282
rect 15710 25230 15762 25282
rect 15762 25230 15764 25282
rect 15708 25228 15764 25230
rect 15260 23772 15316 23828
rect 18172 26460 18228 26516
rect 18222 25898 18278 25900
rect 18222 25846 18224 25898
rect 18224 25846 18276 25898
rect 18276 25846 18278 25898
rect 18222 25844 18278 25846
rect 18326 25898 18382 25900
rect 18326 25846 18328 25898
rect 18328 25846 18380 25898
rect 18380 25846 18382 25898
rect 18326 25844 18382 25846
rect 18430 25898 18486 25900
rect 18430 25846 18432 25898
rect 18432 25846 18484 25898
rect 18484 25846 18486 25898
rect 18430 25844 18486 25846
rect 19068 26460 19124 26516
rect 20300 26236 20356 26292
rect 20412 26348 20468 26404
rect 19404 25282 19460 25284
rect 19404 25230 19406 25282
rect 19406 25230 19458 25282
rect 19458 25230 19460 25282
rect 19404 25228 19460 25230
rect 18222 24330 18278 24332
rect 18222 24278 18224 24330
rect 18224 24278 18276 24330
rect 18276 24278 18278 24330
rect 18222 24276 18278 24278
rect 18326 24330 18382 24332
rect 18326 24278 18328 24330
rect 18328 24278 18380 24330
rect 18380 24278 18382 24330
rect 18326 24276 18382 24278
rect 18430 24330 18486 24332
rect 18430 24278 18432 24330
rect 18432 24278 18484 24330
rect 18484 24278 18486 24330
rect 18430 24276 18486 24278
rect 21624 26682 21680 26684
rect 21624 26630 21626 26682
rect 21626 26630 21678 26682
rect 21678 26630 21680 26682
rect 21624 26628 21680 26630
rect 21728 26682 21784 26684
rect 21728 26630 21730 26682
rect 21730 26630 21782 26682
rect 21782 26630 21784 26682
rect 21728 26628 21784 26630
rect 21832 26682 21888 26684
rect 21832 26630 21834 26682
rect 21834 26630 21886 26682
rect 21886 26630 21888 26682
rect 21832 26628 21888 26630
rect 20972 26290 21028 26292
rect 20972 26238 20974 26290
rect 20974 26238 21026 26290
rect 21026 26238 21028 26290
rect 20972 26236 21028 26238
rect 20860 25452 20916 25508
rect 20748 25340 20804 25396
rect 20636 25228 20692 25284
rect 14820 23546 14876 23548
rect 14820 23494 14822 23546
rect 14822 23494 14874 23546
rect 14874 23494 14876 23546
rect 14820 23492 14876 23494
rect 14924 23546 14980 23548
rect 14924 23494 14926 23546
rect 14926 23494 14978 23546
rect 14978 23494 14980 23546
rect 14924 23492 14980 23494
rect 15028 23546 15084 23548
rect 15028 23494 15030 23546
rect 15030 23494 15082 23546
rect 15082 23494 15084 23546
rect 15028 23492 15084 23494
rect 21196 25004 21252 25060
rect 20972 24444 21028 24500
rect 21532 26348 21588 26404
rect 21644 25506 21700 25508
rect 21644 25454 21646 25506
rect 21646 25454 21698 25506
rect 21698 25454 21700 25506
rect 21644 25452 21700 25454
rect 21624 25114 21680 25116
rect 21624 25062 21626 25114
rect 21626 25062 21678 25114
rect 21678 25062 21680 25114
rect 21624 25060 21680 25062
rect 21728 25114 21784 25116
rect 21728 25062 21730 25114
rect 21730 25062 21782 25114
rect 21782 25062 21784 25114
rect 21728 25060 21784 25062
rect 21832 25114 21888 25116
rect 21832 25062 21834 25114
rect 21834 25062 21886 25114
rect 21886 25062 21888 25114
rect 21832 25060 21888 25062
rect 22876 25676 22932 25732
rect 23548 25676 23604 25732
rect 24220 25676 24276 25732
rect 24444 28924 24500 28980
rect 23100 25394 23156 25396
rect 23100 25342 23102 25394
rect 23102 25342 23154 25394
rect 23154 25342 23156 25394
rect 23100 25340 23156 25342
rect 27804 28252 27860 28308
rect 26124 26908 26180 26964
rect 22428 24444 22484 24500
rect 24332 24444 24388 24500
rect 21644 23826 21700 23828
rect 21644 23774 21646 23826
rect 21646 23774 21698 23826
rect 21698 23774 21700 23826
rect 21644 23772 21700 23774
rect 21624 23546 21680 23548
rect 21624 23494 21626 23546
rect 21626 23494 21678 23546
rect 21678 23494 21680 23546
rect 21624 23492 21680 23494
rect 21728 23546 21784 23548
rect 21728 23494 21730 23546
rect 21730 23494 21782 23546
rect 21782 23494 21784 23546
rect 21728 23492 21784 23494
rect 21832 23546 21888 23548
rect 21832 23494 21834 23546
rect 21834 23494 21886 23546
rect 21886 23494 21888 23546
rect 21832 23492 21888 23494
rect 25026 25898 25082 25900
rect 25026 25846 25028 25898
rect 25028 25846 25080 25898
rect 25080 25846 25082 25898
rect 25026 25844 25082 25846
rect 25130 25898 25186 25900
rect 25130 25846 25132 25898
rect 25132 25846 25184 25898
rect 25184 25846 25186 25898
rect 25130 25844 25186 25846
rect 25234 25898 25290 25900
rect 25234 25846 25236 25898
rect 25236 25846 25288 25898
rect 25288 25846 25290 25898
rect 25234 25844 25290 25846
rect 25340 25676 25396 25732
rect 24668 25282 24724 25284
rect 24668 25230 24670 25282
rect 24670 25230 24722 25282
rect 24722 25230 24724 25282
rect 24668 25228 24724 25230
rect 24556 23772 24612 23828
rect 25340 24444 25396 24500
rect 25788 24668 25844 24724
rect 25026 24330 25082 24332
rect 25026 24278 25028 24330
rect 25028 24278 25080 24330
rect 25080 24278 25082 24330
rect 25026 24276 25082 24278
rect 25130 24330 25186 24332
rect 25130 24278 25132 24330
rect 25132 24278 25184 24330
rect 25184 24278 25186 24330
rect 25130 24276 25186 24278
rect 25234 24330 25290 24332
rect 25234 24278 25236 24330
rect 25236 24278 25288 24330
rect 25288 24278 25290 24330
rect 25234 24276 25290 24278
rect 24668 23212 24724 23268
rect 24108 23100 24164 23156
rect 11418 22762 11474 22764
rect 11418 22710 11420 22762
rect 11420 22710 11472 22762
rect 11472 22710 11474 22762
rect 11418 22708 11474 22710
rect 11522 22762 11578 22764
rect 11522 22710 11524 22762
rect 11524 22710 11576 22762
rect 11576 22710 11578 22762
rect 11522 22708 11578 22710
rect 11626 22762 11682 22764
rect 11626 22710 11628 22762
rect 11628 22710 11680 22762
rect 11680 22710 11682 22762
rect 11626 22708 11682 22710
rect 18222 22762 18278 22764
rect 18222 22710 18224 22762
rect 18224 22710 18276 22762
rect 18276 22710 18278 22762
rect 18222 22708 18278 22710
rect 18326 22762 18382 22764
rect 18326 22710 18328 22762
rect 18328 22710 18380 22762
rect 18380 22710 18382 22762
rect 18326 22708 18382 22710
rect 18430 22762 18486 22764
rect 18430 22710 18432 22762
rect 18432 22710 18484 22762
rect 18484 22710 18486 22762
rect 18430 22708 18486 22710
rect 8016 21978 8072 21980
rect 8016 21926 8018 21978
rect 8018 21926 8070 21978
rect 8070 21926 8072 21978
rect 8016 21924 8072 21926
rect 8120 21978 8176 21980
rect 8120 21926 8122 21978
rect 8122 21926 8174 21978
rect 8174 21926 8176 21978
rect 8120 21924 8176 21926
rect 8224 21978 8280 21980
rect 8224 21926 8226 21978
rect 8226 21926 8278 21978
rect 8278 21926 8280 21978
rect 8224 21924 8280 21926
rect 14820 21978 14876 21980
rect 14820 21926 14822 21978
rect 14822 21926 14874 21978
rect 14874 21926 14876 21978
rect 14820 21924 14876 21926
rect 14924 21978 14980 21980
rect 14924 21926 14926 21978
rect 14926 21926 14978 21978
rect 14978 21926 14980 21978
rect 14924 21924 14980 21926
rect 15028 21978 15084 21980
rect 15028 21926 15030 21978
rect 15030 21926 15082 21978
rect 15082 21926 15084 21978
rect 15028 21924 15084 21926
rect 21624 21978 21680 21980
rect 21624 21926 21626 21978
rect 21626 21926 21678 21978
rect 21678 21926 21680 21978
rect 21624 21924 21680 21926
rect 21728 21978 21784 21980
rect 21728 21926 21730 21978
rect 21730 21926 21782 21978
rect 21782 21926 21784 21978
rect 21728 21924 21784 21926
rect 21832 21978 21888 21980
rect 21832 21926 21834 21978
rect 21834 21926 21886 21978
rect 21886 21926 21888 21978
rect 21832 21924 21888 21926
rect 20636 21644 20692 21700
rect 11418 21194 11474 21196
rect 11418 21142 11420 21194
rect 11420 21142 11472 21194
rect 11472 21142 11474 21194
rect 11418 21140 11474 21142
rect 11522 21194 11578 21196
rect 11522 21142 11524 21194
rect 11524 21142 11576 21194
rect 11576 21142 11578 21194
rect 11522 21140 11578 21142
rect 11626 21194 11682 21196
rect 11626 21142 11628 21194
rect 11628 21142 11680 21194
rect 11680 21142 11682 21194
rect 11626 21140 11682 21142
rect 18222 21194 18278 21196
rect 18222 21142 18224 21194
rect 18224 21142 18276 21194
rect 18276 21142 18278 21194
rect 18222 21140 18278 21142
rect 18326 21194 18382 21196
rect 18326 21142 18328 21194
rect 18328 21142 18380 21194
rect 18380 21142 18382 21194
rect 18326 21140 18382 21142
rect 18430 21194 18486 21196
rect 18430 21142 18432 21194
rect 18432 21142 18484 21194
rect 18484 21142 18486 21194
rect 18430 21140 18486 21142
rect 6076 20636 6132 20692
rect 12124 20860 12180 20916
rect 8016 20410 8072 20412
rect 8016 20358 8018 20410
rect 8018 20358 8070 20410
rect 8070 20358 8072 20410
rect 8016 20356 8072 20358
rect 8120 20410 8176 20412
rect 8120 20358 8122 20410
rect 8122 20358 8174 20410
rect 8174 20358 8176 20410
rect 8120 20356 8176 20358
rect 8224 20410 8280 20412
rect 8224 20358 8226 20410
rect 8226 20358 8278 20410
rect 8278 20358 8280 20410
rect 8224 20356 8280 20358
rect 1820 20242 1876 20244
rect 1820 20190 1822 20242
rect 1822 20190 1874 20242
rect 1874 20190 1876 20242
rect 1820 20188 1876 20190
rect 4614 19626 4670 19628
rect 4614 19574 4616 19626
rect 4616 19574 4668 19626
rect 4668 19574 4670 19626
rect 4614 19572 4670 19574
rect 4718 19626 4774 19628
rect 4718 19574 4720 19626
rect 4720 19574 4772 19626
rect 4772 19574 4774 19626
rect 4718 19572 4774 19574
rect 4822 19626 4878 19628
rect 4822 19574 4824 19626
rect 4824 19574 4876 19626
rect 4876 19574 4878 19626
rect 4822 19572 4878 19574
rect 7756 19292 7812 19348
rect 6300 18508 6356 18564
rect 4614 18058 4670 18060
rect 4614 18006 4616 18058
rect 4616 18006 4668 18058
rect 4668 18006 4670 18058
rect 4614 18004 4670 18006
rect 4718 18058 4774 18060
rect 4718 18006 4720 18058
rect 4720 18006 4772 18058
rect 4772 18006 4774 18058
rect 4718 18004 4774 18006
rect 4822 18058 4878 18060
rect 4822 18006 4824 18058
rect 4824 18006 4876 18058
rect 4876 18006 4878 18058
rect 4822 18004 4878 18006
rect 4844 17554 4900 17556
rect 4844 17502 4846 17554
rect 4846 17502 4898 17554
rect 4898 17502 4900 17554
rect 4844 17500 4900 17502
rect 4844 16940 4900 16996
rect 3164 16882 3220 16884
rect 3164 16830 3166 16882
rect 3166 16830 3218 16882
rect 3218 16830 3220 16882
rect 3164 16828 3220 16830
rect 4956 16828 5012 16884
rect 5404 16828 5460 16884
rect 4614 16490 4670 16492
rect 4614 16438 4616 16490
rect 4616 16438 4668 16490
rect 4668 16438 4670 16490
rect 4614 16436 4670 16438
rect 4718 16490 4774 16492
rect 4718 16438 4720 16490
rect 4720 16438 4772 16490
rect 4772 16438 4774 16490
rect 4718 16436 4774 16438
rect 4822 16490 4878 16492
rect 4822 16438 4824 16490
rect 4824 16438 4876 16490
rect 4876 16438 4878 16490
rect 4822 16436 4878 16438
rect 4956 16156 5012 16212
rect 7644 18562 7700 18564
rect 7644 18510 7646 18562
rect 7646 18510 7698 18562
rect 7698 18510 7700 18562
rect 7644 18508 7700 18510
rect 5852 17500 5908 17556
rect 6860 16940 6916 16996
rect 7084 17666 7140 17668
rect 7084 17614 7086 17666
rect 7086 17614 7138 17666
rect 7138 17614 7140 17666
rect 7084 17612 7140 17614
rect 8652 19346 8708 19348
rect 8652 19294 8654 19346
rect 8654 19294 8706 19346
rect 8706 19294 8708 19346
rect 8652 19292 8708 19294
rect 10444 19292 10500 19348
rect 8016 18842 8072 18844
rect 8016 18790 8018 18842
rect 8018 18790 8070 18842
rect 8070 18790 8072 18842
rect 8016 18788 8072 18790
rect 8120 18842 8176 18844
rect 8120 18790 8122 18842
rect 8122 18790 8174 18842
rect 8174 18790 8176 18842
rect 8120 18788 8176 18790
rect 8224 18842 8280 18844
rect 8224 18790 8226 18842
rect 8226 18790 8278 18842
rect 8278 18790 8280 18842
rect 8224 18788 8280 18790
rect 9436 18450 9492 18452
rect 9436 18398 9438 18450
rect 9438 18398 9490 18450
rect 9490 18398 9492 18450
rect 9436 18396 9492 18398
rect 10780 19068 10836 19124
rect 14476 20914 14532 20916
rect 14476 20862 14478 20914
rect 14478 20862 14530 20914
rect 14530 20862 14532 20914
rect 14476 20860 14532 20862
rect 14820 20410 14876 20412
rect 14820 20358 14822 20410
rect 14822 20358 14874 20410
rect 14874 20358 14876 20410
rect 14820 20356 14876 20358
rect 14924 20410 14980 20412
rect 14924 20358 14926 20410
rect 14926 20358 14978 20410
rect 14978 20358 14980 20410
rect 14924 20356 14980 20358
rect 15028 20410 15084 20412
rect 15028 20358 15030 20410
rect 15030 20358 15082 20410
rect 15082 20358 15084 20410
rect 15028 20356 15084 20358
rect 11418 19626 11474 19628
rect 11418 19574 11420 19626
rect 11420 19574 11472 19626
rect 11472 19574 11474 19626
rect 11418 19572 11474 19574
rect 11522 19626 11578 19628
rect 11522 19574 11524 19626
rect 11524 19574 11576 19626
rect 11576 19574 11578 19626
rect 11522 19572 11578 19574
rect 11626 19626 11682 19628
rect 11626 19574 11628 19626
rect 11628 19574 11680 19626
rect 11680 19574 11682 19626
rect 11626 19572 11682 19574
rect 11452 19346 11508 19348
rect 11452 19294 11454 19346
rect 11454 19294 11506 19346
rect 11506 19294 11508 19346
rect 11452 19292 11508 19294
rect 13916 19292 13972 19348
rect 12460 19122 12516 19124
rect 12460 19070 12462 19122
rect 12462 19070 12514 19122
rect 12514 19070 12516 19122
rect 12460 19068 12516 19070
rect 11228 18396 11284 18452
rect 11418 18058 11474 18060
rect 11418 18006 11420 18058
rect 11420 18006 11472 18058
rect 11472 18006 11474 18058
rect 11418 18004 11474 18006
rect 11522 18058 11578 18060
rect 11522 18006 11524 18058
rect 11524 18006 11576 18058
rect 11576 18006 11578 18058
rect 11522 18004 11578 18006
rect 11626 18058 11682 18060
rect 11626 18006 11628 18058
rect 11628 18006 11680 18058
rect 11680 18006 11682 18058
rect 11626 18004 11682 18006
rect 13244 18450 13300 18452
rect 13244 18398 13246 18450
rect 13246 18398 13298 18450
rect 13298 18398 13300 18450
rect 13244 18396 13300 18398
rect 13132 18338 13188 18340
rect 13132 18286 13134 18338
rect 13134 18286 13186 18338
rect 13186 18286 13188 18338
rect 13132 18284 13188 18286
rect 15372 19628 15428 19684
rect 15260 19346 15316 19348
rect 15260 19294 15262 19346
rect 15262 19294 15314 19346
rect 15314 19294 15316 19346
rect 15260 19292 15316 19294
rect 14252 18956 14308 19012
rect 9436 17612 9492 17668
rect 8016 17274 8072 17276
rect 8016 17222 8018 17274
rect 8018 17222 8070 17274
rect 8070 17222 8072 17274
rect 8016 17220 8072 17222
rect 8120 17274 8176 17276
rect 8120 17222 8122 17274
rect 8122 17222 8174 17274
rect 8174 17222 8176 17274
rect 8120 17220 8176 17222
rect 8224 17274 8280 17276
rect 8224 17222 8226 17274
rect 8226 17222 8278 17274
rect 8278 17222 8280 17274
rect 8224 17220 8280 17222
rect 7084 16828 7140 16884
rect 7532 16882 7588 16884
rect 7532 16830 7534 16882
rect 7534 16830 7586 16882
rect 7586 16830 7588 16882
rect 7532 16828 7588 16830
rect 6300 16604 6356 16660
rect 5516 15372 5572 15428
rect 4614 14922 4670 14924
rect 4614 14870 4616 14922
rect 4616 14870 4668 14922
rect 4668 14870 4670 14922
rect 4614 14868 4670 14870
rect 4718 14922 4774 14924
rect 4718 14870 4720 14922
rect 4720 14870 4772 14922
rect 4772 14870 4774 14922
rect 4718 14868 4774 14870
rect 4822 14922 4878 14924
rect 4822 14870 4824 14922
rect 4824 14870 4876 14922
rect 4876 14870 4878 14922
rect 4822 14868 4878 14870
rect 2716 14700 2772 14756
rect 3948 14754 4004 14756
rect 3948 14702 3950 14754
rect 3950 14702 4002 14754
rect 4002 14702 4004 14754
rect 3948 14700 4004 14702
rect 3500 14364 3556 14420
rect 2380 13132 2436 13188
rect 3276 13186 3332 13188
rect 3276 13134 3278 13186
rect 3278 13134 3330 13186
rect 3330 13134 3332 13186
rect 3276 13132 3332 13134
rect 2380 12908 2436 12964
rect 1596 12348 1652 12404
rect 1708 12684 1764 12740
rect 1708 12124 1764 12180
rect 3388 12796 3444 12852
rect 2492 12738 2548 12740
rect 2492 12686 2494 12738
rect 2494 12686 2546 12738
rect 2546 12686 2548 12738
rect 2492 12684 2548 12686
rect 2604 12348 2660 12404
rect 2044 10332 2100 10388
rect 1820 10108 1876 10164
rect 7308 16658 7364 16660
rect 7308 16606 7310 16658
rect 7310 16606 7362 16658
rect 7362 16606 7364 16658
rect 7308 16604 7364 16606
rect 6636 15932 6692 15988
rect 7308 15986 7364 15988
rect 7308 15934 7310 15986
rect 7310 15934 7362 15986
rect 7362 15934 7364 15986
rect 7308 15932 7364 15934
rect 8016 15706 8072 15708
rect 8016 15654 8018 15706
rect 8018 15654 8070 15706
rect 8070 15654 8072 15706
rect 8016 15652 8072 15654
rect 8120 15706 8176 15708
rect 8120 15654 8122 15706
rect 8122 15654 8174 15706
rect 8174 15654 8176 15706
rect 8120 15652 8176 15654
rect 8224 15706 8280 15708
rect 8224 15654 8226 15706
rect 8226 15654 8278 15706
rect 8278 15654 8280 15706
rect 8224 15652 8280 15654
rect 7980 15426 8036 15428
rect 7980 15374 7982 15426
rect 7982 15374 8034 15426
rect 8034 15374 8036 15426
rect 7980 15372 8036 15374
rect 6748 14418 6804 14420
rect 6748 14366 6750 14418
rect 6750 14366 6802 14418
rect 6802 14366 6804 14418
rect 6748 14364 6804 14366
rect 4732 13468 4788 13524
rect 4614 13354 4670 13356
rect 4614 13302 4616 13354
rect 4616 13302 4668 13354
rect 4668 13302 4670 13354
rect 4614 13300 4670 13302
rect 4718 13354 4774 13356
rect 4718 13302 4720 13354
rect 4720 13302 4772 13354
rect 4772 13302 4774 13354
rect 4718 13300 4774 13302
rect 4822 13354 4878 13356
rect 4822 13302 4824 13354
rect 4824 13302 4876 13354
rect 4876 13302 4878 13354
rect 4822 13300 4878 13302
rect 4172 12796 4228 12852
rect 6524 13468 6580 13524
rect 6188 13356 6244 13412
rect 5180 12908 5236 12964
rect 5516 12962 5572 12964
rect 5516 12910 5518 12962
rect 5518 12910 5570 12962
rect 5570 12910 5572 12962
rect 5516 12908 5572 12910
rect 4620 12796 4676 12852
rect 4620 11900 4676 11956
rect 4614 11786 4670 11788
rect 4614 11734 4616 11786
rect 4616 11734 4668 11786
rect 4668 11734 4670 11786
rect 4614 11732 4670 11734
rect 4718 11786 4774 11788
rect 4718 11734 4720 11786
rect 4720 11734 4772 11786
rect 4772 11734 4774 11786
rect 4718 11732 4774 11734
rect 4822 11786 4878 11788
rect 4822 11734 4824 11786
rect 4824 11734 4876 11786
rect 4876 11734 4878 11786
rect 4822 11732 4878 11734
rect 5964 11676 6020 11732
rect 3164 11004 3220 11060
rect 3052 10610 3108 10612
rect 3052 10558 3054 10610
rect 3054 10558 3106 10610
rect 3106 10558 3108 10610
rect 3052 10556 3108 10558
rect 4844 11004 4900 11060
rect 3724 10556 3780 10612
rect 4614 10218 4670 10220
rect 4614 10166 4616 10218
rect 4616 10166 4668 10218
rect 4668 10166 4670 10218
rect 4614 10164 4670 10166
rect 4718 10218 4774 10220
rect 4718 10166 4720 10218
rect 4720 10166 4772 10218
rect 4772 10166 4774 10218
rect 4718 10164 4774 10166
rect 4822 10218 4878 10220
rect 4822 10166 4824 10218
rect 4824 10166 4876 10218
rect 4876 10166 4878 10218
rect 4822 10164 4878 10166
rect 10220 16828 10276 16884
rect 9996 16210 10052 16212
rect 9996 16158 9998 16210
rect 9998 16158 10050 16210
rect 10050 16158 10052 16210
rect 9996 16156 10052 16158
rect 11418 16490 11474 16492
rect 11418 16438 11420 16490
rect 11420 16438 11472 16490
rect 11472 16438 11474 16490
rect 11418 16436 11474 16438
rect 11522 16490 11578 16492
rect 11522 16438 11524 16490
rect 11524 16438 11576 16490
rect 11576 16438 11578 16490
rect 11522 16436 11578 16438
rect 11626 16490 11682 16492
rect 11626 16438 11628 16490
rect 11628 16438 11680 16490
rect 11680 16438 11682 16490
rect 11626 16436 11682 16438
rect 13692 16716 13748 16772
rect 12908 16098 12964 16100
rect 12908 16046 12910 16098
rect 12910 16046 12962 16098
rect 12962 16046 12964 16098
rect 12908 16044 12964 16046
rect 14140 16716 14196 16772
rect 13692 16098 13748 16100
rect 13692 16046 13694 16098
rect 13694 16046 13746 16098
rect 13746 16046 13748 16098
rect 13692 16044 13748 16046
rect 11900 15820 11956 15876
rect 8016 14138 8072 14140
rect 8016 14086 8018 14138
rect 8018 14086 8070 14138
rect 8070 14086 8072 14138
rect 8016 14084 8072 14086
rect 8120 14138 8176 14140
rect 8120 14086 8122 14138
rect 8122 14086 8174 14138
rect 8174 14086 8176 14138
rect 8120 14084 8176 14086
rect 8224 14138 8280 14140
rect 8224 14086 8226 14138
rect 8226 14086 8278 14138
rect 8278 14086 8280 14138
rect 8224 14084 8280 14086
rect 9212 13804 9268 13860
rect 6972 13356 7028 13412
rect 6972 12908 7028 12964
rect 7868 12908 7924 12964
rect 6636 10444 6692 10500
rect 7532 10498 7588 10500
rect 7532 10446 7534 10498
rect 7534 10446 7586 10498
rect 7586 10446 7588 10498
rect 7532 10444 7588 10446
rect 9996 13580 10052 13636
rect 8988 12908 9044 12964
rect 8016 12570 8072 12572
rect 8016 12518 8018 12570
rect 8018 12518 8070 12570
rect 8070 12518 8072 12570
rect 8016 12516 8072 12518
rect 8120 12570 8176 12572
rect 8120 12518 8122 12570
rect 8122 12518 8174 12570
rect 8174 12518 8176 12570
rect 8120 12516 8176 12518
rect 8224 12570 8280 12572
rect 8224 12518 8226 12570
rect 8226 12518 8278 12570
rect 8278 12518 8280 12570
rect 8224 12516 8280 12518
rect 8988 12236 9044 12292
rect 8540 11676 8596 11732
rect 9100 11676 9156 11732
rect 8016 11002 8072 11004
rect 8016 10950 8018 11002
rect 8018 10950 8070 11002
rect 8070 10950 8072 11002
rect 8016 10948 8072 10950
rect 8120 11002 8176 11004
rect 8120 10950 8122 11002
rect 8122 10950 8174 11002
rect 8174 10950 8176 11002
rect 8120 10948 8176 10950
rect 8224 11002 8280 11004
rect 8224 10950 8226 11002
rect 8226 10950 8278 11002
rect 8278 10950 8280 11002
rect 8224 10948 8280 10950
rect 9772 12290 9828 12292
rect 9772 12238 9774 12290
rect 9774 12238 9826 12290
rect 9826 12238 9828 12290
rect 9772 12236 9828 12238
rect 11418 14922 11474 14924
rect 11418 14870 11420 14922
rect 11420 14870 11472 14922
rect 11472 14870 11474 14922
rect 11418 14868 11474 14870
rect 11522 14922 11578 14924
rect 11522 14870 11524 14922
rect 11524 14870 11576 14922
rect 11576 14870 11578 14922
rect 11522 14868 11578 14870
rect 11626 14922 11682 14924
rect 11626 14870 11628 14922
rect 11628 14870 11680 14922
rect 11680 14870 11682 14922
rect 11626 14868 11682 14870
rect 13580 15874 13636 15876
rect 13580 15822 13582 15874
rect 13582 15822 13634 15874
rect 13634 15822 13636 15874
rect 13580 15820 13636 15822
rect 13020 14306 13076 14308
rect 13020 14254 13022 14306
rect 13022 14254 13074 14306
rect 13074 14254 13076 14306
rect 13020 14252 13076 14254
rect 13916 14252 13972 14308
rect 11788 13858 11844 13860
rect 11788 13806 11790 13858
rect 11790 13806 11842 13858
rect 11842 13806 11844 13858
rect 11788 13804 11844 13806
rect 10780 13634 10836 13636
rect 10780 13582 10782 13634
rect 10782 13582 10834 13634
rect 10834 13582 10836 13634
rect 10780 13580 10836 13582
rect 14820 18842 14876 18844
rect 14820 18790 14822 18842
rect 14822 18790 14874 18842
rect 14874 18790 14876 18842
rect 14820 18788 14876 18790
rect 14924 18842 14980 18844
rect 14924 18790 14926 18842
rect 14926 18790 14978 18842
rect 14978 18790 14980 18842
rect 14924 18788 14980 18790
rect 15028 18842 15084 18844
rect 15028 18790 15030 18842
rect 15030 18790 15082 18842
rect 15082 18790 15084 18842
rect 15028 18788 15084 18790
rect 15484 18284 15540 18340
rect 15932 19740 15988 19796
rect 14588 17612 14644 17668
rect 15260 17666 15316 17668
rect 15260 17614 15262 17666
rect 15262 17614 15314 17666
rect 15314 17614 15316 17666
rect 15260 17612 15316 17614
rect 16268 19628 16324 19684
rect 17612 19852 17668 19908
rect 16940 18620 16996 18676
rect 18396 19740 18452 19796
rect 18222 19626 18278 19628
rect 18222 19574 18224 19626
rect 18224 19574 18276 19626
rect 18276 19574 18278 19626
rect 18222 19572 18278 19574
rect 18326 19626 18382 19628
rect 18326 19574 18328 19626
rect 18328 19574 18380 19626
rect 18380 19574 18382 19626
rect 18326 19572 18382 19574
rect 18430 19626 18486 19628
rect 18430 19574 18432 19626
rect 18432 19574 18484 19626
rect 18484 19574 18486 19626
rect 18430 19572 18486 19574
rect 18956 18956 19012 19012
rect 17164 18396 17220 18452
rect 16380 18284 16436 18340
rect 14820 17274 14876 17276
rect 14820 17222 14822 17274
rect 14822 17222 14874 17274
rect 14874 17222 14876 17274
rect 14820 17220 14876 17222
rect 14924 17274 14980 17276
rect 14924 17222 14926 17274
rect 14926 17222 14978 17274
rect 14978 17222 14980 17274
rect 14924 17220 14980 17222
rect 15028 17274 15084 17276
rect 15028 17222 15030 17274
rect 15030 17222 15082 17274
rect 15082 17222 15084 17274
rect 15028 17220 15084 17222
rect 14252 13580 14308 13636
rect 11418 13354 11474 13356
rect 11418 13302 11420 13354
rect 11420 13302 11472 13354
rect 11472 13302 11474 13354
rect 11418 13300 11474 13302
rect 11522 13354 11578 13356
rect 11522 13302 11524 13354
rect 11524 13302 11576 13354
rect 11576 13302 11578 13354
rect 11522 13300 11578 13302
rect 11626 13354 11682 13356
rect 11626 13302 11628 13354
rect 11628 13302 11680 13354
rect 11680 13302 11682 13354
rect 11626 13300 11682 13302
rect 12460 12962 12516 12964
rect 12460 12910 12462 12962
rect 12462 12910 12514 12962
rect 12514 12910 12516 12962
rect 12460 12908 12516 12910
rect 10220 11676 10276 11732
rect 11418 11786 11474 11788
rect 11418 11734 11420 11786
rect 11420 11734 11472 11786
rect 11472 11734 11474 11786
rect 11418 11732 11474 11734
rect 11522 11786 11578 11788
rect 11522 11734 11524 11786
rect 11524 11734 11576 11786
rect 11576 11734 11578 11786
rect 11522 11732 11578 11734
rect 11626 11786 11682 11788
rect 11626 11734 11628 11786
rect 11628 11734 11680 11786
rect 11680 11734 11682 11786
rect 11626 11732 11682 11734
rect 10108 10780 10164 10836
rect 12348 10780 12404 10836
rect 9324 10668 9380 10724
rect 11788 10722 11844 10724
rect 11788 10670 11790 10722
rect 11790 10670 11842 10722
rect 11842 10670 11844 10722
rect 11788 10668 11844 10670
rect 9996 10444 10052 10500
rect 7868 9884 7924 9940
rect 9772 10332 9828 10388
rect 9548 9826 9604 9828
rect 9548 9774 9550 9826
rect 9550 9774 9602 9826
rect 9602 9774 9604 9826
rect 9548 9772 9604 9774
rect 5516 9660 5572 9716
rect 7644 9714 7700 9716
rect 7644 9662 7646 9714
rect 7646 9662 7698 9714
rect 7698 9662 7700 9714
rect 7644 9660 7700 9662
rect 8016 9434 8072 9436
rect 8016 9382 8018 9434
rect 8018 9382 8070 9434
rect 8070 9382 8072 9434
rect 8016 9380 8072 9382
rect 8120 9434 8176 9436
rect 8120 9382 8122 9434
rect 8122 9382 8174 9434
rect 8174 9382 8176 9434
rect 8120 9380 8176 9382
rect 8224 9434 8280 9436
rect 8224 9382 8226 9434
rect 8226 9382 8278 9434
rect 8278 9382 8280 9434
rect 8224 9380 8280 9382
rect 10780 10498 10836 10500
rect 10780 10446 10782 10498
rect 10782 10446 10834 10498
rect 10834 10446 10836 10498
rect 10780 10444 10836 10446
rect 11418 10218 11474 10220
rect 11418 10166 11420 10218
rect 11420 10166 11472 10218
rect 11472 10166 11474 10218
rect 11418 10164 11474 10166
rect 11522 10218 11578 10220
rect 11522 10166 11524 10218
rect 11524 10166 11576 10218
rect 11576 10166 11578 10218
rect 11522 10164 11578 10166
rect 11626 10218 11682 10220
rect 11626 10166 11628 10218
rect 11628 10166 11680 10218
rect 11680 10166 11682 10218
rect 11626 10164 11682 10166
rect 12460 9660 12516 9716
rect 18732 18450 18788 18452
rect 18732 18398 18734 18450
rect 18734 18398 18786 18450
rect 18786 18398 18788 18450
rect 18732 18396 18788 18398
rect 18172 18284 18228 18340
rect 17164 17612 17220 17668
rect 18222 18058 18278 18060
rect 18222 18006 18224 18058
rect 18224 18006 18276 18058
rect 18276 18006 18278 18058
rect 18222 18004 18278 18006
rect 18326 18058 18382 18060
rect 18326 18006 18328 18058
rect 18328 18006 18380 18058
rect 18380 18006 18382 18058
rect 18326 18004 18382 18006
rect 18430 18058 18486 18060
rect 18430 18006 18432 18058
rect 18432 18006 18484 18058
rect 18484 18006 18486 18058
rect 18430 18004 18486 18006
rect 19292 20076 19348 20132
rect 22204 21698 22260 21700
rect 22204 21646 22206 21698
rect 22206 21646 22258 21698
rect 22258 21646 22260 21698
rect 22204 21644 22260 21646
rect 21624 20410 21680 20412
rect 21624 20358 21626 20410
rect 21626 20358 21678 20410
rect 21678 20358 21680 20410
rect 21624 20356 21680 20358
rect 21728 20410 21784 20412
rect 21728 20358 21730 20410
rect 21730 20358 21782 20410
rect 21782 20358 21784 20410
rect 21728 20356 21784 20358
rect 21832 20410 21888 20412
rect 21832 20358 21834 20410
rect 21834 20358 21886 20410
rect 21886 20358 21888 20410
rect 21832 20356 21888 20358
rect 21196 20076 21252 20132
rect 21196 19906 21252 19908
rect 21196 19854 21198 19906
rect 21198 19854 21250 19906
rect 21250 19854 21252 19906
rect 21196 19852 21252 19854
rect 22204 18956 22260 19012
rect 21624 18842 21680 18844
rect 21624 18790 21626 18842
rect 21626 18790 21678 18842
rect 21678 18790 21680 18842
rect 21624 18788 21680 18790
rect 21728 18842 21784 18844
rect 21728 18790 21730 18842
rect 21730 18790 21782 18842
rect 21782 18790 21784 18842
rect 21728 18788 21784 18790
rect 21832 18842 21888 18844
rect 21832 18790 21834 18842
rect 21834 18790 21886 18842
rect 21886 18790 21888 18842
rect 21832 18788 21888 18790
rect 19404 18620 19460 18676
rect 20076 18508 20132 18564
rect 19404 18396 19460 18452
rect 19068 18284 19124 18340
rect 19404 17612 19460 17668
rect 16380 16716 16436 16772
rect 15932 15874 15988 15876
rect 15932 15822 15934 15874
rect 15934 15822 15986 15874
rect 15986 15822 15988 15874
rect 15932 15820 15988 15822
rect 14820 15706 14876 15708
rect 14820 15654 14822 15706
rect 14822 15654 14874 15706
rect 14874 15654 14876 15706
rect 14820 15652 14876 15654
rect 14924 15706 14980 15708
rect 14924 15654 14926 15706
rect 14926 15654 14978 15706
rect 14978 15654 14980 15706
rect 14924 15652 14980 15654
rect 15028 15706 15084 15708
rect 15028 15654 15030 15706
rect 15030 15654 15082 15706
rect 15082 15654 15084 15706
rect 15028 15652 15084 15654
rect 18222 16490 18278 16492
rect 18222 16438 18224 16490
rect 18224 16438 18276 16490
rect 18276 16438 18278 16490
rect 18222 16436 18278 16438
rect 18326 16490 18382 16492
rect 18326 16438 18328 16490
rect 18328 16438 18380 16490
rect 18380 16438 18382 16490
rect 18326 16436 18382 16438
rect 18430 16490 18486 16492
rect 18430 16438 18432 16490
rect 18432 16438 18484 16490
rect 18484 16438 18486 16490
rect 18430 16436 18486 16438
rect 17500 15820 17556 15876
rect 14820 14138 14876 14140
rect 14820 14086 14822 14138
rect 14822 14086 14874 14138
rect 14874 14086 14876 14138
rect 14820 14084 14876 14086
rect 14924 14138 14980 14140
rect 14924 14086 14926 14138
rect 14926 14086 14978 14138
rect 14978 14086 14980 14138
rect 14924 14084 14980 14086
rect 15028 14138 15084 14140
rect 15028 14086 15030 14138
rect 15030 14086 15082 14138
rect 15082 14086 15084 14138
rect 15028 14084 15084 14086
rect 15036 13634 15092 13636
rect 15036 13582 15038 13634
rect 15038 13582 15090 13634
rect 15090 13582 15092 13634
rect 15036 13580 15092 13582
rect 18222 14922 18278 14924
rect 18222 14870 18224 14922
rect 18224 14870 18276 14922
rect 18276 14870 18278 14922
rect 18222 14868 18278 14870
rect 18326 14922 18382 14924
rect 18326 14870 18328 14922
rect 18328 14870 18380 14922
rect 18380 14870 18382 14922
rect 18326 14868 18382 14870
rect 18430 14922 18486 14924
rect 18430 14870 18432 14922
rect 18432 14870 18484 14922
rect 18484 14870 18486 14922
rect 18430 14868 18486 14870
rect 19628 18284 19684 18340
rect 21644 18562 21700 18564
rect 21644 18510 21646 18562
rect 21646 18510 21698 18562
rect 21698 18510 21700 18562
rect 21644 18508 21700 18510
rect 22428 18450 22484 18452
rect 22428 18398 22430 18450
rect 22430 18398 22482 18450
rect 22482 18398 22484 18450
rect 22428 18396 22484 18398
rect 21868 18284 21924 18340
rect 19068 15148 19124 15204
rect 14820 12570 14876 12572
rect 14820 12518 14822 12570
rect 14822 12518 14874 12570
rect 14874 12518 14876 12570
rect 14820 12516 14876 12518
rect 14924 12570 14980 12572
rect 14924 12518 14926 12570
rect 14926 12518 14978 12570
rect 14978 12518 14980 12570
rect 14924 12516 14980 12518
rect 15028 12570 15084 12572
rect 15028 12518 15030 12570
rect 15030 12518 15082 12570
rect 15082 12518 15084 12570
rect 15028 12516 15084 12518
rect 14812 12178 14868 12180
rect 14812 12126 14814 12178
rect 14814 12126 14866 12178
rect 14866 12126 14868 12178
rect 14812 12124 14868 12126
rect 13916 11452 13972 11508
rect 11900 8930 11956 8932
rect 11900 8878 11902 8930
rect 11902 8878 11954 8930
rect 11954 8878 11956 8930
rect 11900 8876 11956 8878
rect 13244 10610 13300 10612
rect 13244 10558 13246 10610
rect 13246 10558 13298 10610
rect 13298 10558 13300 10610
rect 13244 10556 13300 10558
rect 12908 9772 12964 9828
rect 12684 8876 12740 8932
rect 4614 8650 4670 8652
rect 4614 8598 4616 8650
rect 4616 8598 4668 8650
rect 4668 8598 4670 8650
rect 4614 8596 4670 8598
rect 4718 8650 4774 8652
rect 4718 8598 4720 8650
rect 4720 8598 4772 8650
rect 4772 8598 4774 8650
rect 4718 8596 4774 8598
rect 4822 8650 4878 8652
rect 4822 8598 4824 8650
rect 4824 8598 4876 8650
rect 4876 8598 4878 8650
rect 4822 8596 4878 8598
rect 11418 8650 11474 8652
rect 11418 8598 11420 8650
rect 11420 8598 11472 8650
rect 11472 8598 11474 8650
rect 11418 8596 11474 8598
rect 11522 8650 11578 8652
rect 11522 8598 11524 8650
rect 11524 8598 11576 8650
rect 11576 8598 11578 8650
rect 11522 8596 11578 8598
rect 11626 8650 11682 8652
rect 11626 8598 11628 8650
rect 11628 8598 11680 8650
rect 11680 8598 11682 8650
rect 11626 8596 11682 8598
rect 3388 8092 3444 8148
rect 4060 8146 4116 8148
rect 4060 8094 4062 8146
rect 4062 8094 4114 8146
rect 4114 8094 4116 8146
rect 4060 8092 4116 8094
rect 16268 11506 16324 11508
rect 16268 11454 16270 11506
rect 16270 11454 16322 11506
rect 16322 11454 16324 11506
rect 16268 11452 16324 11454
rect 16268 11228 16324 11284
rect 14820 11002 14876 11004
rect 14820 10950 14822 11002
rect 14822 10950 14874 11002
rect 14874 10950 14876 11002
rect 14820 10948 14876 10950
rect 14924 11002 14980 11004
rect 14924 10950 14926 11002
rect 14926 10950 14978 11002
rect 14978 10950 14980 11002
rect 14924 10948 14980 10950
rect 15028 11002 15084 11004
rect 15028 10950 15030 11002
rect 15030 10950 15082 11002
rect 15082 10950 15084 11002
rect 15028 10948 15084 10950
rect 17276 11282 17332 11284
rect 17276 11230 17278 11282
rect 17278 11230 17330 11282
rect 17330 11230 17332 11282
rect 17276 11228 17332 11230
rect 14476 10556 14532 10612
rect 14140 9826 14196 9828
rect 14140 9774 14142 9826
rect 14142 9774 14194 9826
rect 14194 9774 14196 9826
rect 14140 9772 14196 9774
rect 13916 9714 13972 9716
rect 13916 9662 13918 9714
rect 13918 9662 13970 9714
rect 13970 9662 13972 9714
rect 13916 9660 13972 9662
rect 14140 8876 14196 8932
rect 21196 17666 21252 17668
rect 21196 17614 21198 17666
rect 21198 17614 21250 17666
rect 21250 17614 21252 17666
rect 21196 17612 21252 17614
rect 23100 18172 23156 18228
rect 23212 17612 23268 17668
rect 21624 17274 21680 17276
rect 21624 17222 21626 17274
rect 21626 17222 21678 17274
rect 21678 17222 21680 17274
rect 21624 17220 21680 17222
rect 21728 17274 21784 17276
rect 21728 17222 21730 17274
rect 21730 17222 21782 17274
rect 21782 17222 21784 17274
rect 21728 17220 21784 17222
rect 21832 17274 21888 17276
rect 21832 17222 21834 17274
rect 21834 17222 21886 17274
rect 21886 17222 21888 17274
rect 21832 17220 21888 17222
rect 22764 16044 22820 16100
rect 18222 13354 18278 13356
rect 18222 13302 18224 13354
rect 18224 13302 18276 13354
rect 18276 13302 18278 13354
rect 18222 13300 18278 13302
rect 18326 13354 18382 13356
rect 18326 13302 18328 13354
rect 18328 13302 18380 13354
rect 18380 13302 18382 13354
rect 18326 13300 18382 13302
rect 18430 13354 18486 13356
rect 18430 13302 18432 13354
rect 18432 13302 18484 13354
rect 18484 13302 18486 13354
rect 18430 13300 18486 13302
rect 21196 15874 21252 15876
rect 21196 15822 21198 15874
rect 21198 15822 21250 15874
rect 21250 15822 21252 15874
rect 21196 15820 21252 15822
rect 21624 15706 21680 15708
rect 21624 15654 21626 15706
rect 21626 15654 21678 15706
rect 21678 15654 21680 15706
rect 21624 15652 21680 15654
rect 21728 15706 21784 15708
rect 21728 15654 21730 15706
rect 21730 15654 21782 15706
rect 21782 15654 21784 15706
rect 21728 15652 21784 15654
rect 21832 15706 21888 15708
rect 21832 15654 21834 15706
rect 21834 15654 21886 15706
rect 21886 15654 21888 15706
rect 21832 15652 21888 15654
rect 21308 15202 21364 15204
rect 21308 15150 21310 15202
rect 21310 15150 21362 15202
rect 21362 15150 21364 15202
rect 21308 15148 21364 15150
rect 22316 15820 22372 15876
rect 21980 15148 22036 15204
rect 20860 14252 20916 14308
rect 19516 12178 19572 12180
rect 19516 12126 19518 12178
rect 19518 12126 19570 12178
rect 19570 12126 19572 12178
rect 19516 12124 19572 12126
rect 20748 12908 20804 12964
rect 18222 11786 18278 11788
rect 18222 11734 18224 11786
rect 18224 11734 18276 11786
rect 18276 11734 18278 11786
rect 18222 11732 18278 11734
rect 18326 11786 18382 11788
rect 18326 11734 18328 11786
rect 18328 11734 18380 11786
rect 18380 11734 18382 11786
rect 18326 11732 18382 11734
rect 18430 11786 18486 11788
rect 18430 11734 18432 11786
rect 18432 11734 18484 11786
rect 18484 11734 18486 11786
rect 18430 11732 18486 11734
rect 17948 11452 18004 11508
rect 14700 9826 14756 9828
rect 14700 9774 14702 9826
rect 14702 9774 14754 9826
rect 14754 9774 14756 9826
rect 14700 9772 14756 9774
rect 15484 9826 15540 9828
rect 15484 9774 15486 9826
rect 15486 9774 15538 9826
rect 15538 9774 15540 9826
rect 15484 9772 15540 9774
rect 14820 9434 14876 9436
rect 14820 9382 14822 9434
rect 14822 9382 14874 9434
rect 14874 9382 14876 9434
rect 14820 9380 14876 9382
rect 14924 9434 14980 9436
rect 14924 9382 14926 9434
rect 14926 9382 14978 9434
rect 14978 9382 14980 9434
rect 14924 9380 14980 9382
rect 15028 9434 15084 9436
rect 15028 9382 15030 9434
rect 15030 9382 15082 9434
rect 15082 9382 15084 9434
rect 15028 9380 15084 9382
rect 16828 9884 16884 9940
rect 18222 10218 18278 10220
rect 18222 10166 18224 10218
rect 18224 10166 18276 10218
rect 18276 10166 18278 10218
rect 18222 10164 18278 10166
rect 18326 10218 18382 10220
rect 18326 10166 18328 10218
rect 18328 10166 18380 10218
rect 18380 10166 18382 10218
rect 18326 10164 18382 10166
rect 18430 10218 18486 10220
rect 18430 10166 18432 10218
rect 18432 10166 18484 10218
rect 18484 10166 18486 10218
rect 18430 10164 18486 10166
rect 17276 9772 17332 9828
rect 17948 9884 18004 9940
rect 18956 11228 19012 11284
rect 19292 11506 19348 11508
rect 19292 11454 19294 11506
rect 19294 11454 19346 11506
rect 19346 11454 19348 11506
rect 19292 11452 19348 11454
rect 20300 11282 20356 11284
rect 20300 11230 20302 11282
rect 20302 11230 20354 11282
rect 20354 11230 20356 11282
rect 20300 11228 20356 11230
rect 19068 10780 19124 10836
rect 20188 10834 20244 10836
rect 20188 10782 20190 10834
rect 20190 10782 20242 10834
rect 20242 10782 20244 10834
rect 20188 10780 20244 10782
rect 18732 9884 18788 9940
rect 19180 9938 19236 9940
rect 19180 9886 19182 9938
rect 19182 9886 19234 9938
rect 19234 9886 19236 9938
rect 19180 9884 19236 9886
rect 19964 9826 20020 9828
rect 19964 9774 19966 9826
rect 19966 9774 20018 9826
rect 20018 9774 20020 9826
rect 19964 9772 20020 9774
rect 18396 9602 18452 9604
rect 18396 9550 18398 9602
rect 18398 9550 18450 9602
rect 18450 9550 18452 9602
rect 18396 9548 18452 9550
rect 19292 9602 19348 9604
rect 19292 9550 19294 9602
rect 19294 9550 19346 9602
rect 19346 9550 19348 9602
rect 19292 9548 19348 9550
rect 15932 8316 15988 8372
rect 13356 8092 13412 8148
rect 15484 8146 15540 8148
rect 15484 8094 15486 8146
rect 15486 8094 15538 8146
rect 15538 8094 15540 8146
rect 15484 8092 15540 8094
rect 18222 8650 18278 8652
rect 18222 8598 18224 8650
rect 18224 8598 18276 8650
rect 18276 8598 18278 8650
rect 18222 8596 18278 8598
rect 18326 8650 18382 8652
rect 18326 8598 18328 8650
rect 18328 8598 18380 8650
rect 18380 8598 18382 8650
rect 18326 8596 18382 8598
rect 18430 8650 18486 8652
rect 18430 8598 18432 8650
rect 18432 8598 18484 8650
rect 18484 8598 18486 8650
rect 18430 8596 18486 8598
rect 17612 8370 17668 8372
rect 17612 8318 17614 8370
rect 17614 8318 17666 8370
rect 17666 8318 17668 8370
rect 17612 8316 17668 8318
rect 16940 8092 16996 8148
rect 18620 8146 18676 8148
rect 18620 8094 18622 8146
rect 18622 8094 18674 8146
rect 18674 8094 18676 8146
rect 18620 8092 18676 8094
rect 2940 7644 2996 7700
rect 3836 7644 3892 7700
rect 2044 7420 2100 7476
rect 1932 6748 1988 6804
rect 2940 6748 2996 6804
rect 2044 6578 2100 6580
rect 2044 6526 2046 6578
rect 2046 6526 2098 6578
rect 2098 6526 2100 6578
rect 2044 6524 2100 6526
rect 1708 6076 1764 6132
rect 2492 6076 2548 6132
rect 1932 5404 1988 5460
rect 2044 5628 2100 5684
rect 8016 7866 8072 7868
rect 8016 7814 8018 7866
rect 8018 7814 8070 7866
rect 8070 7814 8072 7866
rect 8016 7812 8072 7814
rect 8120 7866 8176 7868
rect 8120 7814 8122 7866
rect 8122 7814 8174 7866
rect 8174 7814 8176 7866
rect 8120 7812 8176 7814
rect 8224 7866 8280 7868
rect 8224 7814 8226 7866
rect 8226 7814 8278 7866
rect 8278 7814 8280 7866
rect 8224 7812 8280 7814
rect 14820 7866 14876 7868
rect 14820 7814 14822 7866
rect 14822 7814 14874 7866
rect 14874 7814 14876 7866
rect 14820 7812 14876 7814
rect 14924 7866 14980 7868
rect 14924 7814 14926 7866
rect 14926 7814 14978 7866
rect 14978 7814 14980 7866
rect 14924 7812 14980 7814
rect 15028 7866 15084 7868
rect 15028 7814 15030 7866
rect 15030 7814 15082 7866
rect 15082 7814 15084 7866
rect 15028 7812 15084 7814
rect 23772 18172 23828 18228
rect 23212 16044 23268 16100
rect 23324 16716 23380 16772
rect 25026 22762 25082 22764
rect 25026 22710 25028 22762
rect 25028 22710 25080 22762
rect 25080 22710 25082 22762
rect 25026 22708 25082 22710
rect 25130 22762 25186 22764
rect 25130 22710 25132 22762
rect 25132 22710 25184 22762
rect 25184 22710 25186 22762
rect 25130 22708 25186 22710
rect 25234 22762 25290 22764
rect 25234 22710 25236 22762
rect 25236 22710 25288 22762
rect 25288 22710 25290 22762
rect 25234 22708 25290 22710
rect 26124 23436 26180 23492
rect 26236 23324 26292 23380
rect 27580 26236 27636 26292
rect 27468 24780 27524 24836
rect 26908 24722 26964 24724
rect 26908 24670 26910 24722
rect 26910 24670 26962 24722
rect 26962 24670 26964 24722
rect 26908 24668 26964 24670
rect 26908 23436 26964 23492
rect 25564 22540 25620 22596
rect 25452 21756 25508 21812
rect 25026 21194 25082 21196
rect 25026 21142 25028 21194
rect 25028 21142 25080 21194
rect 25080 21142 25082 21194
rect 25026 21140 25082 21142
rect 25130 21194 25186 21196
rect 25130 21142 25132 21194
rect 25132 21142 25184 21194
rect 25184 21142 25186 21194
rect 25130 21140 25186 21142
rect 25234 21194 25290 21196
rect 25234 21142 25236 21194
rect 25236 21142 25288 21194
rect 25288 21142 25290 21194
rect 25234 21140 25290 21142
rect 26124 23266 26180 23268
rect 26124 23214 26126 23266
rect 26126 23214 26178 23266
rect 26178 23214 26180 23266
rect 26124 23212 26180 23214
rect 26796 22876 26852 22932
rect 26460 22258 26516 22260
rect 26460 22206 26462 22258
rect 26462 22206 26514 22258
rect 26514 22206 26516 22258
rect 26460 22204 26516 22206
rect 27132 23378 27188 23380
rect 27132 23326 27134 23378
rect 27134 23326 27186 23378
rect 27186 23326 27188 23378
rect 27132 23324 27188 23326
rect 27692 25564 27748 25620
rect 27692 24892 27748 24948
rect 28140 27580 28196 27636
rect 28428 26682 28484 26684
rect 28428 26630 28430 26682
rect 28430 26630 28482 26682
rect 28482 26630 28484 26682
rect 28428 26628 28484 26630
rect 28532 26682 28588 26684
rect 28532 26630 28534 26682
rect 28534 26630 28586 26682
rect 28586 26630 28588 26682
rect 28532 26628 28588 26630
rect 28636 26682 28692 26684
rect 28636 26630 28638 26682
rect 28638 26630 28690 26682
rect 28690 26630 28692 26682
rect 28636 26628 28692 26630
rect 28140 24780 28196 24836
rect 28428 25114 28484 25116
rect 28428 25062 28430 25114
rect 28430 25062 28482 25114
rect 28482 25062 28484 25114
rect 28428 25060 28484 25062
rect 28532 25114 28588 25116
rect 28532 25062 28534 25114
rect 28534 25062 28586 25114
rect 28586 25062 28588 25114
rect 28532 25060 28588 25062
rect 28636 25114 28692 25116
rect 28636 25062 28638 25114
rect 28638 25062 28690 25114
rect 28690 25062 28692 25114
rect 28636 25060 28692 25062
rect 28252 24220 28308 24276
rect 27580 23660 27636 23716
rect 27468 22258 27524 22260
rect 27468 22206 27470 22258
rect 27470 22206 27522 22258
rect 27522 22206 27524 22258
rect 27468 22204 27524 22206
rect 27804 23100 27860 23156
rect 27804 22540 27860 22596
rect 28428 23546 28484 23548
rect 28428 23494 28430 23546
rect 28430 23494 28482 23546
rect 28482 23494 28484 23546
rect 28428 23492 28484 23494
rect 28532 23546 28588 23548
rect 28532 23494 28534 23546
rect 28534 23494 28586 23546
rect 28586 23494 28588 23546
rect 28532 23492 28588 23494
rect 28636 23546 28692 23548
rect 28636 23494 28638 23546
rect 28638 23494 28690 23546
rect 28690 23494 28692 23546
rect 28636 23492 28692 23494
rect 27804 21810 27860 21812
rect 27804 21758 27806 21810
rect 27806 21758 27858 21810
rect 27858 21758 27860 21810
rect 27804 21756 27860 21758
rect 28428 21978 28484 21980
rect 28428 21926 28430 21978
rect 28430 21926 28482 21978
rect 28482 21926 28484 21978
rect 28428 21924 28484 21926
rect 28532 21978 28588 21980
rect 28532 21926 28534 21978
rect 28534 21926 28586 21978
rect 28586 21926 28588 21978
rect 28532 21924 28588 21926
rect 28636 21978 28692 21980
rect 28636 21926 28638 21978
rect 28638 21926 28690 21978
rect 28690 21926 28692 21978
rect 28636 21924 28692 21926
rect 28028 21532 28084 21588
rect 27132 21474 27188 21476
rect 27132 21422 27134 21474
rect 27134 21422 27186 21474
rect 27186 21422 27188 21474
rect 27132 21420 27188 21422
rect 28140 21420 28196 21476
rect 28140 20860 28196 20916
rect 25788 20748 25844 20804
rect 26908 20802 26964 20804
rect 26908 20750 26910 20802
rect 26910 20750 26962 20802
rect 26962 20750 26964 20802
rect 26908 20748 26964 20750
rect 28428 20410 28484 20412
rect 28428 20358 28430 20410
rect 28430 20358 28482 20410
rect 28482 20358 28484 20410
rect 28428 20356 28484 20358
rect 28532 20410 28588 20412
rect 28532 20358 28534 20410
rect 28534 20358 28586 20410
rect 28586 20358 28588 20410
rect 28532 20356 28588 20358
rect 28636 20410 28692 20412
rect 28636 20358 28638 20410
rect 28638 20358 28690 20410
rect 28690 20358 28692 20410
rect 28636 20356 28692 20358
rect 28028 20188 28084 20244
rect 24892 19964 24948 20020
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 25026 19626 25082 19628
rect 25026 19574 25028 19626
rect 25028 19574 25080 19626
rect 25080 19574 25082 19626
rect 25026 19572 25082 19574
rect 25130 19626 25186 19628
rect 25130 19574 25132 19626
rect 25132 19574 25184 19626
rect 25184 19574 25186 19626
rect 25130 19572 25186 19574
rect 25234 19626 25290 19628
rect 25234 19574 25236 19626
rect 25236 19574 25288 19626
rect 25288 19574 25290 19626
rect 25234 19572 25290 19574
rect 28028 19516 28084 19572
rect 24780 19068 24836 19124
rect 23884 17612 23940 17668
rect 24556 18172 24612 18228
rect 24332 17724 24388 17780
rect 26236 18338 26292 18340
rect 26236 18286 26238 18338
rect 26238 18286 26290 18338
rect 26290 18286 26292 18338
rect 26236 18284 26292 18286
rect 26124 18172 26180 18228
rect 27244 18396 27300 18452
rect 25026 18058 25082 18060
rect 25026 18006 25028 18058
rect 25028 18006 25080 18058
rect 25080 18006 25082 18058
rect 25026 18004 25082 18006
rect 25130 18058 25186 18060
rect 25130 18006 25132 18058
rect 25132 18006 25184 18058
rect 25184 18006 25186 18058
rect 25130 18004 25186 18006
rect 25234 18058 25290 18060
rect 25234 18006 25236 18058
rect 25236 18006 25288 18058
rect 25288 18006 25290 18058
rect 25234 18004 25290 18006
rect 26124 17778 26180 17780
rect 26124 17726 26126 17778
rect 26126 17726 26178 17778
rect 26178 17726 26180 17778
rect 26124 17724 26180 17726
rect 26684 17612 26740 17668
rect 24892 17442 24948 17444
rect 24892 17390 24894 17442
rect 24894 17390 24946 17442
rect 24946 17390 24948 17442
rect 24892 17388 24948 17390
rect 26236 16770 26292 16772
rect 26236 16718 26238 16770
rect 26238 16718 26290 16770
rect 26290 16718 26292 16770
rect 26236 16716 26292 16718
rect 25026 16490 25082 16492
rect 25026 16438 25028 16490
rect 25028 16438 25080 16490
rect 25080 16438 25082 16490
rect 25026 16436 25082 16438
rect 25130 16490 25186 16492
rect 25130 16438 25132 16490
rect 25132 16438 25184 16490
rect 25184 16438 25186 16490
rect 25130 16436 25186 16438
rect 25234 16490 25290 16492
rect 25234 16438 25236 16490
rect 25236 16438 25288 16490
rect 25288 16438 25290 16490
rect 25234 16436 25290 16438
rect 27244 17388 27300 17444
rect 24668 16098 24724 16100
rect 24668 16046 24670 16098
rect 24670 16046 24722 16098
rect 24722 16046 24724 16098
rect 24668 16044 24724 16046
rect 26348 15932 26404 15988
rect 23548 15260 23604 15316
rect 24332 15314 24388 15316
rect 24332 15262 24334 15314
rect 24334 15262 24386 15314
rect 24386 15262 24388 15314
rect 24332 15260 24388 15262
rect 25228 15260 25284 15316
rect 25676 15314 25732 15316
rect 25676 15262 25678 15314
rect 25678 15262 25730 15314
rect 25730 15262 25732 15314
rect 25676 15260 25732 15262
rect 22092 14252 22148 14308
rect 21624 14138 21680 14140
rect 21624 14086 21626 14138
rect 21626 14086 21678 14138
rect 21678 14086 21680 14138
rect 21624 14084 21680 14086
rect 21728 14138 21784 14140
rect 21728 14086 21730 14138
rect 21730 14086 21782 14138
rect 21782 14086 21784 14138
rect 21728 14084 21784 14086
rect 21832 14138 21888 14140
rect 21832 14086 21834 14138
rect 21834 14086 21886 14138
rect 21886 14086 21888 14138
rect 21832 14084 21888 14086
rect 21308 13858 21364 13860
rect 21308 13806 21310 13858
rect 21310 13806 21362 13858
rect 21362 13806 21364 13858
rect 21308 13804 21364 13806
rect 21624 12570 21680 12572
rect 21624 12518 21626 12570
rect 21626 12518 21678 12570
rect 21678 12518 21680 12570
rect 21624 12516 21680 12518
rect 21728 12570 21784 12572
rect 21728 12518 21730 12570
rect 21730 12518 21782 12570
rect 21782 12518 21784 12570
rect 21728 12516 21784 12518
rect 21832 12570 21888 12572
rect 21832 12518 21834 12570
rect 21834 12518 21886 12570
rect 21886 12518 21888 12570
rect 21832 12516 21888 12518
rect 21420 12012 21476 12068
rect 25026 14922 25082 14924
rect 25026 14870 25028 14922
rect 25028 14870 25080 14922
rect 25080 14870 25082 14922
rect 25026 14868 25082 14870
rect 25130 14922 25186 14924
rect 25130 14870 25132 14922
rect 25132 14870 25184 14922
rect 25184 14870 25186 14922
rect 25130 14868 25186 14870
rect 25234 14922 25290 14924
rect 25234 14870 25236 14922
rect 25236 14870 25288 14922
rect 25288 14870 25290 14922
rect 25234 14868 25290 14870
rect 27804 19122 27860 19124
rect 27804 19070 27806 19122
rect 27806 19070 27858 19122
rect 27858 19070 27860 19122
rect 27804 19068 27860 19070
rect 28428 18842 28484 18844
rect 28428 18790 28430 18842
rect 28430 18790 28482 18842
rect 28482 18790 28484 18842
rect 28428 18788 28484 18790
rect 28532 18842 28588 18844
rect 28532 18790 28534 18842
rect 28534 18790 28586 18842
rect 28586 18790 28588 18842
rect 28532 18788 28588 18790
rect 28636 18842 28692 18844
rect 28636 18790 28638 18842
rect 28638 18790 28690 18842
rect 28690 18790 28692 18842
rect 28636 18788 28692 18790
rect 28252 18674 28308 18676
rect 28252 18622 28254 18674
rect 28254 18622 28306 18674
rect 28306 18622 28308 18674
rect 28252 18620 28308 18622
rect 27804 17500 27860 17556
rect 27692 15986 27748 15988
rect 27692 15934 27694 15986
rect 27694 15934 27746 15986
rect 27746 15934 27748 15986
rect 27692 15932 27748 15934
rect 28428 17274 28484 17276
rect 28428 17222 28430 17274
rect 28430 17222 28482 17274
rect 28482 17222 28484 17274
rect 28428 17220 28484 17222
rect 28532 17274 28588 17276
rect 28532 17222 28534 17274
rect 28534 17222 28586 17274
rect 28586 17222 28588 17274
rect 28532 17220 28588 17222
rect 28636 17274 28692 17276
rect 28636 17222 28638 17274
rect 28638 17222 28690 17274
rect 28690 17222 28692 17274
rect 28636 17220 28692 17222
rect 28140 16828 28196 16884
rect 26908 15148 26964 15204
rect 23436 14252 23492 14308
rect 22764 13858 22820 13860
rect 22764 13806 22766 13858
rect 22766 13806 22818 13858
rect 22818 13806 22820 13858
rect 22764 13804 22820 13806
rect 25026 13354 25082 13356
rect 25026 13302 25028 13354
rect 25028 13302 25080 13354
rect 25080 13302 25082 13354
rect 25026 13300 25082 13302
rect 25130 13354 25186 13356
rect 25130 13302 25132 13354
rect 25132 13302 25184 13354
rect 25184 13302 25186 13354
rect 25130 13300 25186 13302
rect 25234 13354 25290 13356
rect 25234 13302 25236 13354
rect 25236 13302 25288 13354
rect 25288 13302 25290 13354
rect 25234 13300 25290 13302
rect 22316 12684 22372 12740
rect 22652 12460 22708 12516
rect 24108 12684 24164 12740
rect 22204 12012 22260 12068
rect 25116 12738 25172 12740
rect 25116 12686 25118 12738
rect 25118 12686 25170 12738
rect 25170 12686 25172 12738
rect 25116 12684 25172 12686
rect 28428 15706 28484 15708
rect 28428 15654 28430 15706
rect 28430 15654 28482 15706
rect 28482 15654 28484 15706
rect 28428 15652 28484 15654
rect 28532 15706 28588 15708
rect 28532 15654 28534 15706
rect 28534 15654 28586 15706
rect 28586 15654 28588 15706
rect 28532 15652 28588 15654
rect 28636 15706 28692 15708
rect 28636 15654 28638 15706
rect 28638 15654 28690 15706
rect 28690 15654 28692 15706
rect 28636 15652 28692 15654
rect 28428 14138 28484 14140
rect 28428 14086 28430 14138
rect 28430 14086 28482 14138
rect 28482 14086 28484 14138
rect 28428 14084 28484 14086
rect 28532 14138 28588 14140
rect 28532 14086 28534 14138
rect 28534 14086 28586 14138
rect 28586 14086 28588 14138
rect 28532 14084 28588 14086
rect 28636 14138 28692 14140
rect 28636 14086 28638 14138
rect 28638 14086 28690 14138
rect 28690 14086 28692 14138
rect 28636 14084 28692 14086
rect 24444 12066 24500 12068
rect 24444 12014 24446 12066
rect 24446 12014 24498 12066
rect 24498 12014 24500 12066
rect 24444 12012 24500 12014
rect 24892 11788 24948 11844
rect 25026 11786 25082 11788
rect 25026 11734 25028 11786
rect 25028 11734 25080 11786
rect 25080 11734 25082 11786
rect 25026 11732 25082 11734
rect 25130 11786 25186 11788
rect 25130 11734 25132 11786
rect 25132 11734 25184 11786
rect 25184 11734 25186 11786
rect 25130 11732 25186 11734
rect 25234 11786 25290 11788
rect 25234 11734 25236 11786
rect 25236 11734 25288 11786
rect 25288 11734 25290 11786
rect 25234 11732 25290 11734
rect 21624 11002 21680 11004
rect 21624 10950 21626 11002
rect 21626 10950 21678 11002
rect 21678 10950 21680 11002
rect 21624 10948 21680 10950
rect 21728 11002 21784 11004
rect 21728 10950 21730 11002
rect 21730 10950 21782 11002
rect 21782 10950 21784 11002
rect 21728 10948 21784 10950
rect 21832 11002 21888 11004
rect 21832 10950 21834 11002
rect 21834 10950 21886 11002
rect 21886 10950 21888 11002
rect 21832 10948 21888 10950
rect 25676 11228 25732 11284
rect 26012 12738 26068 12740
rect 26012 12686 26014 12738
rect 26014 12686 26066 12738
rect 26066 12686 26068 12738
rect 26012 12684 26068 12686
rect 28428 12570 28484 12572
rect 26236 12460 26292 12516
rect 28428 12518 28430 12570
rect 28430 12518 28482 12570
rect 28482 12518 28484 12570
rect 28428 12516 28484 12518
rect 28532 12570 28588 12572
rect 28532 12518 28534 12570
rect 28534 12518 28586 12570
rect 28586 12518 28588 12570
rect 28532 12516 28588 12518
rect 28636 12570 28692 12572
rect 28636 12518 28638 12570
rect 28638 12518 28690 12570
rect 28690 12518 28692 12570
rect 28636 12516 28692 12518
rect 27244 11900 27300 11956
rect 20972 10386 21028 10388
rect 20972 10334 20974 10386
rect 20974 10334 21026 10386
rect 21026 10334 21028 10386
rect 20972 10332 21028 10334
rect 21756 10444 21812 10500
rect 23772 9996 23828 10052
rect 21308 9884 21364 9940
rect 21868 9826 21924 9828
rect 21868 9774 21870 9826
rect 21870 9774 21922 9826
rect 21922 9774 21924 9826
rect 21868 9772 21924 9774
rect 21624 9434 21680 9436
rect 21624 9382 21626 9434
rect 21626 9382 21678 9434
rect 21678 9382 21680 9434
rect 21624 9380 21680 9382
rect 21728 9434 21784 9436
rect 21728 9382 21730 9434
rect 21730 9382 21782 9434
rect 21782 9382 21784 9434
rect 21728 9380 21784 9382
rect 21832 9434 21888 9436
rect 21832 9382 21834 9434
rect 21834 9382 21886 9434
rect 21886 9382 21888 9434
rect 21832 9380 21888 9382
rect 20860 9212 20916 9268
rect 21644 9266 21700 9268
rect 21644 9214 21646 9266
rect 21646 9214 21698 9266
rect 21698 9214 21700 9266
rect 21644 9212 21700 9214
rect 22540 8876 22596 8932
rect 22988 9772 23044 9828
rect 23548 9266 23604 9268
rect 23548 9214 23550 9266
rect 23550 9214 23602 9266
rect 23602 9214 23604 9266
rect 23548 9212 23604 9214
rect 21624 7866 21680 7868
rect 21624 7814 21626 7866
rect 21626 7814 21678 7866
rect 21678 7814 21680 7866
rect 21624 7812 21680 7814
rect 21728 7866 21784 7868
rect 21728 7814 21730 7866
rect 21730 7814 21782 7866
rect 21782 7814 21784 7866
rect 21728 7812 21784 7814
rect 21832 7866 21888 7868
rect 21832 7814 21834 7866
rect 21834 7814 21886 7866
rect 21886 7814 21888 7866
rect 21832 7812 21888 7814
rect 22092 7586 22148 7588
rect 22092 7534 22094 7586
rect 22094 7534 22146 7586
rect 22146 7534 22148 7586
rect 22092 7532 22148 7534
rect 4614 7082 4670 7084
rect 4614 7030 4616 7082
rect 4616 7030 4668 7082
rect 4668 7030 4670 7082
rect 4614 7028 4670 7030
rect 4718 7082 4774 7084
rect 4718 7030 4720 7082
rect 4720 7030 4772 7082
rect 4772 7030 4774 7082
rect 4718 7028 4774 7030
rect 4822 7082 4878 7084
rect 4822 7030 4824 7082
rect 4824 7030 4876 7082
rect 4876 7030 4878 7082
rect 4822 7028 4878 7030
rect 11418 7082 11474 7084
rect 11418 7030 11420 7082
rect 11420 7030 11472 7082
rect 11472 7030 11474 7082
rect 11418 7028 11474 7030
rect 11522 7082 11578 7084
rect 11522 7030 11524 7082
rect 11524 7030 11576 7082
rect 11576 7030 11578 7082
rect 11522 7028 11578 7030
rect 11626 7082 11682 7084
rect 11626 7030 11628 7082
rect 11628 7030 11680 7082
rect 11680 7030 11682 7082
rect 11626 7028 11682 7030
rect 18222 7082 18278 7084
rect 18222 7030 18224 7082
rect 18224 7030 18276 7082
rect 18276 7030 18278 7082
rect 18222 7028 18278 7030
rect 18326 7082 18382 7084
rect 18326 7030 18328 7082
rect 18328 7030 18380 7082
rect 18380 7030 18382 7082
rect 18326 7028 18382 7030
rect 18430 7082 18486 7084
rect 18430 7030 18432 7082
rect 18432 7030 18484 7082
rect 18484 7030 18486 7082
rect 18430 7028 18486 7030
rect 4172 6748 4228 6804
rect 4172 6578 4228 6580
rect 4172 6526 4174 6578
rect 4174 6526 4226 6578
rect 4226 6526 4228 6578
rect 4172 6524 4228 6526
rect 23772 9212 23828 9268
rect 23100 7532 23156 7588
rect 24332 9212 24388 9268
rect 25026 10218 25082 10220
rect 25026 10166 25028 10218
rect 25028 10166 25080 10218
rect 25080 10166 25082 10218
rect 25026 10164 25082 10166
rect 25130 10218 25186 10220
rect 25130 10166 25132 10218
rect 25132 10166 25184 10218
rect 25184 10166 25186 10218
rect 25130 10164 25186 10166
rect 25234 10218 25290 10220
rect 25234 10166 25236 10218
rect 25236 10166 25288 10218
rect 25288 10166 25290 10218
rect 25234 10164 25290 10166
rect 25564 10108 25620 10164
rect 26236 10498 26292 10500
rect 26236 10446 26238 10498
rect 26238 10446 26290 10498
rect 26290 10446 26292 10498
rect 26236 10444 26292 10446
rect 27692 11282 27748 11284
rect 27692 11230 27694 11282
rect 27694 11230 27746 11282
rect 27746 11230 27748 11282
rect 27692 11228 27748 11230
rect 28428 11002 28484 11004
rect 28428 10950 28430 11002
rect 28430 10950 28482 11002
rect 28482 10950 28484 11002
rect 28428 10948 28484 10950
rect 28532 11002 28588 11004
rect 28532 10950 28534 11002
rect 28534 10950 28586 11002
rect 28586 10950 28588 11002
rect 28532 10948 28588 10950
rect 28636 11002 28692 11004
rect 28636 10950 28638 11002
rect 28638 10950 28690 11002
rect 28690 10950 28692 11002
rect 28636 10948 28692 10950
rect 26684 9996 26740 10052
rect 26908 10332 26964 10388
rect 27244 10108 27300 10164
rect 27692 10050 27748 10052
rect 27692 9998 27694 10050
rect 27694 9998 27746 10050
rect 27746 9998 27748 10050
rect 27692 9996 27748 9998
rect 25452 9266 25508 9268
rect 25452 9214 25454 9266
rect 25454 9214 25506 9266
rect 25506 9214 25508 9266
rect 25452 9212 25508 9214
rect 25026 8650 25082 8652
rect 25026 8598 25028 8650
rect 25028 8598 25080 8650
rect 25080 8598 25082 8650
rect 25026 8596 25082 8598
rect 25130 8650 25186 8652
rect 25130 8598 25132 8650
rect 25132 8598 25184 8650
rect 25184 8598 25186 8650
rect 25130 8596 25186 8598
rect 25234 8650 25290 8652
rect 25234 8598 25236 8650
rect 25236 8598 25288 8650
rect 25288 8598 25290 8650
rect 25234 8596 25290 8598
rect 28428 9434 28484 9436
rect 28428 9382 28430 9434
rect 28430 9382 28482 9434
rect 28482 9382 28484 9434
rect 28428 9380 28484 9382
rect 28532 9434 28588 9436
rect 28532 9382 28534 9434
rect 28534 9382 28586 9434
rect 28586 9382 28588 9434
rect 28532 9380 28588 9382
rect 28636 9434 28692 9436
rect 28636 9382 28638 9434
rect 28638 9382 28690 9434
rect 28690 9382 28692 9434
rect 28636 9380 28692 9382
rect 26236 8930 26292 8932
rect 26236 8878 26238 8930
rect 26238 8878 26290 8930
rect 26290 8878 26292 8930
rect 26236 8876 26292 8878
rect 27692 8370 27748 8372
rect 27692 8318 27694 8370
rect 27694 8318 27746 8370
rect 27746 8318 27748 8370
rect 27692 8316 27748 8318
rect 23772 6860 23828 6916
rect 22988 6690 23044 6692
rect 22988 6638 22990 6690
rect 22990 6638 23042 6690
rect 23042 6638 23044 6690
rect 22988 6636 23044 6638
rect 8016 6298 8072 6300
rect 8016 6246 8018 6298
rect 8018 6246 8070 6298
rect 8070 6246 8072 6298
rect 8016 6244 8072 6246
rect 8120 6298 8176 6300
rect 8120 6246 8122 6298
rect 8122 6246 8174 6298
rect 8174 6246 8176 6298
rect 8120 6244 8176 6246
rect 8224 6298 8280 6300
rect 8224 6246 8226 6298
rect 8226 6246 8278 6298
rect 8278 6246 8280 6298
rect 8224 6244 8280 6246
rect 14820 6298 14876 6300
rect 14820 6246 14822 6298
rect 14822 6246 14874 6298
rect 14874 6246 14876 6298
rect 14820 6244 14876 6246
rect 14924 6298 14980 6300
rect 14924 6246 14926 6298
rect 14926 6246 14978 6298
rect 14978 6246 14980 6298
rect 14924 6244 14980 6246
rect 15028 6298 15084 6300
rect 15028 6246 15030 6298
rect 15030 6246 15082 6298
rect 15082 6246 15084 6298
rect 15028 6244 15084 6246
rect 21624 6298 21680 6300
rect 21624 6246 21626 6298
rect 21626 6246 21678 6298
rect 21678 6246 21680 6298
rect 21624 6244 21680 6246
rect 21728 6298 21784 6300
rect 21728 6246 21730 6298
rect 21730 6246 21782 6298
rect 21782 6246 21784 6298
rect 21728 6244 21784 6246
rect 21832 6298 21888 6300
rect 21832 6246 21834 6298
rect 21834 6246 21886 6298
rect 21886 6246 21888 6298
rect 21832 6244 21888 6246
rect 3388 5628 3444 5684
rect 9212 5852 9268 5908
rect 4614 5514 4670 5516
rect 4614 5462 4616 5514
rect 4616 5462 4668 5514
rect 4668 5462 4670 5514
rect 4614 5460 4670 5462
rect 4718 5514 4774 5516
rect 4718 5462 4720 5514
rect 4720 5462 4772 5514
rect 4772 5462 4774 5514
rect 4718 5460 4774 5462
rect 4822 5514 4878 5516
rect 4822 5462 4824 5514
rect 4824 5462 4876 5514
rect 4876 5462 4878 5514
rect 4822 5460 4878 5462
rect 1708 4732 1764 4788
rect 2492 4732 2548 4788
rect 8016 4730 8072 4732
rect 8016 4678 8018 4730
rect 8018 4678 8070 4730
rect 8070 4678 8072 4730
rect 8016 4676 8072 4678
rect 8120 4730 8176 4732
rect 8120 4678 8122 4730
rect 8122 4678 8174 4730
rect 8174 4678 8176 4730
rect 8120 4676 8176 4678
rect 8224 4730 8280 4732
rect 8224 4678 8226 4730
rect 8226 4678 8278 4730
rect 8278 4678 8280 4730
rect 8224 4676 8280 4678
rect 4614 3946 4670 3948
rect 4614 3894 4616 3946
rect 4616 3894 4668 3946
rect 4668 3894 4670 3946
rect 4614 3892 4670 3894
rect 4718 3946 4774 3948
rect 4718 3894 4720 3946
rect 4720 3894 4772 3946
rect 4772 3894 4774 3946
rect 4718 3892 4774 3894
rect 4822 3946 4878 3948
rect 4822 3894 4824 3946
rect 4824 3894 4876 3946
rect 4876 3894 4878 3946
rect 4822 3892 4878 3894
rect 8016 3162 8072 3164
rect 8016 3110 8018 3162
rect 8018 3110 8070 3162
rect 8070 3110 8072 3162
rect 8016 3108 8072 3110
rect 8120 3162 8176 3164
rect 8120 3110 8122 3162
rect 8122 3110 8174 3162
rect 8174 3110 8176 3162
rect 8120 3108 8176 3110
rect 8224 3162 8280 3164
rect 8224 3110 8226 3162
rect 8226 3110 8278 3162
rect 8278 3110 8280 3162
rect 8224 3108 8280 3110
rect 9996 5906 10052 5908
rect 9996 5854 9998 5906
rect 9998 5854 10050 5906
rect 10050 5854 10052 5906
rect 9996 5852 10052 5854
rect 23324 5852 23380 5908
rect 11418 5514 11474 5516
rect 11418 5462 11420 5514
rect 11420 5462 11472 5514
rect 11472 5462 11474 5514
rect 11418 5460 11474 5462
rect 11522 5514 11578 5516
rect 11522 5462 11524 5514
rect 11524 5462 11576 5514
rect 11576 5462 11578 5514
rect 11522 5460 11578 5462
rect 11626 5514 11682 5516
rect 11626 5462 11628 5514
rect 11628 5462 11680 5514
rect 11680 5462 11682 5514
rect 11626 5460 11682 5462
rect 18222 5514 18278 5516
rect 18222 5462 18224 5514
rect 18224 5462 18276 5514
rect 18276 5462 18278 5514
rect 18222 5460 18278 5462
rect 18326 5514 18382 5516
rect 18326 5462 18328 5514
rect 18328 5462 18380 5514
rect 18380 5462 18382 5514
rect 18326 5460 18382 5462
rect 18430 5514 18486 5516
rect 18430 5462 18432 5514
rect 18432 5462 18484 5514
rect 18484 5462 18486 5514
rect 18430 5460 18486 5462
rect 14820 4730 14876 4732
rect 11116 4620 11172 4676
rect 13132 4620 13188 4676
rect 14820 4678 14822 4730
rect 14822 4678 14874 4730
rect 14874 4678 14876 4730
rect 14820 4676 14876 4678
rect 14924 4730 14980 4732
rect 14924 4678 14926 4730
rect 14926 4678 14978 4730
rect 14978 4678 14980 4730
rect 14924 4676 14980 4678
rect 15028 4730 15084 4732
rect 15028 4678 15030 4730
rect 15030 4678 15082 4730
rect 15082 4678 15084 4730
rect 15028 4676 15084 4678
rect 10892 4508 10948 4564
rect 11900 4562 11956 4564
rect 11900 4510 11902 4562
rect 11902 4510 11954 4562
rect 11954 4510 11956 4562
rect 11900 4508 11956 4510
rect 11418 3946 11474 3948
rect 11418 3894 11420 3946
rect 11420 3894 11472 3946
rect 11472 3894 11474 3946
rect 11418 3892 11474 3894
rect 11522 3946 11578 3948
rect 11522 3894 11524 3946
rect 11524 3894 11576 3946
rect 11576 3894 11578 3946
rect 11522 3892 11578 3894
rect 11626 3946 11682 3948
rect 11626 3894 11628 3946
rect 11628 3894 11680 3946
rect 11680 3894 11682 3946
rect 11626 3892 11682 3894
rect 12124 3612 12180 3668
rect 18222 3946 18278 3948
rect 18222 3894 18224 3946
rect 18224 3894 18276 3946
rect 18276 3894 18278 3946
rect 18222 3892 18278 3894
rect 18326 3946 18382 3948
rect 18326 3894 18328 3946
rect 18328 3894 18380 3946
rect 18380 3894 18382 3946
rect 18326 3892 18382 3894
rect 18430 3946 18486 3948
rect 18430 3894 18432 3946
rect 18432 3894 18484 3946
rect 18484 3894 18486 3946
rect 18430 3892 18486 3894
rect 13580 3666 13636 3668
rect 13580 3614 13582 3666
rect 13582 3614 13634 3666
rect 13634 3614 13636 3666
rect 13580 3612 13636 3614
rect 21624 4730 21680 4732
rect 21624 4678 21626 4730
rect 21626 4678 21678 4730
rect 21678 4678 21680 4730
rect 21624 4676 21680 4678
rect 21728 4730 21784 4732
rect 21728 4678 21730 4730
rect 21730 4678 21782 4730
rect 21782 4678 21784 4730
rect 21728 4676 21784 4678
rect 21832 4730 21888 4732
rect 21832 4678 21834 4730
rect 21834 4678 21886 4730
rect 21886 4678 21888 4730
rect 21832 4676 21888 4678
rect 14820 3162 14876 3164
rect 14820 3110 14822 3162
rect 14822 3110 14874 3162
rect 14874 3110 14876 3162
rect 14820 3108 14876 3110
rect 14924 3162 14980 3164
rect 14924 3110 14926 3162
rect 14926 3110 14978 3162
rect 14978 3110 14980 3162
rect 14924 3108 14980 3110
rect 15028 3162 15084 3164
rect 15028 3110 15030 3162
rect 15030 3110 15082 3162
rect 15082 3110 15084 3162
rect 15028 3108 15084 3110
rect 21624 3162 21680 3164
rect 21624 3110 21626 3162
rect 21626 3110 21678 3162
rect 21678 3110 21680 3162
rect 21624 3108 21680 3110
rect 21728 3162 21784 3164
rect 21728 3110 21730 3162
rect 21730 3110 21782 3162
rect 21782 3110 21784 3162
rect 21728 3108 21784 3110
rect 21832 3162 21888 3164
rect 21832 3110 21834 3162
rect 21834 3110 21886 3162
rect 21886 3110 21888 3162
rect 21832 3108 21888 3110
rect 23884 6076 23940 6132
rect 25026 7082 25082 7084
rect 25026 7030 25028 7082
rect 25028 7030 25080 7082
rect 25080 7030 25082 7082
rect 25026 7028 25082 7030
rect 25130 7082 25186 7084
rect 25130 7030 25132 7082
rect 25132 7030 25184 7082
rect 25184 7030 25186 7082
rect 25130 7028 25186 7030
rect 25234 7082 25290 7084
rect 25234 7030 25236 7082
rect 25236 7030 25288 7082
rect 25288 7030 25290 7082
rect 25234 7028 25290 7030
rect 25676 6748 25732 6804
rect 25452 6130 25508 6132
rect 25452 6078 25454 6130
rect 25454 6078 25506 6130
rect 25506 6078 25508 6130
rect 25452 6076 25508 6078
rect 23996 6018 24052 6020
rect 23996 5966 23998 6018
rect 23998 5966 24050 6018
rect 24050 5966 24052 6018
rect 23996 5964 24052 5966
rect 24332 5906 24388 5908
rect 24332 5854 24334 5906
rect 24334 5854 24386 5906
rect 24386 5854 24388 5906
rect 24332 5852 24388 5854
rect 24108 5180 24164 5236
rect 23996 4956 24052 5012
rect 23100 2716 23156 2772
rect 24332 3388 24388 3444
rect 25026 5514 25082 5516
rect 25026 5462 25028 5514
rect 25028 5462 25080 5514
rect 25080 5462 25082 5514
rect 25026 5460 25082 5462
rect 25130 5514 25186 5516
rect 25130 5462 25132 5514
rect 25132 5462 25184 5514
rect 25184 5462 25186 5514
rect 25130 5460 25186 5462
rect 25234 5514 25290 5516
rect 25234 5462 25236 5514
rect 25236 5462 25288 5514
rect 25288 5462 25290 5514
rect 25234 5460 25290 5462
rect 24668 5068 24724 5124
rect 26796 6690 26852 6692
rect 26796 6638 26798 6690
rect 26798 6638 26850 6690
rect 26850 6638 26852 6690
rect 26796 6636 26852 6638
rect 27244 6748 27300 6804
rect 25676 5964 25732 6020
rect 25900 5180 25956 5236
rect 24892 4620 24948 4676
rect 25452 4844 25508 4900
rect 25026 3946 25082 3948
rect 25026 3894 25028 3946
rect 25028 3894 25080 3946
rect 25080 3894 25082 3946
rect 25026 3892 25082 3894
rect 25130 3946 25186 3948
rect 25130 3894 25132 3946
rect 25132 3894 25184 3946
rect 25184 3894 25186 3946
rect 25130 3892 25186 3894
rect 25234 3946 25290 3948
rect 25234 3894 25236 3946
rect 25236 3894 25288 3946
rect 25288 3894 25290 3946
rect 25234 3892 25290 3894
rect 25900 4620 25956 4676
rect 25788 4508 25844 4564
rect 25564 4450 25620 4452
rect 25564 4398 25566 4450
rect 25566 4398 25618 4450
rect 25618 4398 25620 4450
rect 25564 4396 25620 4398
rect 28140 8092 28196 8148
rect 27692 7420 27748 7476
rect 26908 5122 26964 5124
rect 26908 5070 26910 5122
rect 26910 5070 26962 5122
rect 26962 5070 26964 5122
rect 26908 5068 26964 5070
rect 27244 4956 27300 5012
rect 27356 5404 27412 5460
rect 26908 4562 26964 4564
rect 26908 4510 26910 4562
rect 26910 4510 26962 4562
rect 26962 4510 26964 4562
rect 26908 4508 26964 4510
rect 26460 4396 26516 4452
rect 27580 6748 27636 6804
rect 27804 6860 27860 6916
rect 28428 7866 28484 7868
rect 28428 7814 28430 7866
rect 28430 7814 28482 7866
rect 28482 7814 28484 7866
rect 28428 7812 28484 7814
rect 28532 7866 28588 7868
rect 28532 7814 28534 7866
rect 28534 7814 28586 7866
rect 28586 7814 28588 7866
rect 28532 7812 28588 7814
rect 28636 7866 28692 7868
rect 28636 7814 28638 7866
rect 28638 7814 28690 7866
rect 28690 7814 28692 7866
rect 28636 7812 28692 7814
rect 28428 6298 28484 6300
rect 28428 6246 28430 6298
rect 28430 6246 28482 6298
rect 28482 6246 28484 6298
rect 28428 6244 28484 6246
rect 28532 6298 28588 6300
rect 28532 6246 28534 6298
rect 28534 6246 28586 6298
rect 28586 6246 28588 6298
rect 28532 6244 28588 6246
rect 28636 6298 28692 6300
rect 28636 6246 28638 6298
rect 28638 6246 28690 6298
rect 28690 6246 28692 6298
rect 28636 6244 28692 6246
rect 27692 5852 27748 5908
rect 28428 4730 28484 4732
rect 28428 4678 28430 4730
rect 28430 4678 28482 4730
rect 28482 4678 28484 4730
rect 28428 4676 28484 4678
rect 28532 4730 28588 4732
rect 28532 4678 28534 4730
rect 28534 4678 28586 4730
rect 28586 4678 28588 4730
rect 28532 4676 28588 4678
rect 28636 4730 28692 4732
rect 28636 4678 28638 4730
rect 28638 4678 28690 4730
rect 28690 4678 28692 4730
rect 28636 4676 28692 4678
rect 27468 4060 27524 4116
rect 24892 3442 24948 3444
rect 24892 3390 24894 3442
rect 24894 3390 24946 3442
rect 24946 3390 24948 3442
rect 24892 3388 24948 3390
rect 28428 3162 28484 3164
rect 28428 3110 28430 3162
rect 28430 3110 28482 3162
rect 28482 3110 28484 3162
rect 28428 3108 28484 3110
rect 28532 3162 28588 3164
rect 28532 3110 28534 3162
rect 28534 3110 28586 3162
rect 28586 3110 28588 3162
rect 28532 3108 28588 3110
rect 28636 3162 28692 3164
rect 28636 3110 28638 3162
rect 28638 3110 28690 3162
rect 28690 3110 28692 3162
rect 28636 3108 28692 3110
rect 24668 2044 24724 2100
rect 23772 1372 23828 1428
<< metal3 >>
rect 29200 28980 30000 29008
rect 24434 28924 24444 28980
rect 24500 28924 30000 28980
rect 29200 28896 30000 28924
rect 0 28308 800 28336
rect 29200 28308 30000 28336
rect 0 28252 1820 28308
rect 1876 28252 1886 28308
rect 27794 28252 27804 28308
rect 27860 28252 30000 28308
rect 0 28224 800 28252
rect 29200 28224 30000 28252
rect 0 27636 800 27664
rect 29200 27636 30000 27664
rect 0 27580 3724 27636
rect 3780 27580 3790 27636
rect 28130 27580 28140 27636
rect 28196 27580 30000 27636
rect 0 27552 800 27580
rect 29200 27552 30000 27580
rect 0 26964 800 26992
rect 29200 26964 30000 26992
rect 0 26908 3388 26964
rect 3444 26908 3454 26964
rect 26114 26908 26124 26964
rect 26180 26908 30000 26964
rect 0 26880 800 26908
rect 29200 26880 30000 26908
rect 14802 26796 14812 26852
rect 14868 26796 15820 26852
rect 15876 26796 15886 26852
rect 8006 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8290 26684
rect 14810 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15094 26684
rect 21614 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21898 26684
rect 28418 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28702 26684
rect 12786 26460 12796 26516
rect 12852 26460 13580 26516
rect 13636 26460 13646 26516
rect 18162 26460 18172 26516
rect 18228 26460 19068 26516
rect 19124 26460 19134 26516
rect 8754 26348 8764 26404
rect 8820 26348 10108 26404
rect 10164 26348 10174 26404
rect 20402 26348 20412 26404
rect 20468 26348 21532 26404
rect 21588 26348 21598 26404
rect 0 26292 800 26320
rect 29200 26292 30000 26320
rect 0 26236 2044 26292
rect 2100 26236 2110 26292
rect 2930 26236 2940 26292
rect 2996 26236 3948 26292
rect 4004 26236 4014 26292
rect 6402 26236 6412 26292
rect 6468 26236 6972 26292
rect 7028 26236 7038 26292
rect 7858 26236 7868 26292
rect 7924 26236 8316 26292
rect 8372 26236 8382 26292
rect 20290 26236 20300 26292
rect 20356 26236 20972 26292
rect 21028 26236 21038 26292
rect 27570 26236 27580 26292
rect 27636 26236 30000 26292
rect 0 26208 800 26236
rect 29200 26208 30000 26236
rect 11442 26012 11452 26068
rect 11508 26012 12124 26068
rect 12180 26012 12190 26068
rect 4604 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4888 25900
rect 11408 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11692 25900
rect 18212 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18496 25900
rect 25016 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25300 25900
rect 22866 25676 22876 25732
rect 22932 25676 23548 25732
rect 23604 25676 23614 25732
rect 24210 25676 24220 25732
rect 24276 25676 25340 25732
rect 25396 25676 25406 25732
rect 0 25620 800 25648
rect 29200 25620 30000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 7410 25564 7420 25620
rect 7476 25564 11452 25620
rect 11508 25564 11518 25620
rect 27682 25564 27692 25620
rect 27748 25564 30000 25620
rect 0 25536 800 25564
rect 29200 25536 30000 25564
rect 1810 25452 1820 25508
rect 1876 25452 3276 25508
rect 3332 25452 3342 25508
rect 6066 25452 6076 25508
rect 6132 25452 10668 25508
rect 10724 25452 10734 25508
rect 15362 25452 15372 25508
rect 15428 25452 15932 25508
rect 15988 25452 15998 25508
rect 20850 25452 20860 25508
rect 20916 25452 21644 25508
rect 21700 25452 21710 25508
rect 5954 25340 5964 25396
rect 6020 25340 10780 25396
rect 10836 25340 10846 25396
rect 20738 25340 20748 25396
rect 20804 25340 23100 25396
rect 23156 25340 23166 25396
rect 2146 25228 2156 25284
rect 2212 25228 2222 25284
rect 2930 25228 2940 25284
rect 2996 25228 3500 25284
rect 3556 25228 3566 25284
rect 6738 25228 6748 25284
rect 6804 25228 9324 25284
rect 9380 25228 9390 25284
rect 10322 25228 10332 25284
rect 10388 25228 11676 25284
rect 11732 25228 11742 25284
rect 12114 25228 12124 25284
rect 12180 25228 15708 25284
rect 15764 25228 15774 25284
rect 19394 25228 19404 25284
rect 19460 25228 20636 25284
rect 20692 25228 20702 25284
rect 21196 25228 24668 25284
rect 24724 25228 24734 25284
rect 0 24948 800 24976
rect 2156 24948 2212 25228
rect 8006 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8290 25116
rect 14810 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15094 25116
rect 21196 25060 21252 25228
rect 21614 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21898 25116
rect 28418 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28702 25116
rect 21186 25004 21196 25060
rect 21252 25004 21262 25060
rect 29200 24948 30000 24976
rect 0 24892 2212 24948
rect 27682 24892 27692 24948
rect 27748 24892 30000 24948
rect 0 24864 800 24892
rect 29200 24864 30000 24892
rect 2930 24780 2940 24836
rect 2996 24780 4956 24836
rect 5012 24780 5022 24836
rect 27458 24780 27468 24836
rect 27524 24780 28140 24836
rect 28196 24780 28206 24836
rect 2706 24668 2716 24724
rect 2772 24668 4284 24724
rect 4340 24668 4350 24724
rect 25778 24668 25788 24724
rect 25844 24668 26908 24724
rect 26964 24668 26974 24724
rect 20962 24444 20972 24500
rect 21028 24444 22428 24500
rect 22484 24444 22494 24500
rect 24322 24444 24332 24500
rect 24388 24444 25340 24500
rect 25396 24444 25406 24500
rect 0 24276 800 24304
rect 4604 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4888 24332
rect 11408 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11692 24332
rect 18212 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18496 24332
rect 25016 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25300 24332
rect 29200 24276 30000 24304
rect 0 24220 2380 24276
rect 2436 24220 3164 24276
rect 3220 24220 3230 24276
rect 28242 24220 28252 24276
rect 28308 24220 30000 24276
rect 0 24192 800 24220
rect 29200 24192 30000 24220
rect 2258 23884 2268 23940
rect 2324 23884 4956 23940
rect 5012 23884 5022 23940
rect 7858 23884 7868 23940
rect 7924 23884 11340 23940
rect 11396 23884 11406 23940
rect 2034 23772 2044 23828
rect 2100 23772 5180 23828
rect 5236 23772 5246 23828
rect 11666 23772 11676 23828
rect 11732 23772 15260 23828
rect 15316 23772 15326 23828
rect 21634 23772 21644 23828
rect 21700 23772 24556 23828
rect 24612 23772 24622 23828
rect 2930 23660 2940 23716
rect 2996 23660 4732 23716
rect 4788 23660 4798 23716
rect 27570 23660 27580 23716
rect 27636 23660 28868 23716
rect 0 23604 800 23632
rect 28812 23604 28868 23660
rect 29200 23604 30000 23632
rect 0 23548 1708 23604
rect 1764 23548 1774 23604
rect 28812 23548 30000 23604
rect 0 23520 800 23548
rect 8006 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8290 23548
rect 14810 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15094 23548
rect 21614 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21898 23548
rect 28418 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28702 23548
rect 29200 23520 30000 23548
rect 26114 23436 26124 23492
rect 26180 23436 26908 23492
rect 26964 23436 26974 23492
rect 26226 23324 26236 23380
rect 26292 23324 27132 23380
rect 27188 23324 27198 23380
rect 24658 23212 24668 23268
rect 24724 23212 26124 23268
rect 26180 23212 26190 23268
rect 24098 23100 24108 23156
rect 24164 23100 27804 23156
rect 27860 23100 27870 23156
rect 0 22932 800 22960
rect 29200 22932 30000 22960
rect 0 22876 1708 22932
rect 1764 22876 2492 22932
rect 2548 22876 2558 22932
rect 26786 22876 26796 22932
rect 26852 22876 30000 22932
rect 0 22848 800 22876
rect 29200 22848 30000 22876
rect 4604 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4888 22764
rect 11408 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11692 22764
rect 18212 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18496 22764
rect 25016 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25300 22764
rect 25554 22540 25564 22596
rect 25620 22540 27804 22596
rect 27860 22540 27870 22596
rect 0 22260 800 22288
rect 29200 22260 30000 22288
rect 0 22204 2268 22260
rect 2324 22204 2334 22260
rect 26450 22204 26460 22260
rect 26516 22204 27468 22260
rect 27524 22204 30000 22260
rect 0 22176 800 22204
rect 29200 22176 30000 22204
rect 8006 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8290 21980
rect 14810 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15094 21980
rect 21614 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21898 21980
rect 28418 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28702 21980
rect 2930 21756 2940 21812
rect 2996 21756 5740 21812
rect 5796 21756 5806 21812
rect 25442 21756 25452 21812
rect 25508 21756 27804 21812
rect 27860 21756 27870 21812
rect 20626 21644 20636 21700
rect 20692 21644 22204 21700
rect 22260 21644 22270 21700
rect 0 21588 800 21616
rect 29200 21588 30000 21616
rect 0 21532 2156 21588
rect 2212 21532 2222 21588
rect 28018 21532 28028 21588
rect 28084 21532 30000 21588
rect 0 21504 800 21532
rect 29200 21504 30000 21532
rect 27122 21420 27132 21476
rect 27188 21420 28140 21476
rect 28196 21420 28206 21476
rect 4604 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4888 21196
rect 11408 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11692 21196
rect 18212 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18496 21196
rect 25016 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25300 21196
rect 0 20916 800 20944
rect 29200 20916 30000 20944
rect 0 20860 2380 20916
rect 2436 20860 2446 20916
rect 12114 20860 12124 20916
rect 12180 20860 14476 20916
rect 14532 20860 14542 20916
rect 28130 20860 28140 20916
rect 28196 20860 30000 20916
rect 0 20832 800 20860
rect 29200 20832 30000 20860
rect 25778 20748 25788 20804
rect 25844 20748 26908 20804
rect 26964 20748 26974 20804
rect 2034 20636 2044 20692
rect 2100 20636 6076 20692
rect 6132 20636 6142 20692
rect 8006 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8290 20412
rect 14810 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15094 20412
rect 21614 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21898 20412
rect 28418 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28702 20412
rect 0 20244 800 20272
rect 29200 20244 30000 20272
rect 0 20188 1820 20244
rect 1876 20188 1886 20244
rect 28018 20188 28028 20244
rect 28084 20188 30000 20244
rect 0 20160 800 20188
rect 29200 20160 30000 20188
rect 19282 20076 19292 20132
rect 19348 20076 21196 20132
rect 21252 20076 21262 20132
rect 24882 19964 24892 20020
rect 24948 19964 26908 20020
rect 26964 19964 26974 20020
rect 17602 19852 17612 19908
rect 17668 19852 21196 19908
rect 21252 19852 21262 19908
rect 15922 19740 15932 19796
rect 15988 19740 18396 19796
rect 18452 19740 18462 19796
rect 15362 19628 15372 19684
rect 15428 19628 16268 19684
rect 16324 19628 16334 19684
rect 4604 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4888 19628
rect 11408 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11692 19628
rect 18212 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18496 19628
rect 25016 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25300 19628
rect 29200 19572 30000 19600
rect 28018 19516 28028 19572
rect 28084 19516 30000 19572
rect 29200 19488 30000 19516
rect 7746 19292 7756 19348
rect 7812 19292 8652 19348
rect 8708 19292 8718 19348
rect 10434 19292 10444 19348
rect 10500 19292 11452 19348
rect 11508 19292 11518 19348
rect 13906 19292 13916 19348
rect 13972 19292 15260 19348
rect 15316 19292 15326 19348
rect 10770 19068 10780 19124
rect 10836 19068 12460 19124
rect 12516 19068 12526 19124
rect 24770 19068 24780 19124
rect 24836 19068 27804 19124
rect 27860 19068 27870 19124
rect 1708 18956 14252 19012
rect 14308 18956 14318 19012
rect 18946 18956 18956 19012
rect 19012 18956 22204 19012
rect 22260 18956 22270 19012
rect 0 18900 800 18928
rect 1708 18900 1764 18956
rect 29200 18900 30000 18928
rect 0 18844 1764 18900
rect 28812 18844 30000 18900
rect 0 18816 800 18844
rect 8006 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8290 18844
rect 14810 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15094 18844
rect 21614 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21898 18844
rect 28418 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28702 18844
rect 28812 18676 28868 18844
rect 29200 18816 30000 18844
rect 16930 18620 16940 18676
rect 16996 18620 19404 18676
rect 19460 18620 19470 18676
rect 28242 18620 28252 18676
rect 28308 18620 28868 18676
rect 6290 18508 6300 18564
rect 6356 18508 7644 18564
rect 7700 18508 7710 18564
rect 20066 18508 20076 18564
rect 20132 18508 21644 18564
rect 21700 18508 21710 18564
rect 9426 18396 9436 18452
rect 9492 18396 11228 18452
rect 11284 18396 13244 18452
rect 13300 18396 13310 18452
rect 17154 18396 17164 18452
rect 17220 18396 18732 18452
rect 18788 18396 19404 18452
rect 19460 18396 19470 18452
rect 22418 18396 22428 18452
rect 22484 18396 27244 18452
rect 27300 18396 27310 18452
rect 13122 18284 13132 18340
rect 13188 18284 15484 18340
rect 15540 18284 15550 18340
rect 16370 18284 16380 18340
rect 16436 18284 18172 18340
rect 18228 18284 19068 18340
rect 19124 18284 19628 18340
rect 19684 18284 19694 18340
rect 21858 18284 21868 18340
rect 21924 18284 26236 18340
rect 26292 18284 26302 18340
rect 23090 18172 23100 18228
rect 23156 18172 23772 18228
rect 23828 18172 23838 18228
rect 24546 18172 24556 18228
rect 24612 18172 26124 18228
rect 26180 18172 26190 18228
rect 4604 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4888 18060
rect 11408 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11692 18060
rect 18212 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18496 18060
rect 25016 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25300 18060
rect 24322 17724 24332 17780
rect 24388 17724 26124 17780
rect 26180 17724 26190 17780
rect 7074 17612 7084 17668
rect 7140 17612 9436 17668
rect 9492 17612 9502 17668
rect 14578 17612 14588 17668
rect 14644 17612 15260 17668
rect 15316 17612 17164 17668
rect 17220 17612 17230 17668
rect 19394 17612 19404 17668
rect 19460 17612 21196 17668
rect 21252 17612 23212 17668
rect 23268 17612 23278 17668
rect 23874 17612 23884 17668
rect 23940 17612 26684 17668
rect 26740 17612 26750 17668
rect 29200 17556 30000 17584
rect 4834 17500 4844 17556
rect 4900 17500 5852 17556
rect 5908 17500 5918 17556
rect 27794 17500 27804 17556
rect 27860 17500 30000 17556
rect 29200 17472 30000 17500
rect 24882 17388 24892 17444
rect 24948 17388 27244 17444
rect 27300 17388 27310 17444
rect 8006 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8290 17276
rect 14810 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15094 17276
rect 21614 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21898 17276
rect 28418 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28702 17276
rect 4834 16940 4844 16996
rect 4900 16940 6860 16996
rect 6916 16940 7588 16996
rect 7532 16884 7588 16940
rect 29200 16884 30000 16912
rect 3154 16828 3164 16884
rect 3220 16828 4956 16884
rect 5012 16828 5404 16884
rect 5460 16828 7084 16884
rect 7140 16828 7150 16884
rect 7522 16828 7532 16884
rect 7588 16828 10220 16884
rect 10276 16828 10286 16884
rect 28130 16828 28140 16884
rect 28196 16828 30000 16884
rect 29200 16800 30000 16828
rect 13682 16716 13692 16772
rect 13748 16716 14140 16772
rect 14196 16716 16380 16772
rect 16436 16716 16446 16772
rect 23314 16716 23324 16772
rect 23380 16716 26236 16772
rect 26292 16716 26302 16772
rect 6290 16604 6300 16660
rect 6356 16604 7308 16660
rect 7364 16604 7374 16660
rect 4604 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4888 16492
rect 11408 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11692 16492
rect 18212 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18496 16492
rect 25016 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25300 16492
rect 4946 16156 4956 16212
rect 5012 16156 9996 16212
rect 10052 16156 10062 16212
rect 12898 16044 12908 16100
rect 12964 16044 13692 16100
rect 13748 16044 13758 16100
rect 22754 16044 22764 16100
rect 22820 16044 23212 16100
rect 23268 16044 24668 16100
rect 24724 16044 24734 16100
rect 6626 15932 6636 15988
rect 6692 15932 7308 15988
rect 7364 15932 7374 15988
rect 26338 15932 26348 15988
rect 26404 15932 27692 15988
rect 27748 15932 27758 15988
rect 11890 15820 11900 15876
rect 11956 15820 13580 15876
rect 13636 15820 13646 15876
rect 15922 15820 15932 15876
rect 15988 15820 17500 15876
rect 17556 15820 17566 15876
rect 21186 15820 21196 15876
rect 21252 15820 22316 15876
rect 22372 15820 22382 15876
rect 8006 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8290 15708
rect 14810 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15094 15708
rect 21614 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21898 15708
rect 28418 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28702 15708
rect 5506 15372 5516 15428
rect 5572 15372 7980 15428
rect 8036 15372 8046 15428
rect 23538 15260 23548 15316
rect 23604 15260 24332 15316
rect 24388 15260 25228 15316
rect 25284 15260 25676 15316
rect 25732 15260 25742 15316
rect 19058 15148 19068 15204
rect 19124 15148 21308 15204
rect 21364 15148 21374 15204
rect 21970 15148 21980 15204
rect 22036 15148 26908 15204
rect 26964 15148 26974 15204
rect 4604 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4888 14924
rect 11408 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11692 14924
rect 18212 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18496 14924
rect 25016 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25300 14924
rect 2706 14700 2716 14756
rect 2772 14700 3948 14756
rect 4004 14700 4014 14756
rect 3490 14364 3500 14420
rect 3556 14364 6748 14420
rect 6804 14364 6814 14420
rect 13010 14252 13020 14308
rect 13076 14252 13916 14308
rect 13972 14252 13982 14308
rect 20850 14252 20860 14308
rect 20916 14252 22092 14308
rect 22148 14252 23436 14308
rect 23492 14252 23502 14308
rect 8006 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8290 14140
rect 14810 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15094 14140
rect 21614 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21898 14140
rect 28418 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28702 14140
rect 9202 13804 9212 13860
rect 9268 13804 11788 13860
rect 11844 13804 11854 13860
rect 21298 13804 21308 13860
rect 21364 13804 22764 13860
rect 22820 13804 22830 13860
rect 9986 13580 9996 13636
rect 10052 13580 10780 13636
rect 10836 13580 10846 13636
rect 14242 13580 14252 13636
rect 14308 13580 15036 13636
rect 15092 13580 15102 13636
rect 4722 13468 4732 13524
rect 4788 13468 6524 13524
rect 6580 13468 6590 13524
rect 6178 13356 6188 13412
rect 6244 13356 6972 13412
rect 7028 13356 7038 13412
rect 4604 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4888 13356
rect 11408 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11692 13356
rect 18212 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18496 13356
rect 25016 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25300 13356
rect 2370 13132 2380 13188
rect 2436 13132 3276 13188
rect 3332 13132 3342 13188
rect 2370 12908 2380 12964
rect 2436 12908 5180 12964
rect 5236 12908 5516 12964
rect 5572 12908 6972 12964
rect 7028 12908 7868 12964
rect 7924 12908 8988 12964
rect 9044 12908 9054 12964
rect 12450 12908 12460 12964
rect 12516 12908 20748 12964
rect 20804 12908 20814 12964
rect 3378 12796 3388 12852
rect 3444 12796 4172 12852
rect 4228 12796 4620 12852
rect 4676 12796 4686 12852
rect 1698 12684 1708 12740
rect 1764 12684 2492 12740
rect 2548 12684 2558 12740
rect 22306 12684 22316 12740
rect 22372 12684 24108 12740
rect 24164 12684 24174 12740
rect 25106 12684 25116 12740
rect 25172 12684 26012 12740
rect 26068 12684 26078 12740
rect 8006 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8290 12572
rect 14810 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15094 12572
rect 21614 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21898 12572
rect 28418 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28702 12572
rect 22642 12460 22652 12516
rect 22708 12460 26236 12516
rect 26292 12460 26302 12516
rect 1586 12348 1596 12404
rect 1652 12348 2604 12404
rect 2660 12348 2670 12404
rect 8978 12236 8988 12292
rect 9044 12236 9772 12292
rect 9828 12236 9838 12292
rect 0 12180 800 12208
rect 0 12124 1708 12180
rect 1764 12124 1774 12180
rect 14802 12124 14812 12180
rect 14868 12124 19516 12180
rect 19572 12124 19582 12180
rect 0 12096 800 12124
rect 21410 12012 21420 12068
rect 21476 12012 22204 12068
rect 22260 12012 24444 12068
rect 24500 12012 24510 12068
rect 4610 11900 4620 11956
rect 4676 11900 5012 11956
rect 4956 11844 5012 11900
rect 24892 11900 27244 11956
rect 27300 11900 27310 11956
rect 24892 11844 24948 11900
rect 4956 11788 8428 11844
rect 24882 11788 24892 11844
rect 24948 11788 24958 11844
rect 4604 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4888 11788
rect 8372 11732 8428 11788
rect 11408 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11692 11788
rect 18212 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18496 11788
rect 25016 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25300 11788
rect 5954 11676 5964 11732
rect 6020 11676 8540 11732
rect 8596 11676 9100 11732
rect 9156 11676 10220 11732
rect 10276 11676 10286 11732
rect 13906 11452 13916 11508
rect 13972 11452 16268 11508
rect 16324 11452 16334 11508
rect 17938 11452 17948 11508
rect 18004 11452 19292 11508
rect 19348 11452 19358 11508
rect 16258 11228 16268 11284
rect 16324 11228 17276 11284
rect 17332 11228 17342 11284
rect 18946 11228 18956 11284
rect 19012 11228 20300 11284
rect 20356 11228 20366 11284
rect 25666 11228 25676 11284
rect 25732 11228 27692 11284
rect 27748 11228 27758 11284
rect 3154 11004 3164 11060
rect 3220 11004 4844 11060
rect 4900 11004 4910 11060
rect 8006 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8290 11004
rect 14810 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15094 11004
rect 21614 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21898 11004
rect 28418 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28702 11004
rect 10098 10780 10108 10836
rect 10164 10780 12348 10836
rect 12404 10780 12414 10836
rect 19058 10780 19068 10836
rect 19124 10780 20188 10836
rect 20244 10780 20254 10836
rect 9314 10668 9324 10724
rect 9380 10668 11788 10724
rect 11844 10668 11854 10724
rect 3042 10556 3052 10612
rect 3108 10556 3724 10612
rect 3780 10556 3790 10612
rect 13234 10556 13244 10612
rect 13300 10556 14476 10612
rect 14532 10556 14542 10612
rect 6626 10444 6636 10500
rect 6692 10444 7532 10500
rect 7588 10444 7598 10500
rect 9986 10444 9996 10500
rect 10052 10444 10780 10500
rect 10836 10444 10846 10500
rect 21746 10444 21756 10500
rect 21812 10444 26236 10500
rect 26292 10444 26302 10500
rect 2034 10332 2044 10388
rect 2100 10332 9772 10388
rect 9828 10332 9838 10388
rect 20962 10332 20972 10388
rect 21028 10332 26908 10388
rect 26964 10332 26974 10388
rect 0 10164 800 10192
rect 4604 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4888 10220
rect 11408 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11692 10220
rect 18212 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18496 10220
rect 25016 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25300 10220
rect 29200 10164 30000 10192
rect 0 10108 1820 10164
rect 1876 10108 1886 10164
rect 25554 10108 25564 10164
rect 25620 10108 27244 10164
rect 27300 10108 27310 10164
rect 27692 10108 30000 10164
rect 0 10080 800 10108
rect 27692 10052 27748 10108
rect 29200 10080 30000 10108
rect 23762 9996 23772 10052
rect 23828 9996 26684 10052
rect 26740 9996 26750 10052
rect 27682 9996 27692 10052
rect 27748 9996 27758 10052
rect 7858 9884 7868 9940
rect 7924 9884 8428 9940
rect 8372 9828 8428 9884
rect 14700 9884 16828 9940
rect 16884 9884 17948 9940
rect 18004 9884 18732 9940
rect 18788 9884 19180 9940
rect 19236 9884 19246 9940
rect 20132 9884 21308 9940
rect 21364 9884 21374 9940
rect 14700 9828 14756 9884
rect 20132 9828 20188 9884
rect 8372 9772 9548 9828
rect 9604 9772 12908 9828
rect 12964 9772 12974 9828
rect 14130 9772 14140 9828
rect 14196 9772 14700 9828
rect 14756 9772 14766 9828
rect 15474 9772 15484 9828
rect 15540 9772 17276 9828
rect 17332 9772 19964 9828
rect 20020 9772 20188 9828
rect 21858 9772 21868 9828
rect 21924 9772 22988 9828
rect 23044 9772 23054 9828
rect 5506 9660 5516 9716
rect 5572 9660 7644 9716
rect 7700 9660 7710 9716
rect 12450 9660 12460 9716
rect 12516 9660 13916 9716
rect 13972 9660 13982 9716
rect 18386 9548 18396 9604
rect 18452 9548 19292 9604
rect 19348 9548 19358 9604
rect 8006 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8290 9436
rect 14810 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15094 9436
rect 21614 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21898 9436
rect 28418 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28702 9436
rect 20850 9212 20860 9268
rect 20916 9212 21644 9268
rect 21700 9212 23548 9268
rect 23604 9212 23772 9268
rect 23828 9212 24332 9268
rect 24388 9212 25452 9268
rect 25508 9212 25518 9268
rect 11890 8876 11900 8932
rect 11956 8876 12684 8932
rect 12740 8876 14140 8932
rect 14196 8876 14206 8932
rect 22530 8876 22540 8932
rect 22596 8876 26236 8932
rect 26292 8876 26302 8932
rect 29200 8820 30000 8848
rect 29036 8764 30000 8820
rect 4604 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4888 8652
rect 11408 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11692 8652
rect 18212 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18496 8652
rect 25016 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25300 8652
rect 29036 8484 29092 8764
rect 29200 8736 30000 8764
rect 29036 8428 29316 8484
rect 29260 8372 29316 8428
rect 15922 8316 15932 8372
rect 15988 8316 17612 8372
rect 17668 8316 17678 8372
rect 27682 8316 27692 8372
rect 27748 8316 29316 8372
rect 0 8148 800 8176
rect 29200 8148 30000 8176
rect 0 8092 3388 8148
rect 3444 8092 4060 8148
rect 4116 8092 4126 8148
rect 13346 8092 13356 8148
rect 13412 8092 15484 8148
rect 15540 8092 15550 8148
rect 16930 8092 16940 8148
rect 16996 8092 18620 8148
rect 18676 8092 18686 8148
rect 28130 8092 28140 8148
rect 28196 8092 30000 8148
rect 0 8064 800 8092
rect 29200 8064 30000 8092
rect 8006 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8290 7868
rect 14810 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15094 7868
rect 21614 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21898 7868
rect 28418 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28702 7868
rect 2930 7644 2940 7700
rect 2996 7644 3836 7700
rect 3892 7644 3902 7700
rect 22082 7532 22092 7588
rect 22148 7532 23100 7588
rect 23156 7532 23166 7588
rect 0 7476 800 7504
rect 29200 7476 30000 7504
rect 0 7420 2044 7476
rect 2100 7420 2110 7476
rect 27682 7420 27692 7476
rect 27748 7420 30000 7476
rect 0 7392 800 7420
rect 29200 7392 30000 7420
rect 4604 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4888 7084
rect 11408 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11692 7084
rect 18212 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18496 7084
rect 25016 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25300 7084
rect 23762 6860 23772 6916
rect 23828 6860 27804 6916
rect 27860 6860 27870 6916
rect 0 6804 800 6832
rect 29200 6804 30000 6832
rect 0 6748 1932 6804
rect 1988 6748 1998 6804
rect 2930 6748 2940 6804
rect 2996 6748 4172 6804
rect 4228 6748 4238 6804
rect 25666 6748 25676 6804
rect 25732 6748 27244 6804
rect 27300 6748 27310 6804
rect 27570 6748 27580 6804
rect 27636 6748 30000 6804
rect 0 6720 800 6748
rect 29200 6720 30000 6748
rect 22978 6636 22988 6692
rect 23044 6636 26796 6692
rect 26852 6636 26862 6692
rect 2034 6524 2044 6580
rect 2100 6524 4172 6580
rect 4228 6524 4238 6580
rect 8006 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8290 6300
rect 14810 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15094 6300
rect 21614 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21898 6300
rect 28418 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28702 6300
rect 0 6132 800 6160
rect 29200 6132 30000 6160
rect 0 6076 1708 6132
rect 1764 6076 2492 6132
rect 2548 6076 2558 6132
rect 23874 6076 23884 6132
rect 23940 6076 25452 6132
rect 25508 6076 25518 6132
rect 27692 6076 30000 6132
rect 0 6048 800 6076
rect 23986 5964 23996 6020
rect 24052 5964 25676 6020
rect 25732 5964 25742 6020
rect 27692 5908 27748 6076
rect 29200 6048 30000 6076
rect 9202 5852 9212 5908
rect 9268 5852 9996 5908
rect 10052 5852 10062 5908
rect 23314 5852 23324 5908
rect 23380 5852 24332 5908
rect 24388 5852 24398 5908
rect 27682 5852 27692 5908
rect 27748 5852 27758 5908
rect 2034 5628 2044 5684
rect 2100 5628 3388 5684
rect 3444 5628 3454 5684
rect 0 5460 800 5488
rect 4604 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4888 5516
rect 11408 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11692 5516
rect 18212 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18496 5516
rect 25016 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25300 5516
rect 29200 5460 30000 5488
rect 0 5404 1932 5460
rect 1988 5404 1998 5460
rect 27346 5404 27356 5460
rect 27412 5404 30000 5460
rect 0 5376 800 5404
rect 29200 5376 30000 5404
rect 24098 5180 24108 5236
rect 24164 5180 25900 5236
rect 25956 5180 25966 5236
rect 24658 5068 24668 5124
rect 24724 5068 26908 5124
rect 26964 5068 26974 5124
rect 23986 4956 23996 5012
rect 24052 4956 27244 5012
rect 27300 4956 27310 5012
rect 25442 4844 25452 4900
rect 25508 4844 28868 4900
rect 0 4788 800 4816
rect 28812 4788 28868 4844
rect 29200 4788 30000 4816
rect 0 4732 1708 4788
rect 1764 4732 2492 4788
rect 2548 4732 2558 4788
rect 28812 4732 30000 4788
rect 0 4704 800 4732
rect 8006 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8290 4732
rect 14810 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15094 4732
rect 21614 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21898 4732
rect 28418 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28702 4732
rect 29200 4704 30000 4732
rect 11106 4620 11116 4676
rect 11172 4620 13132 4676
rect 13188 4620 13198 4676
rect 24882 4620 24892 4676
rect 24948 4620 25900 4676
rect 25956 4620 25966 4676
rect 10882 4508 10892 4564
rect 10948 4508 11900 4564
rect 11956 4508 11966 4564
rect 25778 4508 25788 4564
rect 25844 4508 26908 4564
rect 26964 4508 26974 4564
rect 25554 4396 25564 4452
rect 25620 4396 26460 4452
rect 26516 4396 26526 4452
rect 29200 4116 30000 4144
rect 27458 4060 27468 4116
rect 27524 4060 30000 4116
rect 29200 4032 30000 4060
rect 4604 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4888 3948
rect 11408 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11692 3948
rect 18212 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18496 3948
rect 25016 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25300 3948
rect 12114 3612 12124 3668
rect 12180 3612 13580 3668
rect 13636 3612 13646 3668
rect 29200 3444 30000 3472
rect 24322 3388 24332 3444
rect 24388 3388 24892 3444
rect 24948 3388 30000 3444
rect 29200 3360 30000 3388
rect 8006 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8290 3164
rect 14810 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15094 3164
rect 21614 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21898 3164
rect 28418 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28702 3164
rect 29200 2772 30000 2800
rect 23090 2716 23100 2772
rect 23156 2716 30000 2772
rect 29200 2688 30000 2716
rect 29200 2100 30000 2128
rect 24658 2044 24668 2100
rect 24724 2044 30000 2100
rect 29200 2016 30000 2044
rect 29200 1428 30000 1456
rect 23762 1372 23772 1428
rect 23828 1372 30000 1428
rect 29200 1344 30000 1372
<< via3 >>
rect 8016 26628 8072 26684
rect 8120 26628 8176 26684
rect 8224 26628 8280 26684
rect 14820 26628 14876 26684
rect 14924 26628 14980 26684
rect 15028 26628 15084 26684
rect 21624 26628 21680 26684
rect 21728 26628 21784 26684
rect 21832 26628 21888 26684
rect 28428 26628 28484 26684
rect 28532 26628 28588 26684
rect 28636 26628 28692 26684
rect 4614 25844 4670 25900
rect 4718 25844 4774 25900
rect 4822 25844 4878 25900
rect 11418 25844 11474 25900
rect 11522 25844 11578 25900
rect 11626 25844 11682 25900
rect 18222 25844 18278 25900
rect 18326 25844 18382 25900
rect 18430 25844 18486 25900
rect 25026 25844 25082 25900
rect 25130 25844 25186 25900
rect 25234 25844 25290 25900
rect 8016 25060 8072 25116
rect 8120 25060 8176 25116
rect 8224 25060 8280 25116
rect 14820 25060 14876 25116
rect 14924 25060 14980 25116
rect 15028 25060 15084 25116
rect 21624 25060 21680 25116
rect 21728 25060 21784 25116
rect 21832 25060 21888 25116
rect 28428 25060 28484 25116
rect 28532 25060 28588 25116
rect 28636 25060 28692 25116
rect 4614 24276 4670 24332
rect 4718 24276 4774 24332
rect 4822 24276 4878 24332
rect 11418 24276 11474 24332
rect 11522 24276 11578 24332
rect 11626 24276 11682 24332
rect 18222 24276 18278 24332
rect 18326 24276 18382 24332
rect 18430 24276 18486 24332
rect 25026 24276 25082 24332
rect 25130 24276 25186 24332
rect 25234 24276 25290 24332
rect 8016 23492 8072 23548
rect 8120 23492 8176 23548
rect 8224 23492 8280 23548
rect 14820 23492 14876 23548
rect 14924 23492 14980 23548
rect 15028 23492 15084 23548
rect 21624 23492 21680 23548
rect 21728 23492 21784 23548
rect 21832 23492 21888 23548
rect 28428 23492 28484 23548
rect 28532 23492 28588 23548
rect 28636 23492 28692 23548
rect 4614 22708 4670 22764
rect 4718 22708 4774 22764
rect 4822 22708 4878 22764
rect 11418 22708 11474 22764
rect 11522 22708 11578 22764
rect 11626 22708 11682 22764
rect 18222 22708 18278 22764
rect 18326 22708 18382 22764
rect 18430 22708 18486 22764
rect 25026 22708 25082 22764
rect 25130 22708 25186 22764
rect 25234 22708 25290 22764
rect 8016 21924 8072 21980
rect 8120 21924 8176 21980
rect 8224 21924 8280 21980
rect 14820 21924 14876 21980
rect 14924 21924 14980 21980
rect 15028 21924 15084 21980
rect 21624 21924 21680 21980
rect 21728 21924 21784 21980
rect 21832 21924 21888 21980
rect 28428 21924 28484 21980
rect 28532 21924 28588 21980
rect 28636 21924 28692 21980
rect 4614 21140 4670 21196
rect 4718 21140 4774 21196
rect 4822 21140 4878 21196
rect 11418 21140 11474 21196
rect 11522 21140 11578 21196
rect 11626 21140 11682 21196
rect 18222 21140 18278 21196
rect 18326 21140 18382 21196
rect 18430 21140 18486 21196
rect 25026 21140 25082 21196
rect 25130 21140 25186 21196
rect 25234 21140 25290 21196
rect 8016 20356 8072 20412
rect 8120 20356 8176 20412
rect 8224 20356 8280 20412
rect 14820 20356 14876 20412
rect 14924 20356 14980 20412
rect 15028 20356 15084 20412
rect 21624 20356 21680 20412
rect 21728 20356 21784 20412
rect 21832 20356 21888 20412
rect 28428 20356 28484 20412
rect 28532 20356 28588 20412
rect 28636 20356 28692 20412
rect 4614 19572 4670 19628
rect 4718 19572 4774 19628
rect 4822 19572 4878 19628
rect 11418 19572 11474 19628
rect 11522 19572 11578 19628
rect 11626 19572 11682 19628
rect 18222 19572 18278 19628
rect 18326 19572 18382 19628
rect 18430 19572 18486 19628
rect 25026 19572 25082 19628
rect 25130 19572 25186 19628
rect 25234 19572 25290 19628
rect 8016 18788 8072 18844
rect 8120 18788 8176 18844
rect 8224 18788 8280 18844
rect 14820 18788 14876 18844
rect 14924 18788 14980 18844
rect 15028 18788 15084 18844
rect 21624 18788 21680 18844
rect 21728 18788 21784 18844
rect 21832 18788 21888 18844
rect 28428 18788 28484 18844
rect 28532 18788 28588 18844
rect 28636 18788 28692 18844
rect 4614 18004 4670 18060
rect 4718 18004 4774 18060
rect 4822 18004 4878 18060
rect 11418 18004 11474 18060
rect 11522 18004 11578 18060
rect 11626 18004 11682 18060
rect 18222 18004 18278 18060
rect 18326 18004 18382 18060
rect 18430 18004 18486 18060
rect 25026 18004 25082 18060
rect 25130 18004 25186 18060
rect 25234 18004 25290 18060
rect 8016 17220 8072 17276
rect 8120 17220 8176 17276
rect 8224 17220 8280 17276
rect 14820 17220 14876 17276
rect 14924 17220 14980 17276
rect 15028 17220 15084 17276
rect 21624 17220 21680 17276
rect 21728 17220 21784 17276
rect 21832 17220 21888 17276
rect 28428 17220 28484 17276
rect 28532 17220 28588 17276
rect 28636 17220 28692 17276
rect 4614 16436 4670 16492
rect 4718 16436 4774 16492
rect 4822 16436 4878 16492
rect 11418 16436 11474 16492
rect 11522 16436 11578 16492
rect 11626 16436 11682 16492
rect 18222 16436 18278 16492
rect 18326 16436 18382 16492
rect 18430 16436 18486 16492
rect 25026 16436 25082 16492
rect 25130 16436 25186 16492
rect 25234 16436 25290 16492
rect 8016 15652 8072 15708
rect 8120 15652 8176 15708
rect 8224 15652 8280 15708
rect 14820 15652 14876 15708
rect 14924 15652 14980 15708
rect 15028 15652 15084 15708
rect 21624 15652 21680 15708
rect 21728 15652 21784 15708
rect 21832 15652 21888 15708
rect 28428 15652 28484 15708
rect 28532 15652 28588 15708
rect 28636 15652 28692 15708
rect 4614 14868 4670 14924
rect 4718 14868 4774 14924
rect 4822 14868 4878 14924
rect 11418 14868 11474 14924
rect 11522 14868 11578 14924
rect 11626 14868 11682 14924
rect 18222 14868 18278 14924
rect 18326 14868 18382 14924
rect 18430 14868 18486 14924
rect 25026 14868 25082 14924
rect 25130 14868 25186 14924
rect 25234 14868 25290 14924
rect 8016 14084 8072 14140
rect 8120 14084 8176 14140
rect 8224 14084 8280 14140
rect 14820 14084 14876 14140
rect 14924 14084 14980 14140
rect 15028 14084 15084 14140
rect 21624 14084 21680 14140
rect 21728 14084 21784 14140
rect 21832 14084 21888 14140
rect 28428 14084 28484 14140
rect 28532 14084 28588 14140
rect 28636 14084 28692 14140
rect 4614 13300 4670 13356
rect 4718 13300 4774 13356
rect 4822 13300 4878 13356
rect 11418 13300 11474 13356
rect 11522 13300 11578 13356
rect 11626 13300 11682 13356
rect 18222 13300 18278 13356
rect 18326 13300 18382 13356
rect 18430 13300 18486 13356
rect 25026 13300 25082 13356
rect 25130 13300 25186 13356
rect 25234 13300 25290 13356
rect 8016 12516 8072 12572
rect 8120 12516 8176 12572
rect 8224 12516 8280 12572
rect 14820 12516 14876 12572
rect 14924 12516 14980 12572
rect 15028 12516 15084 12572
rect 21624 12516 21680 12572
rect 21728 12516 21784 12572
rect 21832 12516 21888 12572
rect 28428 12516 28484 12572
rect 28532 12516 28588 12572
rect 28636 12516 28692 12572
rect 4614 11732 4670 11788
rect 4718 11732 4774 11788
rect 4822 11732 4878 11788
rect 11418 11732 11474 11788
rect 11522 11732 11578 11788
rect 11626 11732 11682 11788
rect 18222 11732 18278 11788
rect 18326 11732 18382 11788
rect 18430 11732 18486 11788
rect 25026 11732 25082 11788
rect 25130 11732 25186 11788
rect 25234 11732 25290 11788
rect 8016 10948 8072 11004
rect 8120 10948 8176 11004
rect 8224 10948 8280 11004
rect 14820 10948 14876 11004
rect 14924 10948 14980 11004
rect 15028 10948 15084 11004
rect 21624 10948 21680 11004
rect 21728 10948 21784 11004
rect 21832 10948 21888 11004
rect 28428 10948 28484 11004
rect 28532 10948 28588 11004
rect 28636 10948 28692 11004
rect 4614 10164 4670 10220
rect 4718 10164 4774 10220
rect 4822 10164 4878 10220
rect 11418 10164 11474 10220
rect 11522 10164 11578 10220
rect 11626 10164 11682 10220
rect 18222 10164 18278 10220
rect 18326 10164 18382 10220
rect 18430 10164 18486 10220
rect 25026 10164 25082 10220
rect 25130 10164 25186 10220
rect 25234 10164 25290 10220
rect 8016 9380 8072 9436
rect 8120 9380 8176 9436
rect 8224 9380 8280 9436
rect 14820 9380 14876 9436
rect 14924 9380 14980 9436
rect 15028 9380 15084 9436
rect 21624 9380 21680 9436
rect 21728 9380 21784 9436
rect 21832 9380 21888 9436
rect 28428 9380 28484 9436
rect 28532 9380 28588 9436
rect 28636 9380 28692 9436
rect 4614 8596 4670 8652
rect 4718 8596 4774 8652
rect 4822 8596 4878 8652
rect 11418 8596 11474 8652
rect 11522 8596 11578 8652
rect 11626 8596 11682 8652
rect 18222 8596 18278 8652
rect 18326 8596 18382 8652
rect 18430 8596 18486 8652
rect 25026 8596 25082 8652
rect 25130 8596 25186 8652
rect 25234 8596 25290 8652
rect 8016 7812 8072 7868
rect 8120 7812 8176 7868
rect 8224 7812 8280 7868
rect 14820 7812 14876 7868
rect 14924 7812 14980 7868
rect 15028 7812 15084 7868
rect 21624 7812 21680 7868
rect 21728 7812 21784 7868
rect 21832 7812 21888 7868
rect 28428 7812 28484 7868
rect 28532 7812 28588 7868
rect 28636 7812 28692 7868
rect 4614 7028 4670 7084
rect 4718 7028 4774 7084
rect 4822 7028 4878 7084
rect 11418 7028 11474 7084
rect 11522 7028 11578 7084
rect 11626 7028 11682 7084
rect 18222 7028 18278 7084
rect 18326 7028 18382 7084
rect 18430 7028 18486 7084
rect 25026 7028 25082 7084
rect 25130 7028 25186 7084
rect 25234 7028 25290 7084
rect 8016 6244 8072 6300
rect 8120 6244 8176 6300
rect 8224 6244 8280 6300
rect 14820 6244 14876 6300
rect 14924 6244 14980 6300
rect 15028 6244 15084 6300
rect 21624 6244 21680 6300
rect 21728 6244 21784 6300
rect 21832 6244 21888 6300
rect 28428 6244 28484 6300
rect 28532 6244 28588 6300
rect 28636 6244 28692 6300
rect 4614 5460 4670 5516
rect 4718 5460 4774 5516
rect 4822 5460 4878 5516
rect 11418 5460 11474 5516
rect 11522 5460 11578 5516
rect 11626 5460 11682 5516
rect 18222 5460 18278 5516
rect 18326 5460 18382 5516
rect 18430 5460 18486 5516
rect 25026 5460 25082 5516
rect 25130 5460 25186 5516
rect 25234 5460 25290 5516
rect 8016 4676 8072 4732
rect 8120 4676 8176 4732
rect 8224 4676 8280 4732
rect 14820 4676 14876 4732
rect 14924 4676 14980 4732
rect 15028 4676 15084 4732
rect 21624 4676 21680 4732
rect 21728 4676 21784 4732
rect 21832 4676 21888 4732
rect 28428 4676 28484 4732
rect 28532 4676 28588 4732
rect 28636 4676 28692 4732
rect 4614 3892 4670 3948
rect 4718 3892 4774 3948
rect 4822 3892 4878 3948
rect 11418 3892 11474 3948
rect 11522 3892 11578 3948
rect 11626 3892 11682 3948
rect 18222 3892 18278 3948
rect 18326 3892 18382 3948
rect 18430 3892 18486 3948
rect 25026 3892 25082 3948
rect 25130 3892 25186 3948
rect 25234 3892 25290 3948
rect 8016 3108 8072 3164
rect 8120 3108 8176 3164
rect 8224 3108 8280 3164
rect 14820 3108 14876 3164
rect 14924 3108 14980 3164
rect 15028 3108 15084 3164
rect 21624 3108 21680 3164
rect 21728 3108 21784 3164
rect 21832 3108 21888 3164
rect 28428 3108 28484 3164
rect 28532 3108 28588 3164
rect 28636 3108 28692 3164
<< metal4 >>
rect 4586 25900 4906 26716
rect 4586 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4906 25900
rect 4586 24332 4906 25844
rect 4586 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4906 24332
rect 4586 22764 4906 24276
rect 4586 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4906 22764
rect 4586 21196 4906 22708
rect 4586 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4906 21196
rect 4586 19628 4906 21140
rect 4586 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4906 19628
rect 4586 18060 4906 19572
rect 4586 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4906 18060
rect 4586 16492 4906 18004
rect 4586 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4906 16492
rect 4586 14924 4906 16436
rect 4586 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4906 14924
rect 4586 13356 4906 14868
rect 4586 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4906 13356
rect 4586 11788 4906 13300
rect 4586 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4906 11788
rect 4586 10220 4906 11732
rect 4586 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4906 10220
rect 4586 8652 4906 10164
rect 4586 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4906 8652
rect 4586 7084 4906 8596
rect 4586 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4906 7084
rect 4586 5516 4906 7028
rect 4586 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4906 5516
rect 4586 3948 4906 5460
rect 4586 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4906 3948
rect 4586 3076 4906 3892
rect 7988 26684 8308 26716
rect 7988 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8308 26684
rect 7988 25116 8308 26628
rect 7988 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8308 25116
rect 7988 23548 8308 25060
rect 7988 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8308 23548
rect 7988 21980 8308 23492
rect 7988 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8308 21980
rect 7988 20412 8308 21924
rect 7988 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8308 20412
rect 7988 18844 8308 20356
rect 7988 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8308 18844
rect 7988 17276 8308 18788
rect 7988 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8308 17276
rect 7988 15708 8308 17220
rect 7988 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8308 15708
rect 7988 14140 8308 15652
rect 7988 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8308 14140
rect 7988 12572 8308 14084
rect 7988 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8308 12572
rect 7988 11004 8308 12516
rect 7988 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8308 11004
rect 7988 9436 8308 10948
rect 7988 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8308 9436
rect 7988 7868 8308 9380
rect 7988 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8308 7868
rect 7988 6300 8308 7812
rect 7988 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8308 6300
rect 7988 4732 8308 6244
rect 7988 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8308 4732
rect 7988 3164 8308 4676
rect 7988 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8308 3164
rect 7988 3076 8308 3108
rect 11390 25900 11710 26716
rect 11390 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11710 25900
rect 11390 24332 11710 25844
rect 11390 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11710 24332
rect 11390 22764 11710 24276
rect 11390 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11710 22764
rect 11390 21196 11710 22708
rect 11390 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11710 21196
rect 11390 19628 11710 21140
rect 11390 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11710 19628
rect 11390 18060 11710 19572
rect 11390 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11710 18060
rect 11390 16492 11710 18004
rect 11390 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11710 16492
rect 11390 14924 11710 16436
rect 11390 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11710 14924
rect 11390 13356 11710 14868
rect 11390 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11710 13356
rect 11390 11788 11710 13300
rect 11390 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11710 11788
rect 11390 10220 11710 11732
rect 11390 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11710 10220
rect 11390 8652 11710 10164
rect 11390 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11710 8652
rect 11390 7084 11710 8596
rect 11390 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11710 7084
rect 11390 5516 11710 7028
rect 11390 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11710 5516
rect 11390 3948 11710 5460
rect 11390 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11710 3948
rect 11390 3076 11710 3892
rect 14792 26684 15112 26716
rect 14792 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15112 26684
rect 14792 25116 15112 26628
rect 14792 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15112 25116
rect 14792 23548 15112 25060
rect 14792 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15112 23548
rect 14792 21980 15112 23492
rect 14792 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15112 21980
rect 14792 20412 15112 21924
rect 14792 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15112 20412
rect 14792 18844 15112 20356
rect 14792 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15112 18844
rect 14792 17276 15112 18788
rect 14792 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15112 17276
rect 14792 15708 15112 17220
rect 14792 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15112 15708
rect 14792 14140 15112 15652
rect 14792 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15112 14140
rect 14792 12572 15112 14084
rect 14792 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15112 12572
rect 14792 11004 15112 12516
rect 14792 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15112 11004
rect 14792 9436 15112 10948
rect 14792 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15112 9436
rect 14792 7868 15112 9380
rect 14792 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15112 7868
rect 14792 6300 15112 7812
rect 14792 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15112 6300
rect 14792 4732 15112 6244
rect 14792 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15112 4732
rect 14792 3164 15112 4676
rect 14792 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15112 3164
rect 14792 3076 15112 3108
rect 18194 25900 18514 26716
rect 18194 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18514 25900
rect 18194 24332 18514 25844
rect 18194 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18514 24332
rect 18194 22764 18514 24276
rect 18194 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18514 22764
rect 18194 21196 18514 22708
rect 18194 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18514 21196
rect 18194 19628 18514 21140
rect 18194 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18514 19628
rect 18194 18060 18514 19572
rect 18194 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18514 18060
rect 18194 16492 18514 18004
rect 18194 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18514 16492
rect 18194 14924 18514 16436
rect 18194 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18514 14924
rect 18194 13356 18514 14868
rect 18194 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18514 13356
rect 18194 11788 18514 13300
rect 18194 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18514 11788
rect 18194 10220 18514 11732
rect 18194 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18514 10220
rect 18194 8652 18514 10164
rect 18194 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18514 8652
rect 18194 7084 18514 8596
rect 18194 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18514 7084
rect 18194 5516 18514 7028
rect 18194 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18514 5516
rect 18194 3948 18514 5460
rect 18194 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18514 3948
rect 18194 3076 18514 3892
rect 21596 26684 21916 26716
rect 21596 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21916 26684
rect 21596 25116 21916 26628
rect 21596 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21916 25116
rect 21596 23548 21916 25060
rect 21596 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21916 23548
rect 21596 21980 21916 23492
rect 21596 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21916 21980
rect 21596 20412 21916 21924
rect 21596 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21916 20412
rect 21596 18844 21916 20356
rect 21596 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21916 18844
rect 21596 17276 21916 18788
rect 21596 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21916 17276
rect 21596 15708 21916 17220
rect 21596 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21916 15708
rect 21596 14140 21916 15652
rect 21596 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21916 14140
rect 21596 12572 21916 14084
rect 21596 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21916 12572
rect 21596 11004 21916 12516
rect 21596 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21916 11004
rect 21596 9436 21916 10948
rect 21596 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21916 9436
rect 21596 7868 21916 9380
rect 21596 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21916 7868
rect 21596 6300 21916 7812
rect 21596 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21916 6300
rect 21596 4732 21916 6244
rect 21596 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21916 4732
rect 21596 3164 21916 4676
rect 21596 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21916 3164
rect 21596 3076 21916 3108
rect 24998 25900 25318 26716
rect 24998 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25318 25900
rect 24998 24332 25318 25844
rect 24998 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25318 24332
rect 24998 22764 25318 24276
rect 24998 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25318 22764
rect 24998 21196 25318 22708
rect 24998 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25318 21196
rect 24998 19628 25318 21140
rect 24998 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25318 19628
rect 24998 18060 25318 19572
rect 24998 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25318 18060
rect 24998 16492 25318 18004
rect 24998 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25318 16492
rect 24998 14924 25318 16436
rect 24998 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25318 14924
rect 24998 13356 25318 14868
rect 24998 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25318 13356
rect 24998 11788 25318 13300
rect 24998 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25318 11788
rect 24998 10220 25318 11732
rect 24998 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25318 10220
rect 24998 8652 25318 10164
rect 24998 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25318 8652
rect 24998 7084 25318 8596
rect 24998 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25318 7084
rect 24998 5516 25318 7028
rect 24998 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25318 5516
rect 24998 3948 25318 5460
rect 24998 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25318 3948
rect 24998 3076 25318 3892
rect 28400 26684 28720 26716
rect 28400 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28720 26684
rect 28400 25116 28720 26628
rect 28400 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28720 25116
rect 28400 23548 28720 25060
rect 28400 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28720 23548
rect 28400 21980 28720 23492
rect 28400 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28720 21980
rect 28400 20412 28720 21924
rect 28400 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28720 20412
rect 28400 18844 28720 20356
rect 28400 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28720 18844
rect 28400 17276 28720 18788
rect 28400 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28720 17276
rect 28400 15708 28720 17220
rect 28400 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28720 15708
rect 28400 14140 28720 15652
rect 28400 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28720 14140
rect 28400 12572 28720 14084
rect 28400 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28720 12572
rect 28400 11004 28720 12516
rect 28400 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28720 11004
rect 28400 9436 28720 10948
rect 28400 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28720 9436
rect 28400 7868 28720 9380
rect 28400 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28720 7868
rect 28400 6300 28720 7812
rect 28400 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28720 6300
rect 28400 4732 28720 6244
rect 28400 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28720 4732
rect 28400 3164 28720 4676
rect 28400 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28720 3164
rect 28400 3076 28720 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _040_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _041_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12992 0 1 10976
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _042_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _043_
timestamp 1698431365
transform 1 0 7056 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _044_
timestamp 1698431365
transform 1 0 4144 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _045_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _046_
timestamp 1698431365
transform 1 0 3024 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _047_
timestamp 1698431365
transform -1 0 3472 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _048_
timestamp 1698431365
transform -1 0 10528 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _049_
timestamp 1698431365
transform -1 0 7056 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _050_
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _051_
timestamp 1698431365
transform 1 0 3696 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _052_
timestamp 1698431365
transform -1 0 18928 0 1 12544
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _053_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _054_
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _055_
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _056_
timestamp 1698431365
transform -1 0 19600 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _057_
timestamp 1698431365
transform -1 0 18368 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _058_
timestamp 1698431365
transform -1 0 16352 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _059_
timestamp 1698431365
transform -1 0 14448 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _060_
timestamp 1698431365
transform -1 0 12880 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _061_
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _062_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _063_
timestamp 1698431365
transform 1 0 17808 0 -1 9408
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _064_
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _065_
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _066_
timestamp 1698431365
transform -1 0 26208 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _067_
timestamp 1698431365
transform -1 0 24304 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _068_
timestamp 1698431365
transform -1 0 26208 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _069_
timestamp 1698431365
transform 1 0 23744 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _070_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _071_
timestamp 1698431365
transform 1 0 25648 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _072_
timestamp 1698431365
transform 1 0 25760 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _073_
timestamp 1698431365
transform -1 0 22624 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _074_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _075_
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _076_
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _077_
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _078_
timestamp 1698431365
transform -1 0 14448 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _079_
timestamp 1698431365
transform -1 0 12992 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _080_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _081_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _082_
timestamp 1698431365
transform -1 0 7280 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _083_
timestamp 1698431365
transform 1 0 2352 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _084_
timestamp 1698431365
transform -1 0 5376 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _085_
timestamp 1698431365
transform 1 0 1792 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _086_
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _087_
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _088_
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _089_
timestamp 1698431365
transform -1 0 5712 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _090_
timestamp 1698431365
transform -1 0 14896 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _091_
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _092_
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _093_
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _094_
timestamp 1698431365
transform 1 0 15232 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _095_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _096_
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _097_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _098_
timestamp 1698431365
transform 1 0 17584 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _099_
timestamp 1698431365
transform -1 0 19712 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _100_
timestamp 1698431365
transform -1 0 24976 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _101_
timestamp 1698431365
transform 1 0 23184 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _102_
timestamp 1698431365
transform 1 0 22624 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _103_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _104_
timestamp 1698431365
transform -1 0 26880 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _105_
timestamp 1698431365
transform 1 0 21056 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _106_
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _107_
timestamp 1698431365
transform 1 0 22848 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _108_
timestamp 1698431365
transform 1 0 21952 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _109_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _110_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _111_
timestamp 1698431365
transform 1 0 15232 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _112_
timestamp 1698431365
transform 1 0 13216 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _113_
timestamp 1698431365
transform 1 0 12544 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _114_
timestamp 1698431365
transform 1 0 9296 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _115_
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_
timestamp 1698431365
transform 1 0 4144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1698431365
transform 1 0 25088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _127_
timestamp 1698431365
transform 1 0 10528 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1698431365
transform -1 0 4368 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _129_
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1698431365
transform 1 0 9744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698431365
transform 1 0 20720 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1698431365
transform -1 0 27664 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1698431365
transform -1 0 5264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698431365
transform 1 0 17696 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _136_
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _137_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_
timestamp 1698431365
transform -1 0 5488 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1698431365
transform 1 0 10640 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _141_
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _142_
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _143_
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _144_
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _145_
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1698431365
transform -1 0 6272 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _147_
timestamp 1698431365
transform -1 0 3696 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _148_
timestamp 1698431365
transform 1 0 25984 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1698431365
transform 1 0 24640 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _150_
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _152_
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _153_
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_
timestamp 1698431365
transform 1 0 25760 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1698431365
transform -1 0 5040 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _156_
timestamp 1698431365
transform -1 0 11760 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _157_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_
timestamp 1698431365
transform -1 0 4144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _159_
timestamp 1698431365
transform 1 0 26096 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _160_
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _161_
timestamp 1698431365
transform -1 0 11088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1698431365
transform -1 0 23184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1698431365
transform 1 0 23968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1698431365
transform 1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1698431365
transform 1 0 25424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__CLK
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__CLK
timestamp 1698431365
transform -1 0 23072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__CLK
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__CLK
timestamp 1698431365
transform -1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__CLK
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__CLK
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__CLK
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform -1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 24192 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 28336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 28112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 1792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 7616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 4032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 23520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 28336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 28336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 27216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 24416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 18928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 3136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 22848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 11536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 8288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 1792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 20384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 17584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 28336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 1792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cby_1__1__84 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cby_1__1__85
timestamp 1698431365
transform -1 0 14672 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cby_1__1__86
timestamp 1698431365
transform 1 0 27216 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cby_1__1__87
timestamp 1698431365
transform -1 0 22288 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cby_1__1__88
timestamp 1698431365
transform -1 0 14000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cby_1__1__89
timestamp 1698431365
transform 1 0 26544 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1698431365
transform 1 0 19264 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_52 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_79 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_83
timestamp 1698431365
transform 1 0 10640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_95
timestamp 1698431365
transform 1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_114
timestamp 1698431365
transform 1 0 14112 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_130
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_134
timestamp 1698431365
transform 1 0 16352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_154
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_162
timestamp 1698431365
transform 1 0 19488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_212
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_234
timestamp 1698431365
transform 1 0 27552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_76
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_78
timestamp 1698431365
transform 1 0 10080 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_89
timestamp 1698431365
transform 1 0 11312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_99
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_131
timestamp 1698431365
transform 1 0 16016 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_172
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_188
timestamp 1698431365
transform 1 0 22400 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_237
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_69
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_73
timestamp 1698431365
transform 1 0 9520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_81
timestamp 1698431365
transform 1 0 10416 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_97
timestamp 1698431365
transform 1 0 12208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_193
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_201
timestamp 1698431365
transform 1 0 23856 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_203
timestamp 1698431365
transform 1 0 24080 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_224
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_237
timestamp 1698431365
transform 1 0 27888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_16
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_48
timestamp 1698431365
transform 1 0 6720 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_64
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_82
timestamp 1698431365
transform 1 0 10528 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_89
timestamp 1698431365
transform 1 0 11312 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_121
timestamp 1698431365
transform 1 0 14896 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_174
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_190
timestamp 1698431365
transform 1 0 22624 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_198
timestamp 1698431365
transform 1 0 23520 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_237
timestamp 1698431365
transform 1 0 27888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 2240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_12
timestamp 1698431365
transform 1 0 2688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_14
timestamp 1698431365
transform 1 0 2912 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_33
timestamp 1698431365
transform 1 0 5040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_228
timestamp 1698431365
transform 1 0 26880 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_16
timestamp 1698431365
transform 1 0 3136 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_48
timestamp 1698431365
transform 1 0 6720 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_158
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_166
timestamp 1698431365
transform 1 0 19936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_170
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_188
timestamp 1698431365
transform 1 0 22400 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_196
timestamp 1698431365
transform 1 0 23296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_232
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_234
timestamp 1698431365
transform 1 0 27552 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_237
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_22
timestamp 1698431365
transform 1 0 3808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_115
timestamp 1698431365
transform 1 0 14224 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_132
timestamp 1698431365
transform 1 0 16128 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_140
timestamp 1698431365
transform 1 0 17024 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_160
timestamp 1698431365
transform 1 0 19264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_191
timestamp 1698431365
transform 1 0 22736 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_226
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_237
timestamp 1698431365
transform 1 0 27888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_38
timestamp 1698431365
transform 1 0 5600 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_104
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_185
timestamp 1698431365
transform 1 0 22064 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_193
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_197
timestamp 1698431365
transform 1 0 23408 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_214
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_217
timestamp 1698431365
transform 1 0 25648 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_237
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_6
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_22
timestamp 1698431365
transform 1 0 3808 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_30
timestamp 1698431365
transform 1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_62
timestamp 1698431365
transform 1 0 8288 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_70
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_117
timestamp 1698431365
transform 1 0 14448 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_164
timestamp 1698431365
transform 1 0 19712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_168
timestamp 1698431365
transform 1 0 20160 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_59
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_82
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_99
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_237
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_6
timestamp 1698431365
transform 1 0 2016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_25
timestamp 1698431365
transform 1 0 4144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_47
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_63
timestamp 1698431365
transform 1 0 8400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_65
timestamp 1698431365
transform 1 0 8624 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_131
timestamp 1698431365
transform 1 0 16016 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_148
timestamp 1698431365
transform 1 0 17920 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_156
timestamp 1698431365
transform 1 0 18816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_158
timestamp 1698431365
transform 1 0 19040 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_211
timestamp 1698431365
transform 1 0 24976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_215
timestamp 1698431365
transform 1 0 25424 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_223
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_8
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_53
timestamp 1698431365
transform 1 0 7280 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_57
timestamp 1698431365
transform 1 0 7728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_237
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_157
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_183
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_228
timestamp 1698431365
transform 1 0 26880 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_236
timestamp 1698431365
transform 1 0 27776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_240
timestamp 1698431365
transform 1 0 28224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_82
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_99
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_107
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_126
timestamp 1698431365
transform 1 0 15456 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_134
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_179
timestamp 1698431365
transform 1 0 21392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_197
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698431365
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_232
timestamp 1698431365
transform 1 0 27328 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_236
timestamp 1698431365
transform 1 0 27776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_238
timestamp 1698431365
transform 1 0 28000 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_20
timestamp 1698431365
transform 1 0 3584 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_62
timestamp 1698431365
transform 1 0 8288 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_70
timestamp 1698431365
transform 1 0 9184 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_113
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_166
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_170
timestamp 1698431365
transform 1 0 20384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_179
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_4
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_39
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_47
timestamp 1698431365
transform 1 0 6608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_82
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_121
timestamp 1698431365
transform 1 0 14896 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_176
timestamp 1698431365
transform 1 0 21056 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_193
timestamp 1698431365
transform 1 0 22960 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_197
timestamp 1698431365
transform 1 0 23408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_222
timestamp 1698431365
transform 1 0 26208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_226
timestamp 1698431365
transform 1 0 26656 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_237
timestamp 1698431365
transform 1 0 27888 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_58
timestamp 1698431365
transform 1 0 7840 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_74
timestamp 1698431365
transform 1 0 9632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_92
timestamp 1698431365
transform 1 0 11648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_94
timestamp 1698431365
transform 1 0 11872 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_117
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_125
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_129
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_211
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_215
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_223
timestamp 1698431365
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_50
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_61
timestamp 1698431365
transform 1 0 8176 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_237
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_22
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_24
timestamp 1698431365
transform 1 0 4032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_117
timestamp 1698431365
transform 1 0 14448 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_121
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_211
timestamp 1698431365
transform 1 0 24976 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_219
timestamp 1698431365
transform 1 0 25872 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_26
timestamp 1698431365
transform 1 0 4256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_64
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_152
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_189
timestamp 1698431365
transform 1 0 22512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_237
timestamp 1698431365
transform 1 0 27888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_63
timestamp 1698431365
transform 1 0 8400 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_80
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_88
timestamp 1698431365
transform 1 0 11200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_193
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_134
timestamp 1698431365
transform 1 0 16352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_175
timestamp 1698431365
transform 1 0 20944 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_192
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_226
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_115
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_132
timestamp 1698431365
transform 1 0 16128 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_148
timestamp 1698431365
transform 1 0 17920 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_152
timestamp 1698431365
transform 1 0 18368 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_163
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_209
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_16
timestamp 1698431365
transform 1 0 3136 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_192
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_228
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_16
timestamp 1698431365
transform 1 0 3136 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_209
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_217
timestamp 1698431365
transform 1 0 25648 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_221
timestamp 1698431365
transform 1 0 26096 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_93
timestamp 1698431365
transform 1 0 11760 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_125
timestamp 1698431365
transform 1 0 15344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_166
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_170
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_228
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_14
timestamp 1698431365
transform 1 0 2912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_44
timestamp 1698431365
transform 1 0 6272 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_60
timestamp 1698431365
transform 1 0 8064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_68
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_139
timestamp 1698431365
transform 1 0 16912 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_152
timestamp 1698431365
transform 1 0 18368 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_199
timestamp 1698431365
transform 1 0 23632 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_207
timestamp 1698431365
transform 1 0 24528 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_226
timestamp 1698431365
transform 1 0 26656 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_237
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_16
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_37
timestamp 1698431365
transform 1 0 5488 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_87
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_119
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_158
timestamp 1698431365
transform 1 0 19040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_166
timestamp 1698431365
transform 1 0 19936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_170
timestamp 1698431365
transform 1 0 20384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_172
timestamp 1698431365
transform 1 0 20608 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_179
timestamp 1698431365
transform 1 0 21392 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_195
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_223
timestamp 1698431365
transform 1 0 26320 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_237
timestamp 1698431365
transform 1 0 27888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_47
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_52
timestamp 1698431365
transform 1 0 7168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_58
timestamp 1698431365
transform 1 0 7840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_64
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_80
timestamp 1698431365
transform 1 0 10304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_113
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_119
timestamp 1698431365
transform 1 0 14672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_163
timestamp 1698431365
transform 1 0 19600 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_191
timestamp 1698431365
transform 1 0 22736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_203
timestamp 1698431365
transform 1 0 24080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_217
timestamp 1698431365
transform 1 0 25648 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_237
timestamp 1698431365
transform 1 0 27888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_16
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_30
timestamp 1698431365
transform 1 0 4704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_70
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_114
timestamp 1698431365
transform 1 0 14112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_118
timestamp 1698431365
transform 1 0 14560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_120
timestamp 1698431365
transform 1 0 14784 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_131
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_135
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_167
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_184
timestamp 1698431365
transform 1 0 21952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_186
timestamp 1698431365
transform 1 0 22176 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_197
timestamp 1698431365
transform 1 0 23408 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_201
timestamp 1698431365
transform 1 0 23856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_203
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_240
timestamp 1698431365
transform 1 0 28224 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20048 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 19264 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 12432 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 11648 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform -1 0 16128 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 27888 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 8624 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 10304 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 22848 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 22960 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 16128 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 16912 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 7840 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform 1 0 6496 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform -1 0 23408 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 22848 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform 1 0 6160 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 12432 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 27888 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform -1 0 17920 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 27776 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 2352 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 27888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform -1 0 28336 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 27888 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 28336 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 8288 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform -1 0 22400 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 21280 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 28336 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 27664 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 28336 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 16240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 27664 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 3136 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 21952 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 6944 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 3136 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 28336 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 28336 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 28336 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 21840 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 9520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 24416 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 5600 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 8288 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 18928 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 27664 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 22848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 12432 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 17584 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 28336 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input42 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 26768 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform 1 0 24528 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform 1 0 10192 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform 1 0 26768 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output48 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3136 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output49
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output50
timestamp 1698431365
transform 1 0 11536 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output51
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform -1 0 4704 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform 1 0 26768 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output55
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output56
timestamp 1698431365
transform 1 0 14896 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output57
timestamp 1698431365
transform -1 0 3136 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform 1 0 26432 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output60
timestamp 1698431365
transform -1 0 3136 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output62
timestamp 1698431365
transform -1 0 3136 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output63
timestamp 1698431365
transform 1 0 26768 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output64
timestamp 1698431365
transform 1 0 10416 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output66
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output67 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output69
timestamp 1698431365
transform -1 0 3136 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output70
timestamp 1698431365
transform -1 0 3136 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output71
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output72
timestamp 1698431365
transform 1 0 10864 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output73
timestamp 1698431365
transform 1 0 17360 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output74
timestamp 1698431365
transform 1 0 25200 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output75
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output76
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output77
timestamp 1698431365
transform -1 0 3136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output78
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output79
timestamp 1698431365
transform -1 0 11088 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output80
timestamp 1698431365
transform -1 0 3136 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output81
timestamp 1698431365
transform -1 0 26432 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output82
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output83
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_30 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 28560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_31
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_32
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_33
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_34
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_35
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_36
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_37
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_38
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_39
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_40
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_41
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 28560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_42
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_43
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_44
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_45
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_46
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_47
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_48
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_49
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_50
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 28560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 28560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_61
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_62
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_63
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_64
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_65
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_66
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_67
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_68
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_69
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_70
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_71
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_72
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_73
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_74
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_75
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_76
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_77
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_78
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_81
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_86
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_87
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_88
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_89
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_90
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_91
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_92
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_93
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_94
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_95
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_96
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_97
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_98
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_99
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_100
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_101
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_102
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_103
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_104
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_105
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_106
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_107
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_108
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_109
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_110
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_111
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_112
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_113
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_114
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_115
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_116
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_117
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_118
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_119
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_120
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_121
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_122
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_123
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_124
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_125
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_126
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_127
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_128
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_129
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_130
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_131
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_132
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_133
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_134
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_135
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_136
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_137
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_138
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_139
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_140
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_141
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_142
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_143
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_144
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_145
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_146
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_147
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_148
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_149
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_150
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_151
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_152
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_153
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_154
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_155
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_156
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_157
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 29200 10080 30000 10192 0 FreeSans 448 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 5376 29200 5488 30000 0 FreeSans 448 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 19488 29200 19600 30000 0 FreeSans 448 90 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal2 s 6720 29200 6832 30000 0 FreeSans 448 90 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal3 s 29200 18816 30000 18928 0 FreeSans 448 0 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal3 s 29200 22176 30000 22288 0 FreeSans 448 0 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal3 s 29200 28896 30000 29008 0 FreeSans 448 0 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal2 s 16128 29200 16240 30000 0 FreeSans 448 90 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal3 s 29200 24192 30000 24304 0 FreeSans 448 0 0 0 chany_bottom_in[19]
port 12 nsew signal input
flabel metal2 s 15456 29200 15568 30000 0 FreeSans 448 90 0 0 chany_bottom_in[1]
port 13 nsew signal input
flabel metal3 s 29200 27552 30000 27664 0 FreeSans 448 0 0 0 chany_bottom_in[2]
port 14 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 chany_bottom_in[3]
port 15 nsew signal input
flabel metal2 s 20160 29200 20272 30000 0 FreeSans 448 90 0 0 chany_bottom_in[4]
port 16 nsew signal input
flabel metal2 s 7392 29200 7504 30000 0 FreeSans 448 90 0 0 chany_bottom_in[5]
port 17 nsew signal input
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 chany_bottom_in[6]
port 18 nsew signal input
flabel metal3 s 29200 1344 30000 1456 0 FreeSans 448 0 0 0 chany_bottom_in[7]
port 19 nsew signal input
flabel metal3 s 29200 8064 30000 8176 0 FreeSans 448 0 0 0 chany_bottom_in[8]
port 20 nsew signal input
flabel metal3 s 29200 21504 30000 21616 0 FreeSans 448 0 0 0 chany_bottom_in[9]
port 21 nsew signal input
flabel metal3 s 29200 28224 30000 28336 0 FreeSans 448 0 0 0 chany_bottom_out[0]
port 22 nsew signal tristate
flabel metal2 s 24192 29200 24304 30000 0 FreeSans 448 90 0 0 chany_bottom_out[10]
port 23 nsew signal tristate
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chany_bottom_out[11]
port 24 nsew signal tristate
flabel metal3 s 29200 7392 30000 7504 0 FreeSans 448 0 0 0 chany_bottom_out[12]
port 25 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 chany_bottom_out[13]
port 26 nsew signal tristate
flabel metal2 s 12096 29200 12208 30000 0 FreeSans 448 90 0 0 chany_bottom_out[14]
port 27 nsew signal tristate
flabel metal2 s 11424 29200 11536 30000 0 FreeSans 448 90 0 0 chany_bottom_out[15]
port 28 nsew signal tristate
flabel metal2 s 22176 29200 22288 30000 0 FreeSans 448 90 0 0 chany_bottom_out[16]
port 29 nsew signal tristate
flabel metal3 s 29200 6048 30000 6160 0 FreeSans 448 0 0 0 chany_bottom_out[17]
port 30 nsew signal tristate
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 chany_bottom_out[18]
port 31 nsew signal tristate
flabel metal3 s 29200 6720 30000 6832 0 FreeSans 448 0 0 0 chany_bottom_out[19]
port 32 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chany_bottom_out[1]
port 33 nsew signal tristate
flabel metal2 s 14784 29200 14896 30000 0 FreeSans 448 90 0 0 chany_bottom_out[2]
port 34 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 chany_bottom_out[3]
port 35 nsew signal tristate
flabel metal3 s 29200 5376 30000 5488 0 FreeSans 448 0 0 0 chany_bottom_out[4]
port 36 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 chany_bottom_out[5]
port 37 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 chany_bottom_out[6]
port 38 nsew signal tristate
flabel metal2 s 18144 29200 18256 30000 0 FreeSans 448 90 0 0 chany_bottom_out[7]
port 39 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 chany_bottom_out[8]
port 40 nsew signal tristate
flabel metal3 s 29200 17472 30000 17584 0 FreeSans 448 0 0 0 chany_bottom_out[9]
port 41 nsew signal tristate
flabel metal3 s 29200 20832 30000 20944 0 FreeSans 448 0 0 0 chany_top_in[0]
port 42 nsew signal input
flabel metal2 s 20832 29200 20944 30000 0 FreeSans 448 90 0 0 chany_top_in[10]
port 43 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 chany_top_in[11]
port 44 nsew signal input
flabel metal3 s 29200 2016 30000 2128 0 FreeSans 448 0 0 0 chany_top_in[12]
port 45 nsew signal input
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 chany_top_in[13]
port 46 nsew signal input
flabel metal2 s 6048 29200 6160 30000 0 FreeSans 448 90 0 0 chany_top_in[14]
port 47 nsew signal input
flabel metal2 s 8736 29200 8848 30000 0 FreeSans 448 90 0 0 chany_top_in[15]
port 48 nsew signal input
flabel metal2 s 18816 29200 18928 30000 0 FreeSans 448 90 0 0 chany_top_in[16]
port 49 nsew signal input
flabel metal3 s 29200 4032 30000 4144 0 FreeSans 448 0 0 0 chany_top_in[17]
port 50 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 chany_top_in[18]
port 51 nsew signal input
flabel metal3 s 29200 2688 30000 2800 0 FreeSans 448 0 0 0 chany_top_in[19]
port 52 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chany_top_in[1]
port 53 nsew signal input
flabel metal2 s 8064 29200 8176 30000 0 FreeSans 448 90 0 0 chany_top_in[2]
port 54 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 chany_top_in[3]
port 55 nsew signal input
flabel metal3 s 29200 3360 30000 3472 0 FreeSans 448 0 0 0 chany_top_in[4]
port 56 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chany_top_in[5]
port 57 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 chany_top_in[6]
port 58 nsew signal input
flabel metal2 s 17472 29200 17584 30000 0 FreeSans 448 90 0 0 chany_top_in[7]
port 59 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 chany_top_in[8]
port 60 nsew signal input
flabel metal3 s 29200 16800 30000 16912 0 FreeSans 448 0 0 0 chany_top_in[9]
port 61 nsew signal input
flabel metal2 s 10080 29200 10192 30000 0 FreeSans 448 90 0 0 chany_top_out[0]
port 62 nsew signal tristate
flabel metal2 s 22848 29200 22960 30000 0 FreeSans 448 90 0 0 chany_top_out[10]
port 63 nsew signal tristate
flabel metal2 s 10752 29200 10864 30000 0 FreeSans 448 90 0 0 chany_top_out[11]
port 64 nsew signal tristate
flabel metal3 s 29200 19488 30000 19600 0 FreeSans 448 0 0 0 chany_top_out[12]
port 65 nsew signal tristate
flabel metal3 s 29200 26208 30000 26320 0 FreeSans 448 0 0 0 chany_top_out[13]
port 66 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 chany_top_out[14]
port 67 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 chany_top_out[15]
port 68 nsew signal tristate
flabel metal3 s 29200 25536 30000 25648 0 FreeSans 448 0 0 0 chany_top_out[16]
port 69 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chany_top_out[17]
port 70 nsew signal tristate
flabel metal2 s 16800 29200 16912 30000 0 FreeSans 448 90 0 0 chany_top_out[18]
port 71 nsew signal tristate
flabel metal3 s 29200 26880 30000 26992 0 FreeSans 448 0 0 0 chany_top_out[19]
port 72 nsew signal tristate
flabel metal2 s 12768 29200 12880 30000 0 FreeSans 448 90 0 0 chany_top_out[1]
port 73 nsew signal tristate
flabel metal3 s 29200 24864 30000 24976 0 FreeSans 448 0 0 0 chany_top_out[2]
port 74 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 chany_top_out[3]
port 75 nsew signal tristate
flabel metal2 s 23520 29200 23632 30000 0 FreeSans 448 90 0 0 chany_top_out[4]
port 76 nsew signal tristate
flabel metal2 s 9408 29200 9520 30000 0 FreeSans 448 90 0 0 chany_top_out[5]
port 77 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 chany_top_out[6]
port 78 nsew signal tristate
flabel metal3 s 29200 4704 30000 4816 0 FreeSans 448 0 0 0 chany_top_out[7]
port 79 nsew signal tristate
flabel metal3 s 29200 8736 30000 8848 0 FreeSans 448 0 0 0 chany_top_out[8]
port 80 nsew signal tristate
flabel metal3 s 29200 20160 30000 20272 0 FreeSans 448 0 0 0 chany_top_out[9]
port 81 nsew signal tristate
flabel metal3 s 29200 23520 30000 23632 0 FreeSans 448 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 82 nsew signal tristate
flabel metal2 s 14112 29200 14224 30000 0 FreeSans 448 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 83 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 84 nsew signal tristate
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 pReset
port 85 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 prog_clk
port 86 nsew signal input
flabel metal2 s 21504 29200 21616 30000 0 FreeSans 448 90 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 87 nsew signal tristate
flabel metal2 s 13440 29200 13552 30000 0 FreeSans 448 90 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 88 nsew signal tristate
flabel metal3 s 29200 22848 30000 22960 0 FreeSans 448 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 89 nsew signal tristate
flabel metal4 s 4586 3076 4906 26716 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 11390 3076 11710 26716 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 18194 3076 18514 26716 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 24998 3076 25318 26716 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 7988 3076 8308 26716 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 14792 3076 15112 26716 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 21596 3076 21916 26716 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 28400 3076 28720 26716 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
rlabel metal1 14952 25872 14952 25872 0 vdd
rlabel via1 15032 26656 15032 26656 0 vss
rlabel metal2 8680 12488 8680 12488 0 _000_
rlabel metal2 6272 13944 6272 13944 0 _001_
rlabel metal2 4368 12376 4368 12376 0 _002_
rlabel metal2 5544 10976 5544 10976 0 _003_
rlabel metal2 2408 13496 2408 13496 0 _004_
rlabel metal2 4984 10136 4984 10136 0 _005_
rlabel metal2 9912 16408 9912 16408 0 _006_
rlabel metal2 6328 18200 6328 18200 0 _007_
rlabel metal2 5880 17304 5880 17304 0 _008_
rlabel metal2 2744 15064 2744 15064 0 _009_
rlabel metal2 11928 15680 11928 15680 0 _010_
rlabel metal2 12376 15064 12376 15064 0 _011_
rlabel metal2 20104 18144 20104 18144 0 _012_
rlabel metal2 19600 20552 19600 20552 0 _013_
rlabel metal2 18144 17528 18144 17528 0 _014_
rlabel metal2 16184 19208 16184 19208 0 _015_
rlabel metal2 14168 18984 14168 18984 0 _016_
rlabel metal2 12600 18256 12600 18256 0 _017_
rlabel metal2 20552 14896 20552 14896 0 _018_
rlabel metal2 16744 15680 16744 15680 0 _019_
rlabel metal2 22008 15512 22008 15512 0 _020_
rlabel metal2 24584 16856 24584 16856 0 _021_
rlabel metal2 25592 14784 25592 14784 0 _022_
rlabel metal2 24136 17864 24136 17864 0 _023_
rlabel metal2 23912 6272 23912 6272 0 _024_
rlabel metal2 24024 9184 24024 9184 0 _025_
rlabel metal2 24584 9408 24584 9408 0 _026_
rlabel metal2 25928 8792 25928 8792 0 _027_
rlabel metal3 25592 12712 25592 12712 0 _028_
rlabel metal2 24136 11984 24136 11984 0 _029_
rlabel metal2 19096 11424 19096 11424 0 _030_
rlabel metal3 18872 9576 18872 9576 0 _031_
rlabel metal2 16408 9856 16408 9856 0 _032_
rlabel metal2 15064 10304 15064 10304 0 _033_
rlabel metal2 12488 9632 12488 9632 0 _034_
rlabel metal2 12432 9128 12432 9128 0 _035_
rlabel metal2 12712 8960 12712 8960 0 _036_
rlabel metal2 4648 12432 4648 12432 0 _037_
rlabel metal2 18200 18368 18200 18368 0 _038_
rlabel metal3 24864 5992 24864 5992 0 _039_
rlabel metal2 1736 12488 1736 12488 0 ccff_head
rlabel metal3 27720 10080 27720 10080 0 ccff_tail
rlabel metal2 5432 28070 5432 28070 0 chany_bottom_in[0]
rlabel metal2 20328 26656 20328 26656 0 chany_bottom_in[10]
rlabel metal2 6776 28070 6776 28070 0 chany_bottom_in[11]
rlabel metal3 28560 18648 28560 18648 0 chany_bottom_in[12]
rlabel metal3 28378 22232 28378 22232 0 chany_bottom_in[13]
rlabel metal2 1736 4928 1736 4928 0 chany_bottom_in[14]
rlabel metal3 1302 20216 1302 20216 0 chany_bottom_in[15]
rlabel metal2 24472 26824 24472 26824 0 chany_bottom_in[16]
rlabel metal2 8568 3024 8568 3024 0 chany_bottom_in[17]
rlabel metal2 16296 25480 16296 25480 0 chany_bottom_in[18]
rlabel metal2 28280 24752 28280 24752 0 chany_bottom_in[19]
rlabel metal2 15400 25760 15400 25760 0 chany_bottom_in[1]
rlabel metal2 28168 26264 28168 26264 0 chany_bottom_in[2]
rlabel metal2 1848 26936 1848 26936 0 chany_bottom_in[3]
rlabel metal2 20440 26320 20440 26320 0 chany_bottom_in[4]
rlabel metal2 7336 26936 7336 26936 0 chany_bottom_in[5]
rlabel metal2 3416 8176 3416 8176 0 chany_bottom_in[6]
rlabel metal2 23800 2464 23800 2464 0 chany_bottom_in[7]
rlabel metal2 28168 7392 28168 7392 0 chany_bottom_in[8]
rlabel metal2 28056 21952 28056 21952 0 chany_bottom_in[9]
rlabel metal2 27776 24696 27776 24696 0 chany_bottom_out[0]
rlabel metal2 25368 25648 25368 25648 0 chany_bottom_out[10]
rlabel metal2 10136 854 10136 854 0 chany_bottom_out[11]
rlabel metal2 27720 6776 27720 6776 0 chany_bottom_out[12]
rlabel metal3 1414 7448 1414 7448 0 chany_bottom_out[13]
rlabel metal2 12152 28070 12152 28070 0 chany_bottom_out[14]
rlabel metal2 12152 25816 12152 25816 0 chany_bottom_out[15]
rlabel metal2 23240 26656 23240 26656 0 chany_bottom_out[16]
rlabel metal2 27720 5208 27720 5208 0 chany_bottom_out[17]
rlabel metal3 2254 27608 2254 27608 0 chany_bottom_out[18]
rlabel metal2 27608 5992 27608 5992 0 chany_bottom_out[19]
rlabel metal2 12152 2198 12152 2198 0 chany_bottom_out[1]
rlabel metal2 15848 26656 15848 26656 0 chany_bottom_out[2]
rlabel metal3 1414 26264 1414 26264 0 chany_bottom_out[3]
rlabel metal2 27384 4592 27384 4592 0 chany_bottom_out[4]
rlabel metal2 20888 854 20888 854 0 chany_bottom_out[5]
rlabel metal3 1358 25592 1358 25592 0 chany_bottom_out[6]
rlabel metal2 19096 26320 19096 26320 0 chany_bottom_out[7]
rlabel metal3 1470 21560 1470 21560 0 chany_bottom_out[8]
rlabel metal2 27776 15512 27776 15512 0 chany_bottom_out[9]
rlabel metal2 28168 21224 28168 21224 0 chany_top_in[0]
rlabel metal2 20888 27426 20888 27426 0 chany_top_in[10]
rlabel metal2 9576 3416 9576 3416 0 chany_top_in[11]
rlabel metal2 24584 3584 24584 3584 0 chany_top_in[12]
rlabel metal2 1736 6328 1736 6328 0 chany_top_in[13]
rlabel metal2 5992 26936 5992 26936 0 chany_top_in[14]
rlabel metal2 8680 27272 8680 27272 0 chany_top_in[15]
rlabel metal2 18872 27426 18872 27426 0 chany_top_in[16]
rlabel metal2 27496 5320 27496 5320 0 chany_top_in[17]
rlabel metal2 2408 24080 2408 24080 0 chany_top_in[18]
rlabel metal2 23128 3136 23128 3136 0 chany_top_in[19]
rlabel metal2 11704 4200 11704 4200 0 chany_top_in[1]
rlabel metal2 8008 26936 8008 26936 0 chany_top_in[2]
rlabel metal2 1736 23688 1736 23688 0 chany_top_in[3]
rlabel metal3 27090 3416 27090 3416 0 chany_top_in[4]
rlabel metal2 20216 1974 20216 1974 0 chany_top_in[5]
rlabel metal3 2086 26936 2086 26936 0 chany_top_in[6]
rlabel metal2 17528 27426 17528 27426 0 chany_top_in[7]
rlabel metal2 1736 23016 1736 23016 0 chany_top_in[8]
rlabel metal2 28168 15680 28168 15680 0 chany_top_in[9]
rlabel metal2 11144 26208 11144 26208 0 chany_top_out[0]
rlabel metal2 23576 25648 23576 25648 0 chany_top_out[10]
rlabel metal2 10808 28070 10808 28070 0 chany_top_out[11]
rlabel metal2 28056 19712 28056 19712 0 chany_top_out[12]
rlabel metal2 27608 25144 27608 25144 0 chany_top_out[13]
rlabel metal3 1358 5432 1358 5432 0 chany_top_out[14]
rlabel metal3 1526 22232 1526 22232 0 chany_top_out[15]
rlabel metal2 27720 25872 27720 25872 0 chany_top_out[16]
rlabel metal2 10808 854 10808 854 0 chany_top_out[17]
rlabel metal2 18312 26656 18312 26656 0 chany_top_out[18]
rlabel metal2 26152 25928 26152 25928 0 chany_top_out[19]
rlabel metal2 13608 26320 13608 26320 0 chany_top_out[1]
rlabel metal2 27720 25088 27720 25088 0 chany_top_out[2]
rlabel metal3 1470 24920 1470 24920 0 chany_top_out[3]
rlabel metal2 25032 26488 25032 26488 0 chany_top_out[4]
rlabel metal2 9744 27048 9744 27048 0 chany_top_out[5]
rlabel metal3 1358 6776 1358 6776 0 chany_top_out[6]
rlabel metal2 25480 4312 25480 4312 0 chany_top_out[7]
rlabel metal3 28504 8344 28504 8344 0 chany_top_out[8]
rlabel metal2 28056 20440 28056 20440 0 chany_top_out[9]
rlabel metal2 19544 15736 19544 15736 0 clknet_0_prog_clk
rlabel metal2 2352 10584 2352 10584 0 clknet_2_0__leaf_prog_clk
rlabel metal2 9632 14504 9632 14504 0 clknet_2_1__leaf_prog_clk
rlabel metal2 27160 7000 27160 7000 0 clknet_2_2__leaf_prog_clk
rlabel metal2 21448 17304 21448 17304 0 clknet_2_3__leaf_prog_clk
rlabel metal2 5544 9464 5544 9464 0 mem_left_ipin_0.DFFR_0_.Q
rlabel metal2 2632 11816 2632 11816 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal2 6272 10696 6272 10696 0 mem_left_ipin_0.DFFR_2_.Q
rlabel metal2 3528 13384 3528 13384 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal2 5432 14532 5432 14532 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal2 9240 13496 9240 13496 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal2 13944 14056 13944 14056 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal2 11144 15736 11144 15736 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal2 1960 15736 1960 15736 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal3 7000 15960 7000 15960 0 mem_left_ipin_1.DFFR_3_.Q
rlabel metal2 8456 18872 8456 18872 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal2 10808 18480 10808 18480 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal2 15512 19488 15512 19488 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal2 15176 19712 15176 19712 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal2 16968 18536 16968 18536 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal2 22232 19544 22232 19544 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal3 21448 21672 21448 21672 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal3 24864 18424 24864 18424 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal2 27272 17192 27272 17192 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal2 26376 15344 26376 15344 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal2 27160 17864 27160 17864 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal2 22344 15624 22344 15624 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal2 17528 15624 17528 15624 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal3 22064 13832 22064 13832 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal2 24920 11704 24920 11704 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal3 26712 11256 26712 11256 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal2 26600 8372 26600 8372 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal2 25592 10080 25592 10080 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal2 25368 7980 25368 7980 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal2 23128 7224 23128 7224 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal3 10584 10696 10584 10696 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal3 14448 8120 14448 8120 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal2 16296 11032 16296 11032 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal3 17808 8120 17808 8120 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal2 18984 10640 18984 10640 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal2 2072 12432 2072 12432 0 net1
rlabel metal2 8792 3360 8792 3360 0 net10
rlabel metal2 10136 18872 10136 18872 0 net100
rlabel metal2 17976 11032 17976 11032 0 net101
rlabel metal2 22568 9352 22568 9352 0 net102
rlabel metal2 21224 20776 21224 20776 0 net103
rlabel metal2 19096 15624 19096 15624 0 net104
rlabel metal2 12152 20440 12152 20440 0 net105
rlabel metal2 13944 18872 13944 18872 0 net106
rlabel metal2 5488 18424 5488 18424 0 net107
rlabel metal2 8120 14448 8120 14448 0 net108
rlabel metal2 21952 11368 21952 11368 0 net109
rlabel metal2 17192 24584 17192 24584 0 net11
rlabel metal2 17640 19544 17640 19544 0 net110
rlabel metal2 3640 16520 3640 16520 0 net111
rlabel metal2 6664 11312 6664 11312 0 net112
rlabel metal2 10024 10136 10024 10136 0 net113
rlabel metal2 22680 12712 22680 12712 0 net114
rlabel metal2 13832 10248 13832 10248 0 net115
rlabel metal2 24360 16912 24360 16912 0 net116
rlabel metal3 3416 10584 3416 10584 0 net117
rlabel metal2 21784 10528 21784 10528 0 net118
rlabel metal2 23912 18424 23912 18424 0 net119
rlabel metal2 27832 23184 27832 23184 0 net12
rlabel metal2 23352 15624 23352 15624 0 net120
rlabel metal2 23576 8316 23576 8316 0 net121
rlabel metal2 26264 7000 26264 7000 0 net122
rlabel metal2 4760 13608 4760 13608 0 net123
rlabel metal2 20776 10136 20776 10136 0 net124
rlabel metal2 12152 24584 12152 24584 0 net13
rlabel metal3 26712 23352 26712 23352 0 net14
rlabel metal2 3864 24976 3864 24976 0 net15
rlabel metal2 21448 25144 21448 25144 0 net16
rlabel metal2 11480 23632 11480 23632 0 net17
rlabel metal2 4592 6664 4592 6664 0 net18
rlabel metal2 24080 3416 24080 3416 0 net19
rlabel metal2 10808 24248 10808 24248 0 net2
rlabel metal2 23800 5600 23800 5600 0 net20
rlabel metal2 27832 22400 27832 22400 0 net21
rlabel metal3 26656 21784 26656 21784 0 net22
rlabel metal2 21000 24976 21000 24976 0 net23
rlabel metal2 10024 4256 10024 4256 0 net24
rlabel metal2 25928 4536 25928 4536 0 net25
rlabel metal3 3136 6552 3136 6552 0 net26
rlabel metal2 10696 24696 10696 24696 0 net27
rlabel metal2 10192 23912 10192 23912 0 net28
rlabel metal2 20664 24248 20664 24248 0 net29
rlabel metal2 20552 25144 20552 25144 0 net3
rlabel metal2 25480 5096 25480 5096 0 net30
rlabel metal2 2744 24248 2744 24248 0 net31
rlabel metal2 23352 4648 23352 4648 0 net32
rlabel metal3 11424 4536 11424 4536 0 net33
rlabel metal3 9632 23912 9632 23912 0 net34
rlabel metal2 5208 24248 5208 24248 0 net35
rlabel metal2 24976 4424 24976 4424 0 net36
rlabel metal2 20216 4200 20216 4200 0 net37
rlabel metal2 4200 24584 4200 24584 0 net38
rlabel metal2 17976 24584 17976 24584 0 net39
rlabel metal2 9352 24584 9352 24584 0 net4
rlabel metal2 2128 23352 2128 23352 0 net40
rlabel metal2 27832 14840 27832 14840 0 net41
rlabel metal2 2072 10528 2072 10528 0 net42
rlabel metal2 26936 10080 26936 10080 0 net43
rlabel metal2 25816 24248 25816 24248 0 net44
rlabel metal2 21224 24976 21224 24976 0 net45
rlabel metal2 10248 4704 10248 4704 0 net46
rlabel metal2 26320 4536 26320 4536 0 net47
rlabel metal2 3864 7112 3864 7112 0 net48
rlabel metal2 11032 24360 11032 24360 0 net49
rlabel metal3 26320 19096 26320 19096 0 net5
rlabel metal2 10360 24528 10360 24528 0 net50
rlabel metal2 21000 23912 21000 23912 0 net51
rlabel metal2 25648 4872 25648 4872 0 net52
rlabel metal2 4536 24920 4536 24920 0 net53
rlabel metal3 25816 5096 25816 5096 0 net54
rlabel metal2 13160 4088 13160 4088 0 net55
rlabel metal2 15288 25032 15288 25032 0 net56
rlabel metal3 3976 24808 3976 24808 0 net57
rlabel metal2 26600 3976 26600 3976 0 net58
rlabel metal2 21112 4200 21112 4200 0 net59
rlabel metal2 27104 22232 27104 22232 0 net6
rlabel metal2 4032 23800 4032 23800 0 net60
rlabel metal2 18144 23800 18144 23800 0 net61
rlabel metal2 2968 23016 2968 23016 0 net62
rlabel metal2 27048 16016 27048 16016 0 net63
rlabel metal2 10584 24304 10584 24304 0 net64
rlabel metal2 20776 24584 20776 24584 0 net65
rlabel metal2 9744 23800 9744 23800 0 net66
rlabel metal2 25032 23688 25032 23688 0 net67
rlabel metal2 26712 23688 26712 23688 0 net68
rlabel metal2 2968 6160 2968 6160 0 net69
rlabel metal2 2072 5320 2072 5320 0 net7
rlabel metal2 5768 22736 5768 22736 0 net70
rlabel metal2 26432 23352 26432 23352 0 net71
rlabel metal2 11032 3920 11032 3920 0 net72
rlabel metal2 17584 23800 17584 23800 0 net73
rlabel metal2 24360 24136 24360 24136 0 net74
rlabel metal2 12376 25032 12376 25032 0 net75
rlabel metal2 26768 25256 26768 25256 0 net76
rlabel metal2 3584 24920 3584 24920 0 net77
rlabel metal3 23128 23800 23128 23800 0 net78
rlabel metal2 11144 23352 11144 23352 0 net79
rlabel metal2 6104 22232 6104 22232 0 net8
rlabel metal2 4536 6496 4536 6496 0 net80
rlabel metal2 26152 4200 26152 4200 0 net81
rlabel metal2 24024 4760 24024 4760 0 net82
rlabel metal2 25816 22008 25816 22008 0 net83
rlabel metal2 2408 20776 2408 20776 0 net84
rlabel metal2 14168 28070 14168 28070 0 net85
rlabel metal2 27552 21784 27552 21784 0 net86
rlabel metal2 22008 26096 22008 26096 0 net87
rlabel metal2 13496 28070 13496 28070 0 net88
rlabel metal2 26824 22568 26824 22568 0 net89
rlabel metal3 25424 23240 25424 23240 0 net9
rlabel metal2 15960 18704 15960 18704 0 net90
rlabel metal2 14224 13608 14224 13608 0 net91
rlabel metal3 16800 8344 16800 8344 0 net92
rlabel metal2 10024 14056 10024 14056 0 net93
rlabel metal2 18312 14224 18312 14224 0 net94
rlabel metal2 4984 15736 4984 15736 0 net95
rlabel metal3 13888 10584 13888 10584 0 net96
rlabel metal2 21896 17976 21896 17976 0 net97
rlabel metal2 6216 13160 6216 13160 0 net98
rlabel metal2 7784 18480 7784 18480 0 net99
rlabel metal2 1848 10024 1848 10024 0 pReset
rlabel metal3 1246 18872 1246 18872 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
