magic
tech gf180mcuD
magscale 1 10
timestamp 1702148883
<< metal1 >>
rect 1344 64314 66640 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 66640 64314
rect 1344 64228 66640 64262
rect 56702 64146 56754 64158
rect 56702 64082 56754 64094
rect 1344 63530 66640 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 66640 63530
rect 1344 63444 66640 63478
rect 66222 62914 66274 62926
rect 66222 62850 66274 62862
rect 1344 62746 66640 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 66640 62746
rect 1344 62660 66640 62694
rect 1344 61962 66640 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 66640 61962
rect 1344 61876 66640 61910
rect 1344 61178 66640 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 66640 61178
rect 1344 61092 66640 61126
rect 1344 60394 66640 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 66640 60394
rect 1344 60308 66640 60342
rect 1344 59610 66640 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 66640 59610
rect 1344 59524 66640 59558
rect 1344 58826 66640 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 66640 58826
rect 1344 58740 66640 58774
rect 1344 58042 66640 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 66640 58042
rect 1344 57956 66640 57990
rect 1344 57258 66640 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 66640 57258
rect 1344 57172 66640 57206
rect 1344 56474 66640 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 66640 56474
rect 1344 56388 66640 56422
rect 1344 55690 66640 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 66640 55690
rect 1344 55604 66640 55638
rect 1344 54906 66640 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 66640 54906
rect 1344 54820 66640 54854
rect 43698 54574 43710 54626
rect 43762 54574 43774 54626
rect 42690 54350 42702 54402
rect 42754 54350 42766 54402
rect 1344 54122 66640 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 66640 54122
rect 1344 54036 66640 54070
rect 30370 53790 30382 53842
rect 30434 53790 30446 53842
rect 33618 53790 33630 53842
rect 33682 53790 33694 53842
rect 38546 53790 38558 53842
rect 38610 53790 38622 53842
rect 41346 53790 41358 53842
rect 41410 53790 41422 53842
rect 45826 53790 45838 53842
rect 45890 53790 45902 53842
rect 31378 53566 31390 53618
rect 31442 53566 31454 53618
rect 34626 53566 34638 53618
rect 34690 53566 34702 53618
rect 39554 53566 39566 53618
rect 39618 53566 39630 53618
rect 42354 53566 42366 53618
rect 42418 53566 42430 53618
rect 47058 53566 47070 53618
rect 47122 53566 47134 53618
rect 1344 53338 66640 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 66640 53338
rect 1344 53252 66640 53286
rect 32050 53006 32062 53058
rect 32114 53006 32126 53058
rect 35858 53006 35870 53058
rect 35922 53006 35934 53058
rect 38658 53006 38670 53058
rect 38722 53006 38734 53058
rect 41234 53006 41246 53058
rect 41298 53006 41310 53058
rect 45938 53006 45950 53058
rect 46002 53006 46014 53058
rect 51090 53006 51102 53058
rect 51154 53006 51166 53058
rect 31042 52782 31054 52834
rect 31106 52782 31118 52834
rect 34850 52782 34862 52834
rect 34914 52782 34926 52834
rect 37650 52782 37662 52834
rect 37714 52782 37726 52834
rect 42578 52782 42590 52834
rect 42642 52782 42654 52834
rect 44930 52782 44942 52834
rect 44994 52782 45006 52834
rect 50082 52782 50094 52834
rect 50146 52782 50158 52834
rect 1344 52554 66640 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 66640 52554
rect 1344 52468 66640 52502
rect 27234 52222 27246 52274
rect 27298 52222 27310 52274
rect 32050 52222 32062 52274
rect 32114 52222 32126 52274
rect 34402 52222 34414 52274
rect 34466 52222 34478 52274
rect 37986 52222 37998 52274
rect 38050 52222 38062 52274
rect 40786 52222 40798 52274
rect 40850 52222 40862 52274
rect 46050 52222 46062 52274
rect 46114 52222 46126 52274
rect 48626 52222 48638 52274
rect 48690 52222 48702 52274
rect 28130 51998 28142 52050
rect 28194 51998 28206 52050
rect 30706 51998 30718 52050
rect 30770 51998 30782 52050
rect 35410 51998 35422 52050
rect 35474 51998 35486 52050
rect 39106 51998 39118 52050
rect 39170 51998 39182 52050
rect 41794 51998 41806 52050
rect 41858 51998 41870 52050
rect 47170 51998 47182 52050
rect 47234 51998 47246 52050
rect 49858 51998 49870 52050
rect 49922 51998 49934 52050
rect 1344 51770 66640 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 66640 51770
rect 1344 51684 66640 51718
rect 23650 51438 23662 51490
rect 23714 51438 23726 51490
rect 28466 51438 28478 51490
rect 28530 51438 28542 51490
rect 29026 51438 29038 51490
rect 29090 51438 29102 51490
rect 37762 51438 37774 51490
rect 37826 51438 37838 51490
rect 43138 51438 43150 51490
rect 43202 51438 43214 51490
rect 45714 51438 45726 51490
rect 45778 51438 45790 51490
rect 50754 51438 50766 51490
rect 50818 51438 50830 51490
rect 53778 51438 53790 51490
rect 53842 51438 53854 51490
rect 22306 51214 22318 51266
rect 22370 51214 22382 51266
rect 27122 51214 27134 51266
rect 27186 51214 27198 51266
rect 30146 51214 30158 51266
rect 30210 51214 30222 51266
rect 36754 51214 36766 51266
rect 36818 51214 36830 51266
rect 41906 51214 41918 51266
rect 41970 51214 41982 51266
rect 44706 51214 44718 51266
rect 44770 51214 44782 51266
rect 49746 51214 49758 51266
rect 49810 51214 49822 51266
rect 52546 51214 52558 51266
rect 52610 51214 52622 51266
rect 1344 50986 66640 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 66640 50986
rect 1344 50900 66640 50934
rect 24546 50654 24558 50706
rect 24610 50654 24622 50706
rect 27570 50654 27582 50706
rect 27634 50654 27646 50706
rect 32610 50654 32622 50706
rect 32674 50654 32686 50706
rect 40002 50654 40014 50706
rect 40066 50654 40078 50706
rect 42578 50654 42590 50706
rect 42642 50654 42654 50706
rect 45826 50654 45838 50706
rect 45890 50654 45902 50706
rect 48626 50654 48638 50706
rect 48690 50654 48702 50706
rect 54002 50654 54014 50706
rect 54066 50654 54078 50706
rect 56802 50654 56814 50706
rect 56866 50654 56878 50706
rect 25330 50430 25342 50482
rect 25394 50430 25406 50482
rect 26562 50430 26574 50482
rect 26626 50430 26638 50482
rect 33954 50430 33966 50482
rect 34018 50430 34030 50482
rect 38882 50430 38894 50482
rect 38946 50430 38958 50482
rect 43922 50430 43934 50482
rect 43986 50430 43998 50482
rect 47058 50430 47070 50482
rect 47122 50430 47134 50482
rect 49634 50430 49646 50482
rect 49698 50430 49710 50482
rect 55122 50430 55134 50482
rect 55186 50430 55198 50482
rect 57810 50430 57822 50482
rect 57874 50430 57886 50482
rect 1344 50202 66640 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 66640 50202
rect 1344 50116 66640 50150
rect 45950 50034 46002 50046
rect 53902 50034 53954 50046
rect 45378 49982 45390 50034
rect 45442 49982 45454 50034
rect 53330 49982 53342 50034
rect 53394 49982 53406 50034
rect 45950 49970 46002 49982
rect 53902 49970 53954 49982
rect 23874 49870 23886 49922
rect 23938 49870 23950 49922
rect 29362 49870 29374 49922
rect 29426 49870 29438 49922
rect 32050 49870 32062 49922
rect 32114 49870 32126 49922
rect 35298 49870 35310 49922
rect 35362 49870 35374 49922
rect 36978 49870 36990 49922
rect 37042 49870 37054 49922
rect 46834 49870 46846 49922
rect 46898 49870 46910 49922
rect 54114 49870 54126 49922
rect 54178 49870 54190 49922
rect 58818 49870 58830 49922
rect 58882 49870 58894 49922
rect 42254 49810 42306 49822
rect 25442 49758 25454 49810
rect 25506 49758 25518 49810
rect 42914 49758 42926 49810
rect 42978 49758 42990 49810
rect 46386 49758 46398 49810
rect 46450 49758 46462 49810
rect 47058 49758 47070 49810
rect 47122 49758 47134 49810
rect 50306 49758 50318 49810
rect 50370 49758 50382 49810
rect 50866 49758 50878 49810
rect 50930 49758 50942 49810
rect 54338 49758 54350 49810
rect 54402 49758 54414 49810
rect 42254 49746 42306 49758
rect 26126 49698 26178 49710
rect 22530 49646 22542 49698
rect 22594 49646 22606 49698
rect 25218 49646 25230 49698
rect 25282 49646 25294 49698
rect 26126 49634 26178 49646
rect 27918 49698 27970 49710
rect 47518 49698 47570 49710
rect 49422 49698 49474 49710
rect 49982 49698 50034 49710
rect 28242 49646 28254 49698
rect 28306 49646 28318 49698
rect 31042 49646 31054 49698
rect 31106 49646 31118 49698
rect 34066 49646 34078 49698
rect 34130 49646 34142 49698
rect 38098 49646 38110 49698
rect 38162 49646 38174 49698
rect 46162 49646 46174 49698
rect 46226 49646 46238 49698
rect 47842 49646 47854 49698
rect 47906 49646 47918 49698
rect 49634 49646 49646 49698
rect 49698 49646 49710 49698
rect 27918 49634 27970 49646
rect 47518 49634 47570 49646
rect 49422 49634 49474 49646
rect 49982 49634 50034 49646
rect 55022 49698 55074 49710
rect 55022 49634 55074 49646
rect 55470 49698 55522 49710
rect 57586 49646 57598 49698
rect 57650 49646 57662 49698
rect 55470 49634 55522 49646
rect 1344 49418 66640 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 66640 49418
rect 1344 49332 66640 49366
rect 27918 49250 27970 49262
rect 27918 49186 27970 49198
rect 35198 49250 35250 49262
rect 35198 49186 35250 49198
rect 41694 49250 41746 49262
rect 41694 49186 41746 49198
rect 48638 49250 48690 49262
rect 55346 49198 55358 49250
rect 55410 49247 55422 49250
rect 55570 49247 55582 49250
rect 55410 49201 55582 49247
rect 55410 49198 55422 49201
rect 55570 49198 55582 49201
rect 55634 49198 55646 49250
rect 48638 49186 48690 49198
rect 28142 49138 28194 49150
rect 55582 49138 55634 49150
rect 19618 49086 19630 49138
rect 19682 49086 19694 49138
rect 22866 49086 22878 49138
rect 22930 49086 22942 49138
rect 49858 49086 49870 49138
rect 49922 49086 49934 49138
rect 53666 49086 53678 49138
rect 53730 49086 53742 49138
rect 56466 49086 56478 49138
rect 56530 49086 56542 49138
rect 28142 49074 28194 49086
rect 55582 49074 55634 49086
rect 31726 49026 31778 49038
rect 37998 49026 38050 49038
rect 44942 49026 44994 49038
rect 52782 49026 52834 49038
rect 24322 48974 24334 49026
rect 24386 48974 24398 49026
rect 24770 48974 24782 49026
rect 24834 48974 24846 49026
rect 32050 48974 32062 49026
rect 32114 48974 32126 49026
rect 36082 48974 36094 49026
rect 36146 48974 36158 49026
rect 38658 48974 38670 49026
rect 38722 48974 38734 49026
rect 43362 48974 43374 49026
rect 43426 48974 43438 49026
rect 45602 48974 45614 49026
rect 45666 48974 45678 49026
rect 51874 48974 51886 49026
rect 51938 48974 51950 49026
rect 31726 48962 31778 48974
rect 37998 48962 38050 48974
rect 44942 48962 44994 48974
rect 52782 48962 52834 48974
rect 29598 48914 29650 48926
rect 18498 48862 18510 48914
rect 18562 48862 18574 48914
rect 21522 48862 21534 48914
rect 21586 48862 21598 48914
rect 29250 48862 29262 48914
rect 29314 48862 29326 48914
rect 29598 48850 29650 48862
rect 30270 48914 30322 48926
rect 30270 48850 30322 48862
rect 42254 48914 42306 48926
rect 42254 48850 42306 48862
rect 42926 48914 42978 48926
rect 47854 48914 47906 48926
rect 43586 48862 43598 48914
rect 43650 48862 43662 48914
rect 50866 48862 50878 48914
rect 50930 48862 50942 48914
rect 51650 48862 51662 48914
rect 51714 48862 51726 48914
rect 54674 48862 54686 48914
rect 54738 48862 54750 48914
rect 57474 48862 57486 48914
rect 57538 48862 57550 48914
rect 42926 48850 42978 48862
rect 47854 48850 47906 48862
rect 28254 48802 28306 48814
rect 27346 48750 27358 48802
rect 27410 48750 27422 48802
rect 28254 48738 28306 48750
rect 30158 48802 30210 48814
rect 36094 48802 36146 48814
rect 42142 48802 42194 48814
rect 34402 48750 34414 48802
rect 34466 48750 34478 48802
rect 41122 48750 41134 48802
rect 41186 48750 41198 48802
rect 30158 48738 30210 48750
rect 36094 48738 36146 48750
rect 42142 48738 42194 48750
rect 42814 48802 42866 48814
rect 42814 48738 42866 48750
rect 1344 48634 66640 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 66640 48634
rect 1344 48548 66640 48582
rect 29934 48466 29986 48478
rect 29250 48414 29262 48466
rect 29314 48414 29326 48466
rect 29934 48402 29986 48414
rect 36094 48466 36146 48478
rect 40462 48466 40514 48478
rect 45390 48466 45442 48478
rect 39890 48414 39902 48466
rect 39954 48414 39966 48466
rect 44818 48414 44830 48466
rect 44882 48414 44894 48466
rect 36094 48402 36146 48414
rect 40462 48402 40514 48414
rect 45390 48402 45442 48414
rect 48638 48466 48690 48478
rect 49410 48414 49422 48466
rect 49474 48414 49486 48466
rect 48638 48402 48690 48414
rect 41246 48354 41298 48366
rect 55358 48354 55410 48366
rect 19506 48302 19518 48354
rect 19570 48302 19582 48354
rect 22642 48302 22654 48354
rect 22706 48302 22718 48354
rect 54562 48302 54574 48354
rect 54626 48302 54638 48354
rect 58818 48302 58830 48354
rect 58882 48302 58894 48354
rect 41246 48290 41298 48302
rect 55358 48290 55410 48302
rect 26462 48242 26514 48254
rect 31950 48242 32002 48254
rect 36766 48242 36818 48254
rect 41918 48242 41970 48254
rect 52334 48242 52386 48254
rect 25890 48190 25902 48242
rect 25954 48190 25966 48242
rect 26898 48190 26910 48242
rect 26962 48190 26974 48242
rect 30818 48190 30830 48242
rect 30882 48190 30894 48242
rect 33058 48190 33070 48242
rect 33122 48190 33134 48242
rect 36082 48190 36094 48242
rect 36146 48190 36158 48242
rect 37426 48190 37438 48242
rect 37490 48190 37502 48242
rect 42242 48190 42254 48242
rect 42306 48190 42318 48242
rect 45602 48190 45614 48242
rect 45666 48190 45678 48242
rect 51762 48190 51774 48242
rect 51826 48190 51838 48242
rect 26462 48178 26514 48190
rect 31950 48178 32002 48190
rect 36766 48178 36818 48190
rect 41918 48178 41970 48190
rect 52334 48178 52386 48190
rect 53118 48242 53170 48254
rect 53118 48178 53170 48190
rect 25342 48130 25394 48142
rect 32622 48130 32674 48142
rect 20850 48078 20862 48130
rect 20914 48078 20926 48130
rect 23650 48078 23662 48130
rect 23714 48078 23726 48130
rect 25666 48078 25678 48130
rect 25730 48078 25742 48130
rect 30930 48078 30942 48130
rect 30994 48078 31006 48130
rect 31602 48078 31614 48130
rect 31666 48078 31678 48130
rect 25342 48066 25394 48078
rect 32622 48066 32674 48078
rect 35422 48130 35474 48142
rect 47966 48130 48018 48142
rect 40898 48078 40910 48130
rect 40962 48078 40974 48130
rect 35422 48066 35474 48078
rect 47966 48066 48018 48078
rect 52670 48130 52722 48142
rect 53554 48078 53566 48130
rect 53618 48078 53630 48130
rect 55570 48078 55582 48130
rect 55634 48078 55646 48130
rect 57586 48078 57598 48130
rect 57650 48078 57662 48130
rect 52670 48066 52722 48078
rect 52658 47966 52670 48018
rect 52722 48015 52734 48018
rect 53106 48015 53118 48018
rect 52722 47969 53118 48015
rect 52722 47966 52734 47969
rect 53106 47966 53118 47969
rect 53170 47966 53182 48018
rect 1344 47850 66640 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 66640 47850
rect 1344 47764 66640 47798
rect 28702 47682 28754 47694
rect 28702 47618 28754 47630
rect 32734 47682 32786 47694
rect 32734 47618 32786 47630
rect 36542 47682 36594 47694
rect 36542 47618 36594 47630
rect 48414 47682 48466 47694
rect 48414 47618 48466 47630
rect 52222 47682 52274 47694
rect 52222 47618 52274 47630
rect 56254 47682 56306 47694
rect 56254 47618 56306 47630
rect 44270 47570 44322 47582
rect 19506 47518 19518 47570
rect 19570 47518 19582 47570
rect 23426 47518 23438 47570
rect 23490 47518 23502 47570
rect 40450 47518 40462 47570
rect 40514 47518 40526 47570
rect 57474 47518 57486 47570
rect 57538 47518 57550 47570
rect 44270 47506 44322 47518
rect 29038 47458 29090 47470
rect 32846 47458 32898 47470
rect 44942 47458 44994 47470
rect 48526 47458 48578 47470
rect 25106 47406 25118 47458
rect 25170 47406 25182 47458
rect 25554 47406 25566 47458
rect 25618 47406 25630 47458
rect 29698 47406 29710 47458
rect 29762 47406 29774 47458
rect 33506 47406 33518 47458
rect 33570 47406 33582 47458
rect 42242 47406 42254 47458
rect 42306 47406 42318 47458
rect 45378 47406 45390 47458
rect 45442 47406 45454 47458
rect 49186 47406 49198 47458
rect 49250 47406 49262 47458
rect 52658 47406 52670 47458
rect 52722 47406 52734 47458
rect 53106 47406 53118 47458
rect 53170 47406 53182 47458
rect 29038 47394 29090 47406
rect 32846 47394 32898 47406
rect 44942 47394 44994 47406
rect 48526 47394 48578 47406
rect 21646 47346 21698 47358
rect 22430 47346 22482 47358
rect 18610 47294 18622 47346
rect 18674 47294 18686 47346
rect 21970 47294 21982 47346
rect 22034 47294 22046 47346
rect 24658 47294 24670 47346
rect 24722 47294 24734 47346
rect 58482 47294 58494 47346
rect 58546 47294 58558 47346
rect 21646 47282 21698 47294
rect 22430 47282 22482 47294
rect 42926 47234 42978 47246
rect 56590 47234 56642 47246
rect 28130 47182 28142 47234
rect 28194 47182 28206 47234
rect 32050 47182 32062 47234
rect 32114 47182 32126 47234
rect 35858 47182 35870 47234
rect 35922 47182 35934 47234
rect 47618 47182 47630 47234
rect 47682 47182 47694 47234
rect 51538 47182 51550 47234
rect 51602 47182 51614 47234
rect 55570 47182 55582 47234
rect 55634 47182 55646 47234
rect 42926 47170 42978 47182
rect 56590 47170 56642 47182
rect 59390 47234 59442 47246
rect 59390 47170 59442 47182
rect 1344 47066 66640 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 66640 47066
rect 1344 46980 66640 47014
rect 31614 46898 31666 46910
rect 39454 46898 39506 46910
rect 44494 46898 44546 46910
rect 23874 46846 23886 46898
rect 23938 46846 23950 46898
rect 30930 46846 30942 46898
rect 30994 46846 31006 46898
rect 38882 46846 38894 46898
rect 38946 46846 38958 46898
rect 43698 46846 43710 46898
rect 43762 46846 43774 46898
rect 31614 46834 31666 46846
rect 39454 46834 39506 46846
rect 44494 46834 44546 46846
rect 44606 46898 44658 46910
rect 44606 46834 44658 46846
rect 52446 46898 52498 46910
rect 52446 46834 52498 46846
rect 40350 46786 40402 46798
rect 17714 46734 17726 46786
rect 17778 46734 17790 46786
rect 25666 46734 25678 46786
rect 25730 46734 25742 46786
rect 35410 46734 35422 46786
rect 35474 46734 35486 46786
rect 40002 46734 40014 46786
rect 40066 46734 40078 46786
rect 40350 46722 40402 46734
rect 45390 46786 45442 46798
rect 45390 46722 45442 46734
rect 51550 46786 51602 46798
rect 51550 46722 51602 46734
rect 53230 46786 53282 46798
rect 58818 46734 58830 46786
rect 58882 46734 58894 46786
rect 59378 46734 59390 46786
rect 59442 46734 59454 46786
rect 53230 46722 53282 46734
rect 28142 46674 28194 46686
rect 35982 46674 36034 46686
rect 40798 46674 40850 46686
rect 48078 46674 48130 46686
rect 20850 46622 20862 46674
rect 20914 46622 20926 46674
rect 21298 46622 21310 46674
rect 21362 46622 21374 46674
rect 28578 46622 28590 46674
rect 28642 46622 28654 46674
rect 32274 46622 32286 46674
rect 32338 46622 32350 46674
rect 36418 46622 36430 46674
rect 36482 46622 36494 46674
rect 41458 46622 41470 46674
rect 41522 46622 41534 46674
rect 47730 46622 47742 46674
rect 47794 46622 47806 46674
rect 28142 46610 28194 46622
rect 35982 46610 36034 46622
rect 40798 46610 40850 46622
rect 48078 46610 48130 46622
rect 48638 46674 48690 46686
rect 56142 46674 56194 46686
rect 49298 46622 49310 46674
rect 49362 46622 49374 46674
rect 55570 46622 55582 46674
rect 55634 46622 55646 46674
rect 59602 46622 59614 46674
rect 59666 46622 59678 46674
rect 48638 46610 48690 46622
rect 56142 46610 56194 46622
rect 56702 46562 56754 46574
rect 18834 46510 18846 46562
rect 18898 46510 18910 46562
rect 26562 46510 26574 46562
rect 26626 46510 26638 46562
rect 32498 46510 32510 46562
rect 32562 46510 32574 46562
rect 34290 46510 34302 46562
rect 34354 46510 34366 46562
rect 56702 46498 56754 46510
rect 57150 46562 57202 46574
rect 57586 46510 57598 46562
rect 57650 46510 57662 46562
rect 57150 46498 57202 46510
rect 24446 46450 24498 46462
rect 24446 46386 24498 46398
rect 52334 46450 52386 46462
rect 52334 46386 52386 46398
rect 1344 46282 66640 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 66640 46282
rect 1344 46196 66640 46230
rect 17166 46114 17218 46126
rect 17166 46050 17218 46062
rect 24894 46114 24946 46126
rect 24894 46050 24946 46062
rect 28702 46114 28754 46126
rect 28702 46050 28754 46062
rect 29038 46114 29090 46126
rect 29038 46050 29090 46062
rect 36542 46114 36594 46126
rect 36542 46050 36594 46062
rect 37438 46114 37490 46126
rect 37438 46050 37490 46062
rect 56254 46114 56306 46126
rect 56254 46050 56306 46062
rect 44942 46002 44994 46014
rect 43586 45950 43598 46002
rect 43650 45950 43662 46002
rect 57474 45950 57486 46002
rect 57538 45950 57550 46002
rect 44942 45938 44994 45950
rect 20862 45890 20914 45902
rect 20290 45838 20302 45890
rect 20354 45838 20366 45890
rect 20862 45826 20914 45838
rect 21422 45890 21474 45902
rect 32734 45890 32786 45902
rect 21746 45838 21758 45890
rect 21810 45838 21822 45890
rect 25106 45838 25118 45890
rect 25170 45838 25182 45890
rect 25554 45838 25566 45890
rect 25618 45838 25630 45890
rect 32050 45838 32062 45890
rect 32114 45838 32126 45890
rect 21422 45826 21474 45838
rect 32734 45826 32786 45838
rect 32846 45890 32898 45902
rect 40910 45890 40962 45902
rect 33394 45838 33406 45890
rect 33458 45838 33470 45890
rect 40450 45838 40462 45890
rect 40514 45838 40526 45890
rect 41794 45838 41806 45890
rect 41858 45838 41870 45890
rect 50418 45838 50430 45890
rect 50482 45838 50494 45890
rect 52658 45838 52670 45890
rect 52722 45838 52734 45890
rect 53106 45838 53118 45890
rect 53170 45838 53182 45890
rect 59266 45838 59278 45890
rect 59330 45838 59342 45890
rect 59490 45838 59502 45890
rect 59554 45838 59566 45890
rect 32846 45826 32898 45838
rect 40910 45826 40962 45838
rect 27918 45778 27970 45790
rect 27918 45714 27970 45726
rect 29822 45778 29874 45790
rect 29822 45714 29874 45726
rect 35758 45778 35810 45790
rect 35758 45714 35810 45726
rect 38222 45778 38274 45790
rect 46274 45726 46286 45778
rect 46338 45726 46350 45778
rect 58482 45726 58494 45778
rect 58546 45726 58558 45778
rect 38222 45714 38274 45726
rect 45726 45666 45778 45678
rect 17714 45614 17726 45666
rect 17778 45614 17790 45666
rect 24210 45614 24222 45666
rect 24274 45614 24286 45666
rect 45726 45602 45778 45614
rect 51886 45666 51938 45678
rect 56590 45666 56642 45678
rect 55682 45614 55694 45666
rect 55746 45614 55758 45666
rect 51886 45602 51938 45614
rect 56590 45602 56642 45614
rect 57038 45666 57090 45678
rect 57038 45602 57090 45614
rect 60622 45666 60674 45678
rect 60622 45602 60674 45614
rect 1344 45498 66640 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 66640 45498
rect 1344 45412 66640 45446
rect 24446 45330 24498 45342
rect 23650 45278 23662 45330
rect 23714 45278 23726 45330
rect 24446 45266 24498 45278
rect 32958 45330 33010 45342
rect 40462 45330 40514 45342
rect 33730 45278 33742 45330
rect 33794 45278 33806 45330
rect 39890 45278 39902 45330
rect 39954 45278 39966 45330
rect 32958 45266 33010 45278
rect 40462 45266 40514 45278
rect 41022 45330 41074 45342
rect 41022 45266 41074 45278
rect 42366 45330 42418 45342
rect 42366 45266 42418 45278
rect 47294 45330 47346 45342
rect 47294 45266 47346 45278
rect 48190 45330 48242 45342
rect 48190 45266 48242 45278
rect 52334 45330 52386 45342
rect 52334 45266 52386 45278
rect 56142 45330 56194 45342
rect 56142 45266 56194 45278
rect 43150 45218 43202 45230
rect 51550 45218 51602 45230
rect 17714 45166 17726 45218
rect 17778 45166 17790 45218
rect 18386 45166 18398 45218
rect 18450 45166 18462 45218
rect 28578 45166 28590 45218
rect 28642 45166 28654 45218
rect 32162 45166 32174 45218
rect 32226 45166 32238 45218
rect 41458 45166 41470 45218
rect 41522 45166 41534 45218
rect 46834 45166 46846 45218
rect 46898 45166 46910 45218
rect 43150 45154 43202 45166
rect 51550 45154 51602 45166
rect 55358 45218 55410 45230
rect 58818 45166 58830 45218
rect 58882 45166 58894 45218
rect 61394 45166 61406 45218
rect 61458 45166 61470 45218
rect 55358 45154 55410 45166
rect 30942 45106 30994 45118
rect 36430 45106 36482 45118
rect 17490 45054 17502 45106
rect 17554 45054 17566 45106
rect 20850 45054 20862 45106
rect 20914 45054 20926 45106
rect 21298 45054 21310 45106
rect 21362 45054 21374 45106
rect 26674 45054 26686 45106
rect 26738 45054 26750 45106
rect 32386 45054 32398 45106
rect 32450 45054 32462 45106
rect 35970 45054 35982 45106
rect 36034 45054 36046 45106
rect 30942 45042 30994 45054
rect 36430 45042 36482 45054
rect 36766 45106 36818 45118
rect 48862 45106 48914 45118
rect 37426 45054 37438 45106
rect 37490 45054 37502 45106
rect 41682 45054 41694 45106
rect 41746 45054 41758 45106
rect 45490 45054 45502 45106
rect 45554 45054 45566 45106
rect 45938 45054 45950 45106
rect 46002 45054 46014 45106
rect 49298 45054 49310 45106
rect 49362 45054 49374 45106
rect 52546 45054 52558 45106
rect 52610 45054 52622 45106
rect 52994 45054 53006 45106
rect 53058 45054 53070 45106
rect 36766 45042 36818 45054
rect 48862 45042 48914 45054
rect 16942 44994 16994 45006
rect 46510 44994 46562 45006
rect 19506 44942 19518 44994
rect 19570 44942 19582 44994
rect 16942 44930 16994 44942
rect 46510 44930 46562 44942
rect 47182 44994 47234 45006
rect 47182 44930 47234 44942
rect 56702 44994 56754 45006
rect 56702 44930 56754 44942
rect 57150 44994 57202 45006
rect 59502 44994 59554 45006
rect 57586 44942 57598 44994
rect 57650 44942 57662 44994
rect 60386 44942 60398 44994
rect 60450 44942 60462 44994
rect 57150 44930 57202 44942
rect 59502 44930 59554 44942
rect 1344 44714 66640 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 66640 44714
rect 1344 44628 66640 44662
rect 17166 44546 17218 44558
rect 17166 44482 17218 44494
rect 28030 44546 28082 44558
rect 28030 44482 28082 44494
rect 35198 44546 35250 44558
rect 35198 44482 35250 44494
rect 40574 44546 40626 44558
rect 40574 44482 40626 44494
rect 49646 44546 49698 44558
rect 49646 44482 49698 44494
rect 24110 44434 24162 44446
rect 29822 44434 29874 44446
rect 49870 44434 49922 44446
rect 51102 44434 51154 44446
rect 14802 44382 14814 44434
rect 14866 44382 14878 44434
rect 23090 44382 23102 44434
rect 23154 44382 23166 44434
rect 29474 44382 29486 44434
rect 29538 44382 29550 44434
rect 41794 44382 41806 44434
rect 41858 44382 41870 44434
rect 45154 44382 45166 44434
rect 45218 44382 45230 44434
rect 50194 44382 50206 44434
rect 50258 44382 50270 44434
rect 24110 44370 24162 44382
rect 29822 44370 29874 44382
rect 49870 44370 49922 44382
rect 51102 44370 51154 44382
rect 51438 44434 51490 44446
rect 57138 44382 57150 44434
rect 57202 44382 57214 44434
rect 58930 44382 58942 44434
rect 58994 44382 59006 44434
rect 61506 44382 61518 44434
rect 61570 44382 61582 44434
rect 51438 44370 51490 44382
rect 20862 44322 20914 44334
rect 20178 44270 20190 44322
rect 20242 44270 20254 44322
rect 20862 44258 20914 44270
rect 24558 44322 24610 44334
rect 31502 44322 31554 44334
rect 45950 44322 46002 44334
rect 24882 44270 24894 44322
rect 24946 44270 24958 44322
rect 30482 44270 30494 44322
rect 30546 44270 30558 44322
rect 32050 44270 32062 44322
rect 32114 44270 32126 44322
rect 36978 44270 36990 44322
rect 37042 44270 37054 44322
rect 37426 44270 37438 44322
rect 37490 44270 37502 44322
rect 45378 44270 45390 44322
rect 45442 44270 45454 44322
rect 46610 44270 46622 44322
rect 46674 44270 46686 44322
rect 52658 44270 52670 44322
rect 52722 44270 52734 44322
rect 58482 44270 58494 44322
rect 58546 44270 58558 44322
rect 24558 44258 24610 44270
rect 31502 44258 31554 44270
rect 45950 44258 46002 44270
rect 28254 44210 28306 44222
rect 36318 44210 36370 44222
rect 43598 44210 43650 44222
rect 59278 44210 59330 44222
rect 16146 44158 16158 44210
rect 16210 44158 16222 44210
rect 22082 44158 22094 44210
rect 22146 44158 22158 44210
rect 30258 44158 30270 44210
rect 30322 44158 30334 44210
rect 35970 44158 35982 44210
rect 36034 44158 36046 44210
rect 42802 44158 42814 44210
rect 42866 44158 42878 44210
rect 58258 44158 58270 44210
rect 58322 44158 58334 44210
rect 62514 44158 62526 44210
rect 62578 44158 62590 44210
rect 28254 44146 28306 44158
rect 36318 44146 36370 44158
rect 43598 44146 43650 44158
rect 59278 44146 59330 44158
rect 28366 44098 28418 44110
rect 40910 44098 40962 44110
rect 17714 44046 17726 44098
rect 17778 44046 17790 44098
rect 27458 44046 27470 44098
rect 27522 44046 27534 44098
rect 34626 44046 34638 44098
rect 34690 44046 34702 44098
rect 39890 44046 39902 44098
rect 39954 44046 39966 44098
rect 28366 44034 28418 44046
rect 40910 44034 40962 44046
rect 43710 44098 43762 44110
rect 50654 44098 50706 44110
rect 49074 44046 49086 44098
rect 49138 44046 49150 44098
rect 43710 44034 43762 44046
rect 50654 44034 50706 44046
rect 51550 44098 51602 44110
rect 51550 44034 51602 44046
rect 59726 44098 59778 44110
rect 59726 44034 59778 44046
rect 1344 43930 66640 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 66640 43930
rect 1344 43844 66640 43878
rect 59502 43762 59554 43774
rect 43698 43710 43710 43762
rect 43762 43710 43774 43762
rect 59502 43698 59554 43710
rect 20750 43650 20802 43662
rect 14802 43598 14814 43650
rect 14866 43598 14878 43650
rect 17714 43598 17726 43650
rect 17778 43598 17790 43650
rect 19394 43598 19406 43650
rect 19458 43598 19470 43650
rect 20750 43586 20802 43598
rect 21534 43650 21586 43662
rect 27918 43650 27970 43662
rect 25666 43598 25678 43650
rect 25730 43598 25742 43650
rect 21534 43586 21586 43598
rect 27918 43586 27970 43598
rect 28702 43650 28754 43662
rect 44494 43650 44546 43662
rect 33058 43598 33070 43650
rect 33122 43598 33134 43650
rect 34178 43598 34190 43650
rect 34242 43598 34254 43650
rect 28702 43586 28754 43598
rect 44494 43586 44546 43598
rect 47742 43650 47794 43662
rect 47742 43586 47794 43598
rect 48190 43650 48242 43662
rect 49534 43650 49586 43662
rect 49186 43598 49198 43650
rect 49250 43598 49262 43650
rect 48190 43586 48242 43598
rect 49534 43586 49586 43598
rect 50766 43650 50818 43662
rect 50766 43586 50818 43598
rect 51774 43650 51826 43662
rect 54898 43598 54910 43650
rect 54962 43598 54974 43650
rect 58818 43598 58830 43650
rect 58882 43598 58894 43650
rect 61394 43598 61406 43650
rect 61458 43598 61470 43650
rect 51774 43586 51826 43598
rect 24446 43538 24498 43550
rect 31390 43538 31442 43550
rect 50990 43538 51042 43550
rect 54686 43538 54738 43550
rect 17490 43486 17502 43538
rect 17554 43486 17566 43538
rect 23762 43486 23774 43538
rect 23826 43486 23838 43538
rect 31042 43486 31054 43538
rect 31106 43486 31118 43538
rect 32386 43486 32398 43538
rect 32450 43486 32462 43538
rect 33282 43486 33294 43538
rect 33346 43486 33358 43538
rect 36530 43486 36542 43538
rect 36594 43486 36606 43538
rect 40898 43486 40910 43538
rect 40962 43486 40974 43538
rect 41458 43486 41470 43538
rect 41522 43486 41534 43538
rect 45154 43486 45166 43538
rect 45218 43486 45230 43538
rect 49970 43486 49982 43538
rect 50034 43486 50046 43538
rect 54114 43486 54126 43538
rect 54178 43486 54190 43538
rect 55122 43486 55134 43538
rect 55186 43486 55198 43538
rect 55906 43486 55918 43538
rect 55970 43486 55982 43538
rect 24446 43474 24498 43486
rect 31390 43474 31442 43486
rect 50990 43474 51042 43486
rect 54686 43474 54738 43486
rect 27694 43426 27746 43438
rect 33854 43426 33906 43438
rect 45726 43426 45778 43438
rect 15810 43374 15822 43426
rect 15874 43374 15886 43426
rect 18050 43374 18062 43426
rect 18114 43374 18126 43426
rect 26674 43374 26686 43426
rect 26738 43374 26750 43426
rect 32162 43374 32174 43426
rect 32226 43374 32238 43426
rect 38994 43374 39006 43426
rect 39058 43374 39070 43426
rect 27694 43362 27746 43374
rect 33854 43362 33906 43374
rect 45726 43362 45778 43374
rect 48862 43426 48914 43438
rect 56702 43426 56754 43438
rect 50194 43374 50206 43426
rect 50258 43374 50270 43426
rect 55682 43374 55694 43426
rect 55746 43374 55758 43426
rect 48862 43362 48914 43374
rect 56702 43362 56754 43374
rect 57150 43426 57202 43438
rect 57586 43374 57598 43426
rect 57650 43374 57662 43426
rect 60386 43374 60398 43426
rect 60450 43374 60462 43426
rect 57150 43362 57202 43374
rect 1344 43146 66640 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 66640 43146
rect 1344 43060 66640 43094
rect 21198 42978 21250 42990
rect 17602 42926 17614 42978
rect 17666 42975 17678 42978
rect 17938 42975 17950 42978
rect 17666 42929 17950 42975
rect 17666 42926 17678 42929
rect 17938 42926 17950 42929
rect 18002 42926 18014 42978
rect 21198 42914 21250 42926
rect 32734 42978 32786 42990
rect 32734 42914 32786 42926
rect 40574 42978 40626 42990
rect 40574 42914 40626 42926
rect 44382 42978 44434 42990
rect 44382 42914 44434 42926
rect 52222 42978 52274 42990
rect 52222 42914 52274 42926
rect 60062 42978 60114 42990
rect 60062 42914 60114 42926
rect 17950 42866 18002 42878
rect 16818 42814 16830 42866
rect 16882 42814 16894 42866
rect 19506 42814 19518 42866
rect 19570 42814 19582 42866
rect 61506 42814 61518 42866
rect 61570 42814 61582 42866
rect 17950 42802 18002 42814
rect 24894 42754 24946 42766
rect 29262 42754 29314 42766
rect 32846 42754 32898 42766
rect 36878 42754 36930 42766
rect 40910 42754 40962 42766
rect 44942 42754 44994 42766
rect 52782 42754 52834 42766
rect 56590 42754 56642 42766
rect 24210 42702 24222 42754
rect 24274 42702 24286 42754
rect 28018 42702 28030 42754
rect 28082 42702 28094 42754
rect 28578 42702 28590 42754
rect 28642 42702 28654 42754
rect 29698 42702 29710 42754
rect 29762 42702 29774 42754
rect 35970 42702 35982 42754
rect 36034 42702 36046 42754
rect 36418 42702 36430 42754
rect 36482 42702 36494 42754
rect 37426 42702 37438 42754
rect 37490 42702 37502 42754
rect 41234 42702 41246 42754
rect 41298 42702 41310 42754
rect 45378 42702 45390 42754
rect 45442 42702 45454 42754
rect 48626 42702 48638 42754
rect 48690 42702 48702 42754
rect 49074 42702 49086 42754
rect 49138 42702 49150 42754
rect 53106 42702 53118 42754
rect 53170 42702 53182 42754
rect 57026 42702 57038 42754
rect 57090 42702 57102 42754
rect 24894 42690 24946 42702
rect 29262 42690 29314 42702
rect 32846 42690 32898 42702
rect 36878 42690 36930 42702
rect 40910 42690 40962 42702
rect 44942 42690 44994 42702
rect 52782 42690 52834 42702
rect 56590 42690 56642 42702
rect 25790 42642 25842 42654
rect 15922 42590 15934 42642
rect 15986 42590 15998 42642
rect 18722 42590 18734 42642
rect 18786 42590 18798 42642
rect 25790 42578 25842 42590
rect 33630 42642 33682 42654
rect 33630 42578 33682 42590
rect 48414 42642 48466 42654
rect 48414 42578 48466 42590
rect 55470 42642 55522 42654
rect 55470 42578 55522 42590
rect 56254 42642 56306 42654
rect 62514 42590 62526 42642
rect 62578 42590 62590 42642
rect 56254 42578 56306 42590
rect 25006 42530 25058 42542
rect 21970 42478 21982 42530
rect 22034 42478 22046 42530
rect 32162 42478 32174 42530
rect 32226 42478 32238 42530
rect 40002 42478 40014 42530
rect 40066 42478 40078 42530
rect 43586 42478 43598 42530
rect 43650 42478 43662 42530
rect 47618 42478 47630 42530
rect 47682 42478 47694 42530
rect 51650 42478 51662 42530
rect 51714 42478 51726 42530
rect 59378 42478 59390 42530
rect 59442 42478 59454 42530
rect 25006 42466 25058 42478
rect 1344 42362 66640 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 66640 42362
rect 1344 42276 66640 42310
rect 23090 42142 23102 42194
rect 23154 42142 23166 42194
rect 43922 42142 43934 42194
rect 43986 42142 43998 42194
rect 51538 42142 51550 42194
rect 51602 42142 51614 42194
rect 55346 42142 55358 42194
rect 55410 42142 55422 42194
rect 30606 42082 30658 42094
rect 12002 42030 12014 42082
rect 12066 42030 12078 42082
rect 16706 42030 16718 42082
rect 16770 42030 16782 42082
rect 17826 42030 17838 42082
rect 17890 42030 17902 42082
rect 30606 42018 30658 42030
rect 36654 42082 36706 42094
rect 36654 42018 36706 42030
rect 47518 42082 47570 42094
rect 58818 42030 58830 42082
rect 58882 42030 58894 42082
rect 61394 42030 61406 42082
rect 61458 42030 61470 42082
rect 47518 42018 47570 42030
rect 20302 41970 20354 41982
rect 23774 41970 23826 41982
rect 27134 41970 27186 41982
rect 27918 41970 27970 41982
rect 31390 41970 31442 41982
rect 32510 41970 32562 41982
rect 35870 41970 35922 41982
rect 39566 41970 39618 41982
rect 20626 41918 20638 41970
rect 20690 41918 20702 41970
rect 23986 41918 23998 41970
rect 24050 41918 24062 41970
rect 27458 41918 27470 41970
rect 27522 41918 27534 41970
rect 28242 41918 28254 41970
rect 28306 41918 28318 41970
rect 31714 41918 31726 41970
rect 31778 41918 31790 41970
rect 33282 41918 33294 41970
rect 33346 41918 33358 41970
rect 38882 41918 38894 41970
rect 38946 41918 38958 41970
rect 20302 41906 20354 41918
rect 23774 41906 23826 41918
rect 27134 41906 27186 41918
rect 27918 41906 27970 41918
rect 31390 41906 31442 41918
rect 32510 41906 32562 41918
rect 35870 41906 35922 41918
rect 39566 41906 39618 41918
rect 40798 41970 40850 41982
rect 44494 41970 44546 41982
rect 41458 41918 41470 41970
rect 41522 41918 41534 41970
rect 40798 41906 40850 41918
rect 44494 41906 44546 41918
rect 44830 41970 44882 41982
rect 48302 41970 48354 41982
rect 45266 41918 45278 41970
rect 45330 41918 45342 41970
rect 44830 41906 44882 41918
rect 48302 41906 48354 41918
rect 48638 41970 48690 41982
rect 52334 41970 52386 41982
rect 49298 41918 49310 41970
rect 49362 41918 49374 41970
rect 48638 41906 48690 41918
rect 52334 41906 52386 41918
rect 52446 41970 52498 41982
rect 56142 41970 56194 41982
rect 52994 41918 53006 41970
rect 53058 41918 53070 41970
rect 52446 41906 52498 41918
rect 56142 41906 56194 41918
rect 56702 41970 56754 41982
rect 56702 41906 56754 41918
rect 59502 41970 59554 41982
rect 62402 41918 62414 41970
rect 62466 41918 62478 41970
rect 59502 41906 59554 41918
rect 24334 41858 24386 41870
rect 13010 41806 13022 41858
rect 13074 41806 13086 41858
rect 15362 41806 15374 41858
rect 15426 41806 15438 41858
rect 18834 41806 18846 41858
rect 18898 41806 18910 41858
rect 24334 41794 24386 41806
rect 25454 41858 25506 41870
rect 25454 41794 25506 41806
rect 25790 41858 25842 41870
rect 26462 41858 26514 41870
rect 40126 41858 40178 41870
rect 26114 41806 26126 41858
rect 26178 41806 26190 41858
rect 26786 41806 26798 41858
rect 26850 41806 26862 41858
rect 31826 41806 31838 41858
rect 31890 41806 31902 41858
rect 39890 41806 39902 41858
rect 39954 41806 39966 41858
rect 25790 41794 25842 41806
rect 26462 41794 26514 41806
rect 40126 41794 40178 41806
rect 57150 41858 57202 41870
rect 62974 41858 63026 41870
rect 57586 41806 57598 41858
rect 57650 41806 57662 41858
rect 60386 41806 60398 41858
rect 60450 41806 60462 41858
rect 62178 41806 62190 41858
rect 62242 41806 62254 41858
rect 57150 41794 57202 41806
rect 62974 41794 63026 41806
rect 34078 41746 34130 41758
rect 34078 41682 34130 41694
rect 1344 41578 66640 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 66640 41578
rect 1344 41492 66640 41526
rect 25006 41410 25058 41422
rect 25006 41346 25058 41358
rect 35870 41410 35922 41422
rect 35870 41346 35922 41358
rect 56254 41410 56306 41422
rect 56254 41346 56306 41358
rect 24782 41298 24834 41310
rect 36094 41298 36146 41310
rect 11890 41246 11902 41298
rect 11954 41246 11966 41298
rect 16818 41246 16830 41298
rect 16882 41246 16894 41298
rect 19730 41246 19742 41298
rect 19794 41246 19806 41298
rect 24434 41246 24446 41298
rect 24498 41246 24510 41298
rect 30930 41246 30942 41298
rect 30994 41246 31006 41298
rect 24782 41234 24834 41246
rect 36094 41234 36146 41246
rect 36990 41298 37042 41310
rect 46174 41298 46226 41310
rect 46846 41298 46898 41310
rect 52110 41298 52162 41310
rect 38210 41246 38222 41298
rect 38274 41246 38286 41298
rect 43362 41246 43374 41298
rect 43426 41246 43438 41298
rect 45490 41246 45502 41298
rect 45554 41246 45566 41298
rect 46498 41246 46510 41298
rect 46562 41246 46574 41298
rect 47170 41246 47182 41298
rect 47234 41246 47246 41298
rect 51650 41246 51662 41298
rect 51714 41246 51726 41298
rect 36990 41234 37042 41246
rect 46174 41234 46226 41246
rect 46846 41234 46898 41246
rect 52110 41234 52162 41246
rect 56702 41298 56754 41310
rect 56702 41234 56754 41246
rect 57038 41298 57090 41310
rect 59614 41298 59666 41310
rect 57474 41246 57486 41298
rect 57538 41246 57550 41298
rect 59266 41246 59278 41298
rect 59330 41246 59342 41298
rect 61730 41246 61742 41298
rect 61794 41246 61806 41298
rect 57038 41234 57090 41246
rect 59614 41234 59666 41246
rect 32174 41186 32226 41198
rect 39006 41186 39058 41198
rect 42478 41186 42530 41198
rect 47630 41186 47682 41198
rect 52558 41186 52610 41198
rect 23538 41134 23550 41186
rect 23602 41134 23614 41186
rect 28018 41134 28030 41186
rect 28082 41134 28094 41186
rect 28578 41134 28590 41186
rect 28642 41134 28654 41186
rect 32722 41134 32734 41186
rect 32786 41134 32798 41186
rect 39442 41134 39454 41186
rect 39506 41134 39518 41186
rect 45714 41134 45726 41186
rect 45778 41134 45790 41186
rect 48066 41134 48078 41186
rect 48130 41134 48142 41186
rect 51426 41134 51438 41186
rect 51490 41134 51502 41186
rect 53218 41134 53230 41186
rect 53282 41134 53294 41186
rect 32174 41122 32226 41134
rect 39006 41122 39058 41134
rect 42478 41122 42530 41134
rect 47630 41122 47682 41134
rect 52558 41122 52610 41134
rect 25790 41074 25842 41086
rect 38558 41074 38610 41086
rect 43038 41074 43090 41086
rect 10770 41022 10782 41074
rect 10834 41022 10846 41074
rect 15922 41022 15934 41074
rect 15986 41022 15998 41074
rect 18722 41022 18734 41074
rect 18786 41022 18798 41074
rect 29922 41022 29934 41074
rect 29986 41022 29998 41074
rect 36418 41022 36430 41074
rect 36482 41022 36494 41074
rect 42690 41022 42702 41074
rect 42754 41022 42766 41074
rect 25790 41010 25842 41022
rect 38558 41010 38610 41022
rect 43038 41010 43090 41022
rect 43710 41074 43762 41086
rect 45166 41074 45218 41086
rect 44818 41022 44830 41074
rect 44882 41022 44894 41074
rect 58482 41022 58494 41074
rect 58546 41022 58558 41074
rect 62514 41022 62526 41074
rect 62578 41022 62590 41074
rect 43710 41010 43762 41022
rect 45166 41010 45218 41022
rect 20750 40962 20802 40974
rect 20750 40898 20802 40910
rect 22878 40962 22930 40974
rect 37102 40962 37154 40974
rect 51102 40962 51154 40974
rect 35186 40910 35198 40962
rect 35250 40910 35262 40962
rect 41682 40910 41694 40962
rect 41746 40910 41758 40962
rect 50306 40910 50318 40962
rect 50370 40910 50382 40962
rect 55682 40910 55694 40962
rect 55746 40910 55758 40962
rect 22878 40898 22930 40910
rect 37102 40898 37154 40910
rect 51102 40898 51154 40910
rect 1344 40794 66640 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 66640 40794
rect 1344 40708 66640 40742
rect 11678 40626 11730 40638
rect 16382 40626 16434 40638
rect 12226 40574 12238 40626
rect 12290 40574 12302 40626
rect 11678 40562 11730 40574
rect 16382 40562 16434 40574
rect 21086 40626 21138 40638
rect 21086 40562 21138 40574
rect 28142 40626 28194 40638
rect 32622 40626 32674 40638
rect 37214 40626 37266 40638
rect 47966 40626 48018 40638
rect 31826 40574 31838 40626
rect 31890 40574 31902 40626
rect 36418 40574 36430 40626
rect 36482 40574 36494 40626
rect 47394 40574 47406 40626
rect 47458 40574 47470 40626
rect 28142 40562 28194 40574
rect 32622 40562 32674 40574
rect 37214 40562 37266 40574
rect 47966 40562 48018 40574
rect 56142 40626 56194 40638
rect 56142 40562 56194 40574
rect 56702 40626 56754 40638
rect 56702 40562 56754 40574
rect 57150 40626 57202 40638
rect 57150 40562 57202 40574
rect 59502 40626 59554 40638
rect 59502 40562 59554 40574
rect 17838 40514 17890 40526
rect 21870 40514 21922 40526
rect 44046 40514 44098 40526
rect 18834 40462 18846 40514
rect 18898 40462 18910 40514
rect 25554 40462 25566 40514
rect 25618 40462 25630 40514
rect 26450 40462 26462 40514
rect 26514 40462 26526 40514
rect 39442 40462 39454 40514
rect 39506 40462 39518 40514
rect 42914 40462 42926 40514
rect 42978 40462 42990 40514
rect 43698 40462 43710 40514
rect 43762 40462 43774 40514
rect 17838 40450 17890 40462
rect 21870 40450 21922 40462
rect 44046 40450 44098 40462
rect 55358 40514 55410 40526
rect 58818 40462 58830 40514
rect 58882 40462 58894 40514
rect 61394 40462 61406 40514
rect 61458 40462 61470 40514
rect 55358 40450 55410 40462
rect 15150 40402 15202 40414
rect 14690 40350 14702 40402
rect 14754 40350 14766 40402
rect 15150 40338 15202 40350
rect 16494 40402 16546 40414
rect 20302 40402 20354 40414
rect 28926 40402 28978 40414
rect 33518 40402 33570 40414
rect 44494 40402 44546 40414
rect 52446 40402 52498 40414
rect 17490 40350 17502 40402
rect 17554 40350 17566 40402
rect 24098 40350 24110 40402
rect 24162 40350 24174 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 25778 40350 25790 40402
rect 25842 40350 25854 40402
rect 29474 40350 29486 40402
rect 29538 40350 29550 40402
rect 34178 40350 34190 40402
rect 34242 40350 34254 40402
rect 44930 40350 44942 40402
rect 44994 40350 45006 40402
rect 49186 40350 49198 40402
rect 49250 40350 49262 40402
rect 51986 40350 51998 40402
rect 52050 40350 52062 40402
rect 53106 40350 53118 40402
rect 53170 40350 53182 40402
rect 16494 40338 16546 40350
rect 20302 40338 20354 40350
rect 28926 40338 28978 40350
rect 33518 40338 33570 40350
rect 44494 40338 44546 40350
rect 52446 40338 52498 40350
rect 51102 40290 51154 40302
rect 19842 40238 19854 40290
rect 19906 40238 19918 40290
rect 27682 40238 27694 40290
rect 27746 40238 27758 40290
rect 38434 40238 38446 40290
rect 38498 40238 38510 40290
rect 41906 40238 41918 40290
rect 41970 40238 41982 40290
rect 52210 40238 52222 40290
rect 52274 40238 52286 40290
rect 57586 40238 57598 40290
rect 57650 40238 57662 40290
rect 60386 40238 60398 40290
rect 60450 40238 60462 40290
rect 51102 40226 51154 40238
rect 1344 40010 66640 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 66640 40010
rect 1344 39924 66640 39958
rect 17054 39842 17106 39854
rect 17054 39778 17106 39790
rect 20862 39842 20914 39854
rect 20862 39778 20914 39790
rect 27470 39842 27522 39854
rect 27470 39778 27522 39790
rect 37774 39842 37826 39854
rect 37774 39778 37826 39790
rect 48414 39842 48466 39854
rect 48414 39778 48466 39790
rect 27918 39730 27970 39742
rect 9090 39678 9102 39730
rect 9154 39678 9166 39730
rect 11890 39678 11902 39730
rect 11954 39678 11966 39730
rect 22194 39678 22206 39730
rect 22258 39678 22270 39730
rect 23090 39678 23102 39730
rect 23154 39678 23166 39730
rect 27918 39666 27970 39678
rect 28590 39730 28642 39742
rect 49198 39730 49250 39742
rect 51774 39730 51826 39742
rect 31154 39678 31166 39730
rect 31218 39678 31230 39730
rect 34738 39678 34750 39730
rect 34802 39678 34814 39730
rect 42690 39678 42702 39730
rect 42754 39678 42766 39730
rect 49634 39678 49646 39730
rect 49698 39678 49710 39730
rect 51426 39678 51438 39730
rect 51490 39678 51502 39730
rect 28590 39666 28642 39678
rect 49198 39666 49250 39678
rect 51774 39666 51826 39678
rect 57038 39730 57090 39742
rect 57922 39678 57934 39730
rect 57986 39678 57998 39730
rect 61506 39678 61518 39730
rect 61570 39678 61582 39730
rect 57038 39666 57090 39678
rect 17166 39618 17218 39630
rect 23998 39618 24050 39630
rect 41246 39618 41298 39630
rect 13458 39566 13470 39618
rect 13522 39566 13534 39618
rect 14018 39566 14030 39618
rect 14082 39566 14094 39618
rect 17714 39566 17726 39618
rect 17778 39566 17790 39618
rect 22418 39566 22430 39618
rect 22482 39566 22494 39618
rect 24322 39566 24334 39618
rect 24386 39566 24398 39618
rect 29138 39566 29150 39618
rect 29202 39566 29214 39618
rect 34962 39566 34974 39618
rect 35026 39566 35038 39618
rect 40898 39566 40910 39618
rect 40962 39566 40974 39618
rect 17166 39554 17218 39566
rect 23998 39554 24050 39566
rect 41246 39554 41298 39566
rect 44942 39618 44994 39630
rect 53006 39618 53058 39630
rect 45378 39566 45390 39618
rect 45442 39566 45454 39618
rect 53666 39566 53678 39618
rect 53730 39566 53742 39618
rect 44942 39554 44994 39566
rect 53006 39554 53058 39566
rect 16270 39506 16322 39518
rect 21646 39506 21698 39518
rect 8082 39454 8094 39506
rect 8146 39454 8158 39506
rect 10770 39454 10782 39506
rect 10834 39454 10846 39506
rect 21298 39454 21310 39506
rect 21362 39454 21374 39506
rect 16270 39442 16322 39454
rect 21646 39442 21698 39454
rect 22878 39506 22930 39518
rect 22878 39442 22930 39454
rect 26686 39506 26738 39518
rect 26686 39442 26738 39454
rect 38558 39506 38610 39518
rect 44034 39454 44046 39506
rect 44098 39454 44110 39506
rect 50866 39454 50878 39506
rect 50930 39454 50942 39506
rect 58930 39454 58942 39506
rect 58994 39454 59006 39506
rect 62514 39454 62526 39506
rect 62578 39454 62590 39506
rect 38558 39442 38610 39454
rect 28478 39394 28530 39406
rect 20178 39342 20190 39394
rect 20242 39342 20254 39394
rect 28478 39330 28530 39342
rect 37438 39394 37490 39406
rect 37438 39330 37490 39342
rect 41806 39394 41858 39406
rect 48750 39394 48802 39406
rect 47842 39342 47854 39394
rect 47906 39342 47918 39394
rect 41806 39330 41858 39342
rect 48750 39330 48802 39342
rect 52782 39394 52834 39406
rect 56702 39394 56754 39406
rect 55906 39342 55918 39394
rect 55970 39342 55982 39394
rect 52782 39330 52834 39342
rect 56702 39330 56754 39342
rect 1344 39226 66640 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 66640 39226
rect 1344 39140 66640 39174
rect 16942 39058 16994 39070
rect 16258 39006 16270 39058
rect 16322 39006 16334 39058
rect 16942 38994 16994 39006
rect 20974 39058 21026 39070
rect 20974 38994 21026 39006
rect 21086 39058 21138 39070
rect 28030 39058 28082 39070
rect 37550 39058 37602 39070
rect 44606 39058 44658 39070
rect 21858 39006 21870 39058
rect 21922 39006 21934 39058
rect 36866 39006 36878 39058
rect 36930 39006 36942 39058
rect 43922 39006 43934 39058
rect 43986 39006 43998 39058
rect 21086 38994 21138 39006
rect 28030 38994 28082 39006
rect 37550 38994 37602 39006
rect 44606 38994 44658 39006
rect 45390 39058 45442 39070
rect 53790 39058 53842 39070
rect 52434 39006 52446 39058
rect 52498 39006 52510 39058
rect 45390 38994 45442 39006
rect 53790 38994 53842 39006
rect 56702 39058 56754 39070
rect 56702 38994 56754 39006
rect 20190 38946 20242 38958
rect 6962 38894 6974 38946
rect 7026 38894 7038 38946
rect 10994 38894 11006 38946
rect 11058 38894 11070 38946
rect 20190 38882 20242 38894
rect 28814 38946 28866 38958
rect 32286 38946 32338 38958
rect 53230 38946 53282 38958
rect 31938 38894 31950 38946
rect 32002 38894 32014 38946
rect 47058 38894 47070 38946
rect 47122 38894 47134 38946
rect 55458 38894 55470 38946
rect 55522 38894 55534 38946
rect 58818 38894 58830 38946
rect 58882 38894 58894 38946
rect 61394 38894 61406 38946
rect 61458 38894 61470 38946
rect 28814 38882 28866 38894
rect 32286 38882 32338 38894
rect 53230 38882 53282 38894
rect 13470 38834 13522 38846
rect 17278 38834 17330 38846
rect 31502 38834 31554 38846
rect 13794 38782 13806 38834
rect 13858 38782 13870 38834
rect 17826 38782 17838 38834
rect 17890 38782 17902 38834
rect 24210 38782 24222 38834
rect 24274 38782 24286 38834
rect 24658 38782 24670 38834
rect 24722 38782 24734 38834
rect 27794 38782 27806 38834
rect 27858 38782 27870 38834
rect 31154 38782 31166 38834
rect 31218 38782 31230 38834
rect 13470 38770 13522 38782
rect 17278 38770 17330 38782
rect 31502 38770 31554 38782
rect 33854 38834 33906 38846
rect 40910 38834 40962 38846
rect 49534 38834 49586 38846
rect 34514 38782 34526 38834
rect 34578 38782 34590 38834
rect 40226 38782 40238 38834
rect 40290 38782 40302 38834
rect 41570 38782 41582 38834
rect 41634 38782 41646 38834
rect 50194 38782 50206 38834
rect 50258 38782 50270 38834
rect 33854 38770 33906 38782
rect 40910 38770 40962 38782
rect 49534 38770 49586 38782
rect 10222 38722 10274 38734
rect 25454 38722 25506 38734
rect 7970 38670 7982 38722
rect 8034 38670 8046 38722
rect 9986 38670 9998 38722
rect 10050 38670 10062 38722
rect 12002 38670 12014 38722
rect 12066 38670 12078 38722
rect 10222 38658 10274 38670
rect 25454 38658 25506 38670
rect 44942 38722 44994 38734
rect 47966 38722 48018 38734
rect 45826 38670 45838 38722
rect 45890 38670 45902 38722
rect 47730 38670 47742 38722
rect 47794 38670 47806 38722
rect 44942 38658 44994 38670
rect 47966 38658 48018 38670
rect 48750 38722 48802 38734
rect 48962 38670 48974 38722
rect 49026 38670 49038 38722
rect 54450 38670 54462 38722
rect 54514 38670 54526 38722
rect 57586 38670 57598 38722
rect 57650 38670 57662 38722
rect 60386 38670 60398 38722
rect 60450 38670 60462 38722
rect 48750 38658 48802 38670
rect 37998 38610 38050 38622
rect 37998 38546 38050 38558
rect 1344 38442 66640 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 66640 38442
rect 1344 38356 66640 38390
rect 27694 38274 27746 38286
rect 27694 38210 27746 38222
rect 35086 38274 35138 38286
rect 35086 38210 35138 38222
rect 42702 38274 42754 38286
rect 42702 38210 42754 38222
rect 28030 38162 28082 38174
rect 7858 38110 7870 38162
rect 7922 38110 7934 38162
rect 15810 38110 15822 38162
rect 15874 38110 15886 38162
rect 22642 38110 22654 38162
rect 22706 38110 22718 38162
rect 28030 38098 28082 38110
rect 37438 38162 37490 38174
rect 38110 38162 38162 38174
rect 37650 38110 37662 38162
rect 37714 38110 37726 38162
rect 43698 38110 43710 38162
rect 43762 38110 43774 38162
rect 56690 38110 56702 38162
rect 56754 38110 56766 38162
rect 61506 38110 61518 38162
rect 61570 38110 61582 38162
rect 37438 38098 37490 38110
rect 38110 38098 38162 38110
rect 9326 38050 9378 38062
rect 23998 38050 24050 38062
rect 31390 38050 31442 38062
rect 39230 38050 39282 38062
rect 48750 38050 48802 38062
rect 9874 37998 9886 38050
rect 9938 37998 9950 38050
rect 15026 37998 15038 38050
rect 15090 37998 15102 38050
rect 20626 37998 20638 38050
rect 20690 37998 20702 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 31938 37998 31950 38050
rect 32002 37998 32014 38050
rect 39666 37998 39678 38050
rect 39730 37998 39742 38050
rect 43138 37998 43150 38050
rect 43202 37998 43214 38050
rect 43810 37998 43822 38050
rect 43874 37998 43886 38050
rect 44818 37998 44830 38050
rect 44882 37998 44894 38050
rect 45378 37998 45390 38050
rect 45442 37998 45454 38050
rect 49186 37998 49198 38050
rect 49250 37998 49262 38050
rect 52770 37998 52782 38050
rect 52834 37998 52846 38050
rect 9326 37986 9378 37998
rect 23998 37986 24050 37998
rect 31390 37986 31442 37998
rect 39230 37986 39282 37998
rect 48750 37986 48802 37998
rect 19742 37938 19794 37950
rect 26910 37938 26962 37950
rect 31166 37938 31218 37950
rect 7074 37886 7086 37938
rect 7138 37886 7150 37938
rect 20066 37886 20078 37938
rect 20130 37886 20142 37938
rect 20402 37886 20414 37938
rect 20466 37886 20478 37938
rect 21522 37886 21534 37938
rect 21586 37886 21598 37938
rect 30818 37886 30830 37938
rect 30882 37886 30894 37938
rect 38434 37886 38446 37938
rect 38498 37886 38510 37938
rect 42914 37886 42926 37938
rect 42978 37886 42990 37938
rect 62514 37886 62526 37938
rect 62578 37886 62590 37938
rect 19742 37874 19794 37886
rect 26910 37874 26962 37886
rect 31166 37874 31218 37886
rect 13022 37826 13074 37838
rect 12450 37774 12462 37826
rect 12514 37774 12526 37826
rect 13022 37762 13074 37774
rect 23326 37826 23378 37838
rect 48414 37826 48466 37838
rect 52222 37826 52274 37838
rect 34290 37774 34302 37826
rect 34354 37774 34366 37826
rect 42130 37774 42142 37826
rect 42194 37774 42206 37826
rect 47618 37774 47630 37826
rect 47682 37774 47694 37826
rect 51426 37774 51438 37826
rect 51490 37774 51502 37826
rect 23326 37762 23378 37774
rect 48414 37762 48466 37774
rect 52222 37762 52274 37774
rect 1344 37658 66640 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 66640 37658
rect 1344 37572 66640 37606
rect 16942 37490 16994 37502
rect 20974 37490 21026 37502
rect 24782 37490 24834 37502
rect 16370 37438 16382 37490
rect 16434 37438 16446 37490
rect 20178 37438 20190 37490
rect 20242 37438 20254 37490
rect 24210 37438 24222 37490
rect 24274 37438 24286 37490
rect 16942 37426 16994 37438
rect 20974 37426 21026 37438
rect 24782 37426 24834 37438
rect 32622 37490 32674 37502
rect 32622 37426 32674 37438
rect 34302 37490 34354 37502
rect 48190 37490 48242 37502
rect 38546 37438 38558 37490
rect 38610 37438 38622 37490
rect 53106 37438 53118 37490
rect 53170 37438 53182 37490
rect 34302 37426 34354 37438
rect 48190 37426 48242 37438
rect 25566 37378 25618 37390
rect 4162 37326 4174 37378
rect 4226 37326 4238 37378
rect 6962 37326 6974 37378
rect 7026 37326 7038 37378
rect 10994 37326 11006 37378
rect 11058 37326 11070 37378
rect 25218 37326 25230 37378
rect 25282 37326 25294 37378
rect 25566 37314 25618 37326
rect 31838 37378 31890 37390
rect 31838 37314 31890 37326
rect 33406 37378 33458 37390
rect 33406 37314 33458 37326
rect 34190 37378 34242 37390
rect 34190 37314 34242 37326
rect 47294 37378 47346 37390
rect 48750 37378 48802 37390
rect 47618 37326 47630 37378
rect 47682 37326 47694 37378
rect 47294 37314 47346 37326
rect 48750 37314 48802 37326
rect 49534 37378 49586 37390
rect 56702 37378 56754 37390
rect 53890 37326 53902 37378
rect 53954 37326 53966 37378
rect 54898 37326 54910 37378
rect 54962 37326 54974 37378
rect 55794 37326 55806 37378
rect 55858 37326 55870 37378
rect 58818 37326 58830 37378
rect 58882 37326 58894 37378
rect 61394 37326 61406 37378
rect 61458 37326 61470 37378
rect 49534 37314 49586 37326
rect 56702 37314 56754 37326
rect 13246 37266 13298 37278
rect 17278 37266 17330 37278
rect 21310 37266 21362 37278
rect 28926 37266 28978 37278
rect 35646 37266 35698 37278
rect 49982 37266 50034 37278
rect 54238 37266 54290 37278
rect 13906 37214 13918 37266
rect 13970 37214 13982 37266
rect 17938 37214 17950 37266
rect 18002 37214 18014 37266
rect 21634 37214 21646 37266
rect 21698 37214 21710 37266
rect 26114 37214 26126 37266
rect 26178 37214 26190 37266
rect 29474 37214 29486 37266
rect 29538 37214 29550 37266
rect 36306 37214 36318 37266
rect 36370 37214 36382 37266
rect 41794 37214 41806 37266
rect 41858 37214 41870 37266
rect 50642 37214 50654 37266
rect 50706 37214 50718 37266
rect 54674 37214 54686 37266
rect 54738 37214 54750 37266
rect 13246 37202 13298 37214
rect 17278 37202 17330 37214
rect 21310 37202 21362 37214
rect 28926 37202 28978 37214
rect 35646 37202 35698 37214
rect 49982 37202 50034 37214
rect 54238 37202 54290 37214
rect 39678 37154 39730 37166
rect 40350 37154 40402 37166
rect 5170 37102 5182 37154
rect 5234 37102 5246 37154
rect 7970 37102 7982 37154
rect 8034 37102 8046 37154
rect 12002 37102 12014 37154
rect 12066 37102 12078 37154
rect 28018 37102 28030 37154
rect 28082 37102 28094 37154
rect 33058 37102 33070 37154
rect 33122 37102 33134 37154
rect 40114 37102 40126 37154
rect 40178 37102 40190 37154
rect 39678 37090 39730 37102
rect 40350 37090 40402 37102
rect 41358 37154 41410 37166
rect 55470 37154 55522 37166
rect 46722 37102 46734 37154
rect 46786 37102 46798 37154
rect 48962 37102 48974 37154
rect 49026 37102 49038 37154
rect 57586 37102 57598 37154
rect 57650 37102 57662 37154
rect 60386 37102 60398 37154
rect 60450 37102 60462 37154
rect 41358 37090 41410 37102
rect 55470 37090 55522 37102
rect 39342 37042 39394 37054
rect 39342 36978 39394 36990
rect 53678 37042 53730 37054
rect 53678 36978 53730 36990
rect 1344 36874 66640 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 66640 36874
rect 1344 36788 66640 36822
rect 13022 36706 13074 36718
rect 13022 36642 13074 36654
rect 27694 36706 27746 36718
rect 27694 36642 27746 36654
rect 36542 36706 36594 36718
rect 36542 36642 36594 36654
rect 41694 36706 41746 36718
rect 56254 36706 56306 36718
rect 45490 36654 45502 36706
rect 45554 36654 45566 36706
rect 41694 36642 41746 36654
rect 56254 36642 56306 36654
rect 14030 36594 14082 36606
rect 3938 36542 3950 36594
rect 4002 36542 4014 36594
rect 8082 36542 8094 36594
rect 8146 36542 8158 36594
rect 14030 36530 14082 36542
rect 19742 36594 19794 36606
rect 37326 36594 37378 36606
rect 20066 36542 20078 36594
rect 20130 36542 20142 36594
rect 22642 36542 22654 36594
rect 22706 36542 22718 36594
rect 19742 36530 19794 36542
rect 37326 36530 37378 36542
rect 42030 36594 42082 36606
rect 42030 36530 42082 36542
rect 42814 36594 42866 36606
rect 42814 36530 42866 36542
rect 43150 36594 43202 36606
rect 43150 36530 43202 36542
rect 44382 36594 44434 36606
rect 50306 36542 50318 36594
rect 50370 36542 50382 36594
rect 51426 36542 51438 36594
rect 51490 36542 51502 36594
rect 57698 36542 57710 36594
rect 57762 36542 57774 36594
rect 61506 36542 61518 36594
rect 61570 36542 61582 36594
rect 44382 36530 44434 36542
rect 9326 36482 9378 36494
rect 18622 36482 18674 36494
rect 9874 36430 9886 36482
rect 9938 36430 9950 36482
rect 14802 36430 14814 36482
rect 14866 36430 14878 36482
rect 18162 36430 18174 36482
rect 18226 36430 18238 36482
rect 9326 36418 9378 36430
rect 18622 36418 18674 36430
rect 24222 36482 24274 36494
rect 29038 36482 29090 36494
rect 32734 36482 32786 36494
rect 24546 36430 24558 36482
rect 24610 36430 24622 36482
rect 29586 36430 29598 36482
rect 29650 36430 29662 36482
rect 24222 36418 24274 36430
rect 29038 36418 29090 36430
rect 32734 36418 32786 36430
rect 33070 36482 33122 36494
rect 37774 36482 37826 36494
rect 33506 36430 33518 36482
rect 33570 36430 33582 36482
rect 33070 36418 33122 36430
rect 37774 36418 37826 36430
rect 37998 36482 38050 36494
rect 48078 36482 48130 36494
rect 52558 36482 52610 36494
rect 56590 36482 56642 36494
rect 38658 36430 38670 36482
rect 38722 36430 38734 36482
rect 47058 36430 47070 36482
rect 47122 36430 47134 36482
rect 48290 36430 48302 36482
rect 48354 36430 48366 36482
rect 51314 36430 51326 36482
rect 51378 36430 51390 36482
rect 53218 36430 53230 36482
rect 53282 36430 53294 36482
rect 37998 36418 38050 36430
rect 48078 36418 48130 36430
rect 52558 36418 52610 36430
rect 56590 36418 56642 36430
rect 1710 36370 1762 36382
rect 19518 36370 19570 36382
rect 3042 36318 3054 36370
rect 3106 36318 3118 36370
rect 7074 36318 7086 36370
rect 7138 36318 7150 36370
rect 13682 36318 13694 36370
rect 13746 36318 13758 36370
rect 14578 36318 14590 36370
rect 14642 36318 14654 36370
rect 1710 36306 1762 36318
rect 19518 36306 19570 36318
rect 20414 36370 20466 36382
rect 40910 36370 40962 36382
rect 20738 36318 20750 36370
rect 20802 36318 20814 36370
rect 21746 36318 21758 36370
rect 21810 36318 21822 36370
rect 36978 36318 36990 36370
rect 37042 36318 37054 36370
rect 43474 36318 43486 36370
rect 43538 36318 43550 36370
rect 58482 36318 58494 36370
rect 58546 36318 58558 36370
rect 62514 36318 62526 36370
rect 62578 36318 62590 36370
rect 20414 36306 20466 36318
rect 40910 36306 40962 36318
rect 2046 36258 2098 36270
rect 15150 36258 15202 36270
rect 23214 36258 23266 36270
rect 12450 36206 12462 36258
rect 12514 36206 12526 36258
rect 15922 36206 15934 36258
rect 15986 36206 15998 36258
rect 2046 36194 2098 36206
rect 15150 36194 15202 36206
rect 23214 36194 23266 36206
rect 23662 36258 23714 36270
rect 28030 36258 28082 36270
rect 27010 36206 27022 36258
rect 27074 36206 27086 36258
rect 32162 36206 32174 36258
rect 32226 36206 32238 36258
rect 35970 36206 35982 36258
rect 36034 36206 36046 36258
rect 55458 36206 55470 36258
rect 55522 36206 55534 36258
rect 23662 36194 23714 36206
rect 28030 36194 28082 36206
rect 1344 36090 66640 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 66640 36090
rect 1344 36004 66640 36038
rect 1822 35922 1874 35934
rect 1822 35858 1874 35870
rect 11454 35922 11506 35934
rect 11454 35858 11506 35870
rect 11902 35922 11954 35934
rect 19182 35922 19234 35934
rect 28366 35922 28418 35934
rect 38558 35922 38610 35934
rect 12674 35870 12686 35922
rect 12738 35870 12750 35922
rect 19730 35870 19742 35922
rect 19794 35870 19806 35922
rect 29138 35870 29150 35922
rect 29202 35870 29214 35922
rect 37762 35870 37774 35922
rect 37826 35870 37838 35922
rect 11902 35858 11954 35870
rect 19182 35858 19234 35870
rect 28366 35858 28418 35870
rect 38558 35858 38610 35870
rect 38894 35922 38946 35934
rect 44494 35922 44546 35934
rect 48302 35922 48354 35934
rect 43698 35870 43710 35922
rect 43762 35870 43774 35922
rect 47730 35870 47742 35922
rect 47794 35870 47806 35922
rect 38894 35858 38946 35870
rect 44494 35858 44546 35870
rect 48302 35858 48354 35870
rect 48862 35922 48914 35934
rect 48862 35858 48914 35870
rect 49310 35922 49362 35934
rect 56702 35922 56754 35934
rect 53666 35870 53678 35922
rect 53730 35870 53742 35922
rect 49310 35858 49362 35870
rect 56702 35858 56754 35870
rect 18174 35810 18226 35822
rect 33406 35810 33458 35822
rect 4162 35758 4174 35810
rect 4226 35758 4238 35810
rect 6962 35758 6974 35810
rect 7026 35758 7038 35810
rect 15810 35758 15822 35810
rect 15874 35758 15886 35810
rect 16482 35758 16494 35810
rect 16546 35758 16558 35810
rect 17378 35758 17390 35810
rect 17442 35758 17454 35810
rect 23426 35758 23438 35810
rect 23490 35758 23502 35810
rect 33058 35758 33070 35810
rect 33122 35758 33134 35810
rect 18174 35746 18226 35758
rect 33406 35746 33458 35758
rect 34078 35810 34130 35822
rect 34078 35746 34130 35758
rect 50318 35810 50370 35822
rect 55122 35758 55134 35810
rect 55186 35758 55198 35810
rect 58818 35758 58830 35810
rect 58882 35758 58894 35810
rect 61394 35758 61406 35810
rect 61458 35758 61470 35810
rect 50318 35746 50370 35758
rect 15374 35698 15426 35710
rect 22878 35698 22930 35710
rect 34862 35698 34914 35710
rect 41022 35698 41074 35710
rect 44830 35698 44882 35710
rect 50542 35698 50594 35710
rect 15026 35646 15038 35698
rect 15090 35646 15102 35698
rect 16034 35646 16046 35698
rect 16098 35646 16110 35698
rect 16706 35646 16718 35698
rect 16770 35646 16782 35698
rect 17602 35646 17614 35698
rect 17666 35646 17678 35698
rect 22194 35646 22206 35698
rect 22258 35646 22270 35698
rect 26002 35646 26014 35698
rect 26066 35646 26078 35698
rect 31378 35646 31390 35698
rect 31442 35646 31454 35698
rect 31938 35646 31950 35698
rect 32002 35646 32014 35698
rect 35522 35646 35534 35698
rect 35586 35646 35598 35698
rect 41458 35646 41470 35698
rect 41522 35646 41534 35698
rect 45266 35646 45278 35698
rect 45330 35646 45342 35698
rect 51090 35646 51102 35698
rect 51154 35646 51166 35698
rect 54898 35646 54910 35698
rect 54962 35646 54974 35698
rect 55570 35646 55582 35698
rect 55634 35646 55646 35698
rect 15374 35634 15426 35646
rect 22878 35634 22930 35646
rect 34862 35634 34914 35646
rect 41022 35634 41074 35646
rect 44830 35634 44882 35646
rect 50542 35634 50594 35646
rect 11342 35586 11394 35598
rect 18958 35586 19010 35598
rect 5170 35534 5182 35586
rect 5234 35534 5246 35586
rect 7970 35534 7982 35586
rect 8034 35534 8046 35586
rect 18386 35534 18398 35586
rect 18450 35534 18462 35586
rect 11342 35522 11394 35534
rect 18958 35522 19010 35534
rect 24446 35586 24498 35598
rect 32622 35586 32674 35598
rect 27794 35534 27806 35586
rect 27858 35534 27870 35586
rect 33730 35534 33742 35586
rect 33794 35534 33806 35586
rect 49970 35534 49982 35586
rect 50034 35534 50046 35586
rect 55682 35534 55694 35586
rect 55746 35534 55758 35586
rect 57586 35534 57598 35586
rect 57650 35534 57662 35586
rect 60386 35534 60398 35586
rect 60450 35534 60462 35586
rect 24446 35522 24498 35534
rect 32622 35522 32674 35534
rect 54238 35474 54290 35486
rect 54238 35410 54290 35422
rect 1344 35306 66640 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 66640 35306
rect 1344 35220 66640 35254
rect 17054 35138 17106 35150
rect 17054 35074 17106 35086
rect 56366 35138 56418 35150
rect 56366 35074 56418 35086
rect 12910 35026 12962 35038
rect 29934 35026 29986 35038
rect 37326 35026 37378 35038
rect 3826 34974 3838 35026
rect 3890 34974 3902 35026
rect 7298 34974 7310 35026
rect 7362 34974 7374 35026
rect 26338 34974 26350 35026
rect 26402 34974 26414 35026
rect 27010 34974 27022 35026
rect 27074 34974 27086 35026
rect 37090 34974 37102 35026
rect 37154 34974 37166 35026
rect 12910 34962 12962 34974
rect 29934 34962 29986 34974
rect 37326 34962 37378 34974
rect 44270 35026 44322 35038
rect 44270 34962 44322 34974
rect 46734 35026 46786 35038
rect 46734 34962 46786 34974
rect 52110 35026 52162 35038
rect 52110 34962 52162 34974
rect 56814 35026 56866 35038
rect 59390 35026 59442 35038
rect 57586 34974 57598 35026
rect 57650 34974 57662 35026
rect 61506 34974 61518 35026
rect 61570 34974 61582 35026
rect 56814 34962 56866 34974
rect 59390 34962 59442 34974
rect 8766 34914 8818 34926
rect 12238 34914 12290 34926
rect 17166 34914 17218 34926
rect 46958 34914 47010 34926
rect 52670 34914 52722 34926
rect 9090 34862 9102 34914
rect 9154 34862 9166 34914
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 13906 34862 13918 34914
rect 13970 34862 13982 34914
rect 17714 34862 17726 34914
rect 17778 34862 17790 34914
rect 22754 34862 22766 34914
rect 22818 34862 22830 34914
rect 30146 34862 30158 34914
rect 30210 34862 30222 34914
rect 37874 34862 37886 34914
rect 37938 34862 37950 34914
rect 46050 34862 46062 34914
rect 46114 34862 46126 34914
rect 47618 34862 47630 34914
rect 47682 34862 47694 34914
rect 50978 34862 50990 34914
rect 51042 34862 51054 34914
rect 53330 34862 53342 34914
rect 53394 34862 53406 34914
rect 8766 34850 8818 34862
rect 12238 34850 12290 34862
rect 17166 34850 17218 34862
rect 46958 34850 47010 34862
rect 52670 34850 52722 34862
rect 27246 34802 27298 34814
rect 3042 34750 3054 34802
rect 3106 34750 3118 34802
rect 6290 34750 6302 34802
rect 6354 34750 6366 34802
rect 12562 34750 12574 34802
rect 12626 34750 12638 34802
rect 27246 34738 27298 34750
rect 27582 34802 27634 34814
rect 45502 34802 45554 34814
rect 35186 34750 35198 34802
rect 35250 34750 35262 34802
rect 42914 34750 42926 34802
rect 42978 34750 42990 34802
rect 45154 34750 45166 34802
rect 45218 34750 45230 34802
rect 46274 34750 46286 34802
rect 46338 34750 46350 34802
rect 51202 34750 51214 34802
rect 51266 34750 51278 34802
rect 51762 34750 51774 34802
rect 51826 34750 51838 34802
rect 58818 34750 58830 34802
rect 58882 34750 58894 34802
rect 62514 34750 62526 34802
rect 62578 34750 62590 34802
rect 27582 34738 27634 34750
rect 45502 34738 45554 34750
rect 20862 34690 20914 34702
rect 11666 34638 11678 34690
rect 11730 34638 11742 34690
rect 16482 34638 16494 34690
rect 16546 34638 16558 34690
rect 20178 34638 20190 34690
rect 20242 34638 20254 34690
rect 20862 34626 20914 34638
rect 27694 34690 27746 34702
rect 27694 34626 27746 34638
rect 28366 34690 28418 34702
rect 28366 34626 28418 34638
rect 29262 34690 29314 34702
rect 29262 34626 29314 34638
rect 36542 34690 36594 34702
rect 36542 34626 36594 34638
rect 43598 34690 43650 34702
rect 50654 34690 50706 34702
rect 59502 34690 59554 34702
rect 49970 34638 49982 34690
rect 50034 34638 50046 34690
rect 55682 34638 55694 34690
rect 55746 34638 55758 34690
rect 43598 34626 43650 34638
rect 50654 34626 50706 34638
rect 59502 34626 59554 34638
rect 1344 34522 66640 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 66640 34522
rect 1344 34436 66640 34470
rect 11118 34354 11170 34366
rect 15262 34354 15314 34366
rect 20974 34354 21026 34366
rect 24782 34354 24834 34366
rect 31838 34354 31890 34366
rect 52334 34354 52386 34366
rect 56142 34354 56194 34366
rect 11890 34302 11902 34354
rect 11954 34302 11966 34354
rect 20402 34302 20414 34354
rect 20466 34302 20478 34354
rect 24210 34302 24222 34354
rect 24274 34302 24286 34354
rect 31266 34302 31278 34354
rect 31330 34302 31342 34354
rect 39890 34302 39902 34354
rect 39954 34302 39966 34354
rect 51538 34302 51550 34354
rect 51602 34302 51614 34354
rect 55346 34302 55358 34354
rect 55410 34302 55422 34354
rect 11118 34290 11170 34302
rect 15262 34290 15314 34302
rect 20974 34290 21026 34302
rect 24782 34290 24834 34302
rect 31838 34290 31890 34302
rect 52334 34290 52386 34302
rect 56142 34290 56194 34302
rect 32398 34242 32450 34254
rect 4162 34190 4174 34242
rect 4226 34190 4238 34242
rect 6962 34190 6974 34242
rect 7026 34190 7038 34242
rect 27122 34190 27134 34242
rect 27186 34190 27198 34242
rect 32050 34190 32062 34242
rect 32114 34190 32126 34242
rect 32398 34178 32450 34190
rect 33742 34242 33794 34254
rect 33742 34178 33794 34190
rect 43710 34242 43762 34254
rect 58818 34190 58830 34242
rect 58882 34190 58894 34242
rect 61394 34190 61406 34242
rect 61458 34190 61470 34242
rect 43710 34178 43762 34190
rect 17278 34130 17330 34142
rect 21086 34130 21138 34142
rect 28366 34130 28418 34142
rect 36430 34130 36482 34142
rect 14130 34078 14142 34130
rect 14194 34078 14206 34130
rect 14690 34078 14702 34130
rect 14754 34078 14766 34130
rect 17826 34078 17838 34130
rect 17890 34078 17902 34130
rect 21634 34078 21646 34130
rect 21698 34078 21710 34130
rect 25330 34078 25342 34130
rect 25394 34078 25406 34130
rect 28690 34078 28702 34130
rect 28754 34078 28766 34130
rect 36082 34078 36094 34130
rect 36146 34078 36158 34130
rect 17278 34066 17330 34078
rect 21086 34066 21138 34078
rect 28366 34066 28418 34078
rect 36430 34066 36482 34078
rect 36766 34130 36818 34142
rect 41022 34130 41074 34142
rect 48862 34130 48914 34142
rect 52446 34130 52498 34142
rect 37426 34078 37438 34130
rect 37490 34078 37502 34130
rect 41458 34078 41470 34130
rect 41522 34078 41534 34130
rect 45602 34078 45614 34130
rect 45666 34078 45678 34130
rect 49298 34078 49310 34130
rect 49362 34078 49374 34130
rect 53106 34078 53118 34130
rect 53170 34078 53182 34130
rect 36766 34066 36818 34078
rect 41022 34066 41074 34078
rect 48862 34066 48914 34078
rect 52446 34066 52498 34078
rect 9998 34018 10050 34030
rect 10558 34018 10610 34030
rect 5170 33966 5182 34018
rect 5234 33966 5246 34018
rect 7970 33966 7982 34018
rect 8034 33966 8046 34018
rect 10210 33966 10222 34018
rect 10274 33966 10286 34018
rect 9998 33954 10050 33966
rect 10558 33954 10610 33966
rect 15822 34018 15874 34030
rect 15822 33954 15874 33966
rect 16270 34018 16322 34030
rect 16830 34018 16882 34030
rect 16482 33966 16494 34018
rect 16546 33966 16558 34018
rect 16270 33954 16322 33966
rect 16830 33954 16882 33966
rect 44494 34018 44546 34030
rect 45054 34018 45106 34030
rect 44706 33966 44718 34018
rect 44770 33966 44782 34018
rect 44494 33954 44546 33966
rect 45054 33954 45106 33966
rect 56814 34018 56866 34030
rect 57586 33966 57598 34018
rect 57650 33966 57662 34018
rect 60386 33966 60398 34018
rect 60450 33966 60462 34018
rect 56814 33954 56866 33966
rect 32958 33906 33010 33918
rect 32958 33842 33010 33854
rect 40462 33906 40514 33918
rect 40462 33842 40514 33854
rect 47966 33906 48018 33918
rect 47966 33842 48018 33854
rect 1344 33738 66640 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 66640 33738
rect 1344 33652 66640 33686
rect 9102 33570 9154 33582
rect 9102 33506 9154 33518
rect 15934 33570 15986 33582
rect 15934 33506 15986 33518
rect 13806 33458 13858 33470
rect 22206 33458 22258 33470
rect 35086 33458 35138 33470
rect 4050 33406 4062 33458
rect 4114 33406 4126 33458
rect 7858 33406 7870 33458
rect 7922 33406 7934 33458
rect 13458 33406 13470 33458
rect 13522 33406 13534 33458
rect 21410 33406 21422 33458
rect 21474 33406 21486 33458
rect 34290 33406 34302 33458
rect 34354 33406 34366 33458
rect 13806 33394 13858 33406
rect 22206 33394 22258 33406
rect 35086 33394 35138 33406
rect 35646 33458 35698 33470
rect 43262 33458 43314 33470
rect 42914 33406 42926 33458
rect 42978 33406 42990 33458
rect 35646 33394 35698 33406
rect 43262 33394 43314 33406
rect 43934 33458 43986 33470
rect 43934 33394 43986 33406
rect 52782 33458 52834 33470
rect 53666 33406 53678 33458
rect 53730 33406 53742 33458
rect 56466 33406 56478 33458
rect 56530 33406 56542 33458
rect 61506 33406 61518 33458
rect 61570 33406 61582 33458
rect 52782 33394 52834 33406
rect 12574 33346 12626 33358
rect 17166 33346 17218 33358
rect 30606 33346 30658 33358
rect 44718 33346 44770 33358
rect 48526 33346 48578 33358
rect 12114 33294 12126 33346
rect 12178 33294 12190 33346
rect 16706 33294 16718 33346
rect 16770 33294 16782 33346
rect 17714 33294 17726 33346
rect 17778 33294 17790 33346
rect 22530 33294 22542 33346
rect 22594 33294 22606 33346
rect 22754 33294 22766 33346
rect 22818 33294 22830 33346
rect 28466 33294 28478 33346
rect 28530 33294 28542 33346
rect 30930 33294 30942 33346
rect 30994 33294 31006 33346
rect 34514 33294 34526 33346
rect 34578 33294 34590 33346
rect 36082 33294 36094 33346
rect 36146 33294 36158 33346
rect 38546 33294 38558 33346
rect 38610 33294 38622 33346
rect 45378 33294 45390 33346
rect 45442 33294 45454 33346
rect 49186 33294 49198 33346
rect 49250 33294 49262 33346
rect 12574 33282 12626 33294
rect 17166 33282 17218 33294
rect 30606 33282 30658 33294
rect 44718 33282 44770 33294
rect 48526 33282 48578 33294
rect 9886 33234 9938 33246
rect 3042 33182 3054 33234
rect 3106 33182 3118 33234
rect 6626 33182 6638 33234
rect 6690 33182 6702 33234
rect 9886 33170 9938 33182
rect 21646 33234 21698 33246
rect 30158 33234 30210 33246
rect 47630 33234 47682 33246
rect 23538 33182 23550 33234
rect 23602 33182 23614 33234
rect 29810 33182 29822 33234
rect 29874 33182 29886 33234
rect 35858 33182 35870 33234
rect 35922 33182 35934 33234
rect 40338 33182 40350 33234
rect 40402 33182 40414 33234
rect 54674 33182 54686 33234
rect 54738 33182 54750 33234
rect 57474 33182 57486 33234
rect 57538 33182 57550 33234
rect 62514 33182 62526 33234
rect 62578 33182 62590 33234
rect 21646 33170 21698 33182
rect 30158 33170 30210 33182
rect 47630 33170 47682 33182
rect 8878 33122 8930 33134
rect 20862 33122 20914 33134
rect 34078 33122 34130 33134
rect 20290 33070 20302 33122
rect 20354 33070 20366 33122
rect 33506 33070 33518 33122
rect 33570 33070 33582 33122
rect 8878 33058 8930 33070
rect 20862 33058 20914 33070
rect 34078 33058 34130 33070
rect 43822 33122 43874 33134
rect 43822 33058 43874 33070
rect 48414 33122 48466 33134
rect 52222 33122 52274 33134
rect 51650 33070 51662 33122
rect 51714 33070 51726 33122
rect 48414 33058 48466 33070
rect 52222 33058 52274 33070
rect 1344 32954 66640 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 66640 32954
rect 1344 32868 66640 32902
rect 16158 32786 16210 32798
rect 41134 32786 41186 32798
rect 44942 32786 44994 32798
rect 29474 32734 29486 32786
rect 29538 32734 29550 32786
rect 39890 32734 39902 32786
rect 39954 32734 39966 32786
rect 44370 32734 44382 32786
rect 44434 32734 44446 32786
rect 16158 32722 16210 32734
rect 41134 32722 41186 32734
rect 44942 32722 44994 32734
rect 15374 32674 15426 32686
rect 33742 32674 33794 32686
rect 4162 32622 4174 32674
rect 4226 32622 4238 32674
rect 6962 32622 6974 32674
rect 7026 32622 7038 32674
rect 24322 32622 24334 32674
rect 24386 32622 24398 32674
rect 27234 32622 27246 32674
rect 27298 32622 27310 32674
rect 47170 32622 47182 32674
rect 47234 32622 47246 32674
rect 50754 32622 50766 32674
rect 50818 32622 50830 32674
rect 53778 32622 53790 32674
rect 53842 32622 53854 32674
rect 58818 32622 58830 32674
rect 58882 32622 58894 32674
rect 61394 32622 61406 32674
rect 61458 32622 61470 32674
rect 15374 32610 15426 32622
rect 33742 32610 33794 32622
rect 9102 32562 9154 32574
rect 28478 32562 28530 32574
rect 32398 32562 32450 32574
rect 36766 32562 36818 32574
rect 41246 32562 41298 32574
rect 45390 32562 45442 32574
rect 9874 32510 9886 32562
rect 9938 32510 9950 32562
rect 12562 32510 12574 32562
rect 12626 32510 12638 32562
rect 13010 32510 13022 32562
rect 13074 32510 13086 32562
rect 18386 32510 18398 32562
rect 18450 32510 18462 32562
rect 23762 32510 23774 32562
rect 23826 32510 23838 32562
rect 25890 32510 25902 32562
rect 25954 32510 25966 32562
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 36082 32510 36094 32562
rect 36146 32510 36158 32562
rect 36530 32510 36542 32562
rect 36594 32510 36606 32562
rect 37426 32510 37438 32562
rect 37490 32510 37502 32562
rect 41906 32510 41918 32562
rect 41970 32510 41982 32562
rect 9102 32498 9154 32510
rect 28478 32498 28530 32510
rect 32398 32498 32450 32510
rect 36766 32498 36818 32510
rect 41246 32498 41298 32510
rect 45390 32498 45442 32510
rect 48078 32562 48130 32574
rect 54562 32510 54574 32562
rect 54626 32510 54638 32562
rect 48078 32498 48130 32510
rect 16830 32450 16882 32462
rect 23326 32450 23378 32462
rect 24670 32450 24722 32462
rect 5170 32398 5182 32450
rect 5234 32398 5246 32450
rect 7970 32398 7982 32450
rect 8034 32398 8046 32450
rect 16482 32398 16494 32450
rect 16546 32398 16558 32450
rect 19506 32398 19518 32450
rect 19570 32398 19582 32450
rect 22978 32398 22990 32450
rect 23042 32398 23054 32450
rect 23874 32398 23886 32450
rect 23938 32398 23950 32450
rect 16830 32386 16882 32398
rect 23326 32386 23378 32398
rect 24670 32386 24722 32398
rect 45726 32450 45778 32462
rect 48862 32450 48914 32462
rect 46162 32398 46174 32450
rect 46226 32398 46238 32450
rect 45726 32386 45778 32398
rect 48862 32386 48914 32398
rect 49310 32450 49362 32462
rect 52222 32450 52274 32462
rect 49746 32398 49758 32450
rect 49810 32398 49822 32450
rect 52546 32398 52558 32450
rect 52610 32398 52622 32450
rect 54450 32398 54462 32450
rect 54514 32398 54526 32450
rect 57586 32398 57598 32450
rect 57650 32398 57662 32450
rect 60386 32398 60398 32450
rect 60450 32398 60462 32450
rect 49310 32386 49362 32398
rect 52222 32386 52274 32398
rect 10670 32338 10722 32350
rect 10670 32274 10722 32286
rect 28702 32338 28754 32350
rect 28702 32274 28754 32286
rect 32958 32338 33010 32350
rect 32958 32274 33010 32286
rect 40462 32338 40514 32350
rect 40462 32274 40514 32286
rect 1344 32170 66640 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 66640 32170
rect 1344 32084 66640 32118
rect 9102 31890 9154 31902
rect 4050 31838 4062 31890
rect 4114 31838 4126 31890
rect 7858 31838 7870 31890
rect 7922 31838 7934 31890
rect 9102 31826 9154 31838
rect 13022 31890 13074 31902
rect 13022 31826 13074 31838
rect 17054 31890 17106 31902
rect 17054 31826 17106 31838
rect 21198 31890 21250 31902
rect 43262 31890 43314 31902
rect 51438 31890 51490 31902
rect 36978 31838 36990 31890
rect 37042 31838 37054 31890
rect 42914 31838 42926 31890
rect 42978 31838 42990 31890
rect 49634 31838 49646 31890
rect 49698 31838 49710 31890
rect 57474 31838 57486 31890
rect 57538 31838 57550 31890
rect 61506 31838 61518 31890
rect 61570 31838 61582 31890
rect 64306 31838 64318 31890
rect 64370 31838 64382 31890
rect 21198 31826 21250 31838
rect 43262 31826 43314 31838
rect 51438 31826 51490 31838
rect 13358 31778 13410 31790
rect 17166 31778 17218 31790
rect 24670 31778 24722 31790
rect 29262 31778 29314 31790
rect 36542 31778 36594 31790
rect 9426 31726 9438 31778
rect 9490 31726 9502 31778
rect 9874 31726 9886 31778
rect 9938 31726 9950 31778
rect 13906 31726 13918 31778
rect 13970 31726 13982 31778
rect 17714 31726 17726 31778
rect 17778 31726 17790 31778
rect 24210 31726 24222 31778
rect 24274 31726 24286 31778
rect 28130 31726 28142 31778
rect 28194 31726 28206 31778
rect 28578 31726 28590 31778
rect 28642 31726 28654 31778
rect 29698 31726 29710 31778
rect 29762 31726 29774 31778
rect 32946 31726 32958 31778
rect 33010 31726 33022 31778
rect 33394 31726 33406 31778
rect 33458 31726 33470 31778
rect 13358 31714 13410 31726
rect 17166 31714 17218 31726
rect 24670 31714 24722 31726
rect 29262 31714 29314 31726
rect 36542 31714 36594 31726
rect 38222 31778 38274 31790
rect 42254 31778 42306 31790
rect 44718 31778 44770 31790
rect 52782 31778 52834 31790
rect 38658 31726 38670 31778
rect 38722 31726 38734 31778
rect 42690 31726 42702 31778
rect 42754 31726 42766 31778
rect 44146 31726 44158 31778
rect 44210 31726 44222 31778
rect 45378 31726 45390 31778
rect 45442 31726 45454 31778
rect 53218 31726 53230 31778
rect 53282 31726 53294 31778
rect 38222 31714 38274 31726
rect 42254 31714 42306 31726
rect 44718 31714 44770 31726
rect 52782 31714 52834 31726
rect 20078 31666 20130 31678
rect 3042 31614 3054 31666
rect 3106 31614 3118 31666
rect 7074 31614 7086 31666
rect 7138 31614 7150 31666
rect 20078 31602 20130 31614
rect 20862 31666 20914 31678
rect 20862 31602 20914 31614
rect 21982 31666 22034 31678
rect 21982 31602 22034 31614
rect 25790 31666 25842 31678
rect 25790 31602 25842 31614
rect 37326 31666 37378 31678
rect 37326 31602 37378 31614
rect 41694 31666 41746 31678
rect 41906 31614 41918 31666
rect 41970 31614 41982 31666
rect 43922 31614 43934 31666
rect 43986 31614 43998 31666
rect 50866 31614 50878 31666
rect 50930 31614 50942 31666
rect 58482 31614 58494 31666
rect 58546 31614 58558 31666
rect 62514 31614 62526 31666
rect 62578 31614 62590 31666
rect 65538 31614 65550 31666
rect 65602 31614 65614 31666
rect 41694 31602 41746 31614
rect 8654 31554 8706 31566
rect 25006 31554 25058 31566
rect 32734 31554 32786 31566
rect 37774 31554 37826 31566
rect 43374 31554 43426 31566
rect 48414 31554 48466 31566
rect 12338 31502 12350 31554
rect 12402 31502 12414 31554
rect 16482 31502 16494 31554
rect 16546 31502 16558 31554
rect 32050 31502 32062 31554
rect 32114 31502 32126 31554
rect 35858 31502 35870 31554
rect 35922 31502 35934 31554
rect 41122 31502 41134 31554
rect 41186 31502 41198 31554
rect 47842 31502 47854 31554
rect 47906 31502 47918 31554
rect 8654 31490 8706 31502
rect 25006 31490 25058 31502
rect 32734 31490 32786 31502
rect 37774 31490 37826 31502
rect 43374 31490 43426 31502
rect 48414 31490 48466 31502
rect 48750 31554 48802 31566
rect 48750 31490 48802 31502
rect 49198 31554 49250 31566
rect 49198 31490 49250 31502
rect 51550 31554 51602 31566
rect 56254 31554 56306 31566
rect 55682 31502 55694 31554
rect 55746 31502 55758 31554
rect 51550 31490 51602 31502
rect 56254 31490 56306 31502
rect 56590 31554 56642 31566
rect 56590 31490 56642 31502
rect 57038 31554 57090 31566
rect 57038 31490 57090 31502
rect 1344 31386 66640 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 66640 31386
rect 1344 31300 66640 31334
rect 8878 31218 8930 31230
rect 13134 31218 13186 31230
rect 17838 31218 17890 31230
rect 23998 31218 24050 31230
rect 12450 31166 12462 31218
rect 12514 31166 12526 31218
rect 16370 31166 16382 31218
rect 16434 31166 16446 31218
rect 22530 31166 22542 31218
rect 22594 31166 22606 31218
rect 8878 31154 8930 31166
rect 13134 31154 13186 31166
rect 17838 31154 17890 31166
rect 23998 31154 24050 31166
rect 25454 31218 25506 31230
rect 39902 31218 39954 31230
rect 48302 31218 48354 31230
rect 36082 31166 36094 31218
rect 36146 31166 36158 31218
rect 43698 31166 43710 31218
rect 43762 31166 43774 31218
rect 47730 31166 47742 31218
rect 47794 31166 47806 31218
rect 25454 31154 25506 31166
rect 39902 31154 39954 31166
rect 48302 31154 48354 31166
rect 56142 31218 56194 31230
rect 60510 31218 60562 31230
rect 59490 31166 59502 31218
rect 59554 31166 59566 31218
rect 56142 31154 56194 31166
rect 60510 31154 60562 31166
rect 5182 31106 5234 31118
rect 2146 31054 2158 31106
rect 2210 31054 2222 31106
rect 5182 31042 5234 31054
rect 8990 31106 9042 31118
rect 8990 31042 9042 31054
rect 16942 31106 16994 31118
rect 16942 31042 16994 31054
rect 17726 31106 17778 31118
rect 17726 31042 17778 31054
rect 26686 31106 26738 31118
rect 26686 31042 26738 31054
rect 51550 31106 51602 31118
rect 51550 31042 51602 31054
rect 55358 31106 55410 31118
rect 62402 31054 62414 31106
rect 62466 31054 62478 31106
rect 55358 31042 55410 31054
rect 9438 30994 9490 31006
rect 13246 30994 13298 31006
rect 19518 30994 19570 31006
rect 32958 30994 33010 31006
rect 39790 30994 39842 31006
rect 7522 30942 7534 30994
rect 7586 30942 7598 30994
rect 7970 30942 7982 30994
rect 8034 30942 8046 30994
rect 10098 30942 10110 30994
rect 10162 30942 10174 30994
rect 13794 30942 13806 30994
rect 13858 30942 13870 30994
rect 20178 30942 20190 30994
rect 20242 30942 20254 30994
rect 27122 30942 27134 30994
rect 27186 30942 27198 30994
rect 33618 30942 33630 30994
rect 33682 30942 33694 30994
rect 37314 30942 37326 30994
rect 37378 30942 37390 30994
rect 9438 30930 9490 30942
rect 13246 30930 13298 30942
rect 19518 30930 19570 30942
rect 32958 30930 33010 30942
rect 39790 30930 39842 30942
rect 41022 30994 41074 31006
rect 52670 30994 52722 31006
rect 56478 30994 56530 31006
rect 60174 30994 60226 31006
rect 66110 30994 66162 31006
rect 41458 30942 41470 30994
rect 41522 30942 41534 30994
rect 44706 30942 44718 30994
rect 44770 30942 44782 30994
rect 45154 30942 45166 30994
rect 45218 30942 45230 30994
rect 48738 30942 48750 30994
rect 48802 30942 48814 30994
rect 49298 30942 49310 30994
rect 49362 30942 49374 30994
rect 53106 30942 53118 30994
rect 53170 30942 53182 30994
rect 57138 30942 57150 30994
rect 57202 30942 57214 30994
rect 64978 30942 64990 30994
rect 65042 30942 65054 30994
rect 41022 30930 41074 30942
rect 52670 30930 52722 30942
rect 56478 30930 56530 30942
rect 60174 30930 60226 30942
rect 66110 30930 66162 30942
rect 18510 30882 18562 30894
rect 3154 30830 3166 30882
rect 3218 30830 3230 30882
rect 18510 30818 18562 30830
rect 19294 30882 19346 30894
rect 19294 30818 19346 30830
rect 23550 30882 23602 30894
rect 23550 30818 23602 30830
rect 26014 30882 26066 30894
rect 26338 30830 26350 30882
rect 26402 30830 26414 30882
rect 32162 30830 32174 30882
rect 32226 30830 32238 30882
rect 61394 30830 61406 30882
rect 61458 30830 61470 30882
rect 26014 30818 26066 30830
rect 4398 30770 4450 30782
rect 4398 30706 4450 30718
rect 23214 30770 23266 30782
rect 23214 30706 23266 30718
rect 36654 30770 36706 30782
rect 44494 30770 44546 30782
rect 38322 30718 38334 30770
rect 38386 30718 38398 30770
rect 36654 30706 36706 30718
rect 44494 30706 44546 30718
rect 52334 30770 52386 30782
rect 52334 30706 52386 30718
rect 1344 30602 66640 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 66640 30602
rect 1344 30516 66640 30550
rect 14702 30322 14754 30334
rect 4050 30270 4062 30322
rect 4114 30270 4126 30322
rect 7074 30270 7086 30322
rect 7138 30270 7150 30322
rect 12450 30270 12462 30322
rect 12514 30270 12526 30322
rect 14702 30258 14754 30270
rect 15038 30322 15090 30334
rect 15038 30258 15090 30270
rect 19630 30322 19682 30334
rect 50766 30322 50818 30334
rect 21410 30270 21422 30322
rect 21474 30270 21486 30322
rect 22530 30270 22542 30322
rect 22594 30270 22606 30322
rect 55458 30270 55470 30322
rect 55522 30270 55534 30322
rect 61506 30270 61518 30322
rect 61570 30270 61582 30322
rect 19630 30258 19682 30270
rect 50766 30258 50818 30270
rect 4510 30210 4562 30222
rect 4510 30146 4562 30158
rect 8318 30210 8370 30222
rect 12014 30210 12066 30222
rect 14030 30210 14082 30222
rect 19070 30210 19122 30222
rect 11330 30158 11342 30210
rect 11394 30158 11406 30210
rect 13682 30158 13694 30210
rect 13746 30158 13758 30210
rect 15362 30158 15374 30210
rect 15426 30158 15438 30210
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 8318 30146 8370 30158
rect 12014 30146 12066 30158
rect 14030 30146 14082 30158
rect 19070 30146 19122 30158
rect 20302 30210 20354 30222
rect 20302 30146 20354 30158
rect 20750 30210 20802 30222
rect 20750 30146 20802 30158
rect 21646 30210 21698 30222
rect 21646 30146 21698 30158
rect 22318 30210 22370 30222
rect 27246 30210 27298 30222
rect 26674 30158 26686 30210
rect 26738 30158 26750 30210
rect 22318 30146 22370 30158
rect 27246 30146 27298 30158
rect 27470 30210 27522 30222
rect 27470 30146 27522 30158
rect 28254 30210 28306 30222
rect 28254 30146 28306 30158
rect 29262 30210 29314 30222
rect 37102 30210 37154 30222
rect 40686 30210 40738 30222
rect 29586 30158 29598 30210
rect 29650 30158 29662 30210
rect 32946 30158 32958 30210
rect 33010 30158 33022 30210
rect 33506 30158 33518 30210
rect 33570 30158 33582 30210
rect 37538 30158 37550 30210
rect 37602 30158 37614 30210
rect 41234 30158 41246 30210
rect 41298 30158 41310 30210
rect 46274 30158 46286 30210
rect 46338 30158 46350 30210
rect 53890 30158 53902 30210
rect 53954 30158 53966 30210
rect 29262 30146 29314 30158
rect 37102 30146 37154 30158
rect 40686 30146 40738 30158
rect 12238 30098 12290 30110
rect 3042 30046 3054 30098
rect 3106 30046 3118 30098
rect 6066 30046 6078 30098
rect 6130 30046 6142 30098
rect 12238 30034 12290 30046
rect 16382 30098 16434 30110
rect 16382 30034 16434 30046
rect 24334 30098 24386 30110
rect 51998 30098 52050 30110
rect 46834 30046 46846 30098
rect 46898 30046 46910 30098
rect 50418 30046 50430 30098
rect 50482 30046 50494 30098
rect 51650 30046 51662 30098
rect 51714 30046 51726 30098
rect 24334 30034 24386 30046
rect 51998 30034 52050 30046
rect 52782 30098 52834 30110
rect 53106 30046 53118 30098
rect 53170 30046 53182 30098
rect 62514 30046 62526 30098
rect 62578 30046 62590 30098
rect 52782 30034 52834 30046
rect 7646 29986 7698 29998
rect 7646 29922 7698 29934
rect 8094 29986 8146 29998
rect 15598 29986 15650 29998
rect 8866 29934 8878 29986
rect 8930 29934 8942 29986
rect 8094 29922 8146 29934
rect 15598 29922 15650 29934
rect 23550 29986 23602 29998
rect 23550 29922 23602 29934
rect 27582 29986 27634 29998
rect 32734 29986 32786 29998
rect 36542 29986 36594 29998
rect 40574 29986 40626 29998
rect 44382 29986 44434 29998
rect 32162 29934 32174 29986
rect 32226 29934 32238 29986
rect 35970 29934 35982 29986
rect 36034 29934 36046 29986
rect 40002 29934 40014 29986
rect 40066 29934 40078 29986
rect 43586 29934 43598 29986
rect 43650 29934 43662 29986
rect 27582 29922 27634 29934
rect 32734 29922 32786 29934
rect 36542 29922 36594 29934
rect 40574 29922 40626 29934
rect 44382 29922 44434 29934
rect 51214 29986 51266 29998
rect 51214 29922 51266 29934
rect 1344 29818 66640 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 66640 29818
rect 1344 29732 66640 29766
rect 13246 29650 13298 29662
rect 12562 29598 12574 29650
rect 12626 29598 12638 29650
rect 13246 29586 13298 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 17950 29650 18002 29662
rect 17950 29586 18002 29598
rect 20302 29650 20354 29662
rect 20302 29586 20354 29598
rect 20862 29650 20914 29662
rect 46286 29650 46338 29662
rect 23986 29598 23998 29650
rect 24050 29598 24062 29650
rect 28130 29598 28142 29650
rect 28194 29598 28206 29650
rect 45266 29598 45278 29650
rect 45330 29598 45342 29650
rect 20862 29586 20914 29598
rect 46286 29586 46338 29598
rect 46734 29650 46786 29662
rect 46734 29586 46786 29598
rect 47182 29650 47234 29662
rect 56702 29650 56754 29662
rect 51650 29598 51662 29650
rect 51714 29598 51726 29650
rect 53106 29598 53118 29650
rect 53170 29598 53182 29650
rect 47182 29586 47234 29598
rect 56702 29586 56754 29598
rect 57150 29650 57202 29662
rect 57150 29586 57202 29598
rect 6190 29538 6242 29550
rect 3154 29486 3166 29538
rect 3218 29486 3230 29538
rect 6190 29474 6242 29486
rect 14030 29538 14082 29550
rect 29710 29538 29762 29550
rect 41246 29538 41298 29550
rect 18834 29486 18846 29538
rect 18898 29486 18910 29538
rect 33058 29486 33070 29538
rect 33122 29486 33134 29538
rect 33730 29486 33742 29538
rect 33794 29486 33806 29538
rect 40898 29486 40910 29538
rect 40962 29486 40974 29538
rect 14030 29474 14082 29486
rect 29710 29474 29762 29486
rect 41246 29474 41298 29486
rect 41918 29538 41970 29550
rect 58818 29486 58830 29538
rect 58882 29486 58894 29538
rect 61394 29486 61406 29538
rect 61458 29486 61470 29538
rect 41918 29474 41970 29486
rect 9102 29426 9154 29438
rect 8418 29374 8430 29426
rect 8482 29374 8494 29426
rect 9102 29362 9154 29374
rect 9662 29426 9714 29438
rect 21310 29426 21362 29438
rect 25342 29426 25394 29438
rect 32622 29426 32674 29438
rect 42254 29426 42306 29438
rect 48862 29426 48914 29438
rect 55918 29426 55970 29438
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 16370 29374 16382 29426
rect 16434 29374 16446 29426
rect 16818 29374 16830 29426
rect 16882 29374 16894 29426
rect 21634 29374 21646 29426
rect 21698 29374 21710 29426
rect 25778 29374 25790 29426
rect 25842 29374 25854 29426
rect 32050 29374 32062 29426
rect 32114 29374 32126 29426
rect 33954 29374 33966 29426
rect 34018 29374 34030 29426
rect 36194 29374 36206 29426
rect 36258 29374 36270 29426
rect 42914 29374 42926 29426
rect 42978 29374 42990 29426
rect 49298 29374 49310 29426
rect 49362 29374 49374 29426
rect 55570 29374 55582 29426
rect 55634 29374 55646 29426
rect 9662 29362 9714 29374
rect 21310 29362 21362 29374
rect 25342 29362 25394 29374
rect 32622 29362 32674 29374
rect 42254 29362 42306 29374
rect 48862 29362 48914 29374
rect 55918 29362 55970 29374
rect 33406 29314 33458 29326
rect 48190 29314 48242 29326
rect 4162 29262 4174 29314
rect 4226 29262 4238 29314
rect 19842 29262 19854 29314
rect 19906 29262 19918 29314
rect 38546 29262 38558 29314
rect 38610 29262 38622 29314
rect 41570 29262 41582 29314
rect 41634 29262 41646 29314
rect 47954 29262 47966 29314
rect 48018 29262 48030 29314
rect 57586 29262 57598 29314
rect 57650 29262 57662 29314
rect 60386 29262 60398 29314
rect 60450 29262 60462 29314
rect 33406 29250 33458 29262
rect 48190 29250 48242 29262
rect 5406 29202 5458 29214
rect 5406 29138 5458 29150
rect 13134 29202 13186 29214
rect 13134 29138 13186 29150
rect 24782 29202 24834 29214
rect 24782 29138 24834 29150
rect 28814 29202 28866 29214
rect 28814 29138 28866 29150
rect 28926 29202 28978 29214
rect 28926 29138 28978 29150
rect 45950 29202 46002 29214
rect 45950 29138 46002 29150
rect 52334 29202 52386 29214
rect 52334 29138 52386 29150
rect 52446 29202 52498 29214
rect 52446 29138 52498 29150
rect 1344 29034 66640 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 66640 29034
rect 1344 28948 66640 28982
rect 25790 28866 25842 28878
rect 25790 28802 25842 28814
rect 48526 28866 48578 28878
rect 48526 28802 48578 28814
rect 4510 28754 4562 28766
rect 12238 28754 12290 28766
rect 12910 28754 12962 28766
rect 16382 28754 16434 28766
rect 4050 28702 4062 28754
rect 4114 28702 4126 28754
rect 6850 28702 6862 28754
rect 6914 28702 6926 28754
rect 7858 28702 7870 28754
rect 7922 28702 7934 28754
rect 12674 28702 12686 28754
rect 12738 28702 12750 28754
rect 15698 28702 15710 28754
rect 15762 28702 15774 28754
rect 4510 28690 4562 28702
rect 12238 28690 12290 28702
rect 12910 28690 12962 28702
rect 16382 28690 16434 28702
rect 28366 28754 28418 28766
rect 28366 28690 28418 28702
rect 29262 28754 29314 28766
rect 30718 28754 30770 28766
rect 51102 28754 51154 28766
rect 51998 28754 52050 28766
rect 30482 28702 30494 28754
rect 30546 28702 30558 28754
rect 36082 28702 36094 28754
rect 36146 28702 36158 28754
rect 51650 28702 51662 28754
rect 51714 28702 51726 28754
rect 29262 28690 29314 28702
rect 30718 28690 30770 28702
rect 51102 28690 51154 28702
rect 51998 28690 52050 28702
rect 56590 28754 56642 28766
rect 57474 28702 57486 28754
rect 57538 28702 57550 28754
rect 59490 28702 59502 28754
rect 59554 28702 59566 28754
rect 61506 28702 61518 28754
rect 61570 28702 61582 28754
rect 56590 28690 56642 28702
rect 6526 28642 6578 28654
rect 6526 28578 6578 28590
rect 7198 28642 7250 28654
rect 11566 28642 11618 28654
rect 17166 28642 17218 28654
rect 22318 28642 22370 28654
rect 34638 28642 34690 28654
rect 36878 28642 36930 28654
rect 40574 28642 40626 28654
rect 44158 28642 44210 28654
rect 7634 28590 7646 28642
rect 7698 28590 7710 28642
rect 11106 28590 11118 28642
rect 11170 28590 11182 28642
rect 13794 28590 13806 28642
rect 13858 28590 13870 28642
rect 17714 28590 17726 28642
rect 17778 28590 17790 28642
rect 21522 28590 21534 28642
rect 21586 28590 21598 28642
rect 22642 28590 22654 28642
rect 22706 28590 22718 28642
rect 26002 28590 26014 28642
rect 26066 28590 26078 28642
rect 29698 28590 29710 28642
rect 29762 28590 29774 28642
rect 29922 28590 29934 28642
rect 29986 28590 29998 28642
rect 34066 28590 34078 28642
rect 34130 28590 34142 28642
rect 35074 28590 35086 28642
rect 35138 28590 35150 28642
rect 36306 28590 36318 28642
rect 36370 28590 36382 28642
rect 40002 28590 40014 28642
rect 40066 28590 40078 28642
rect 43698 28590 43710 28642
rect 43762 28590 43774 28642
rect 7198 28578 7250 28590
rect 11566 28578 11618 28590
rect 17166 28578 17218 28590
rect 22318 28578 22370 28590
rect 34638 28578 34690 28590
rect 36878 28578 36930 28590
rect 40574 28578 40626 28590
rect 44158 28578 44210 28590
rect 44830 28642 44882 28654
rect 59278 28642 59330 28654
rect 45490 28590 45502 28642
rect 45554 28590 45566 28642
rect 48738 28590 48750 28642
rect 48802 28590 48814 28642
rect 52658 28590 52670 28642
rect 52722 28590 52734 28642
rect 53218 28590 53230 28642
rect 53282 28590 53294 28642
rect 44830 28578 44882 28590
rect 59278 28578 59330 28590
rect 8878 28530 8930 28542
rect 41470 28530 41522 28542
rect 3042 28478 3054 28530
rect 3106 28478 3118 28530
rect 34850 28478 34862 28530
rect 34914 28478 34926 28530
rect 58482 28478 58494 28530
rect 58546 28478 58558 28530
rect 62514 28478 62526 28530
rect 62578 28478 62590 28530
rect 8878 28466 8930 28478
rect 41470 28466 41522 28478
rect 6414 28418 6466 28430
rect 6414 28354 6466 28366
rect 8094 28418 8146 28430
rect 8094 28354 8146 28366
rect 16494 28418 16546 28430
rect 20862 28418 20914 28430
rect 30942 28418 30994 28430
rect 40686 28418 40738 28430
rect 56254 28418 56306 28430
rect 20290 28366 20302 28418
rect 20354 28366 20366 28418
rect 21298 28366 21310 28418
rect 21362 28366 21374 28418
rect 25106 28366 25118 28418
rect 25170 28366 25182 28418
rect 31714 28366 31726 28418
rect 31778 28366 31790 28418
rect 37650 28366 37662 28418
rect 37714 28366 37726 28418
rect 47842 28366 47854 28418
rect 47906 28366 47918 28418
rect 55570 28366 55582 28418
rect 55634 28366 55646 28418
rect 16494 28354 16546 28366
rect 20862 28354 20914 28366
rect 30942 28354 30994 28366
rect 40686 28354 40738 28366
rect 56254 28354 56306 28366
rect 1344 28250 66640 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 66640 28250
rect 1344 28164 66640 28198
rect 16830 28082 16882 28094
rect 19294 28082 19346 28094
rect 26238 28082 26290 28094
rect 4722 28030 4734 28082
rect 4786 28030 4798 28082
rect 17938 28030 17950 28082
rect 18002 28030 18014 28082
rect 20738 28030 20750 28082
rect 20802 28030 20814 28082
rect 16830 28018 16882 28030
rect 19294 28018 19346 28030
rect 26238 28018 26290 28030
rect 26686 28082 26738 28094
rect 26686 28018 26738 28030
rect 27246 28082 27298 28094
rect 33182 28082 33234 28094
rect 38894 28082 38946 28094
rect 28242 28030 28254 28082
rect 28306 28030 28318 28082
rect 37314 28030 37326 28082
rect 37378 28030 37390 28082
rect 27246 28018 27298 28030
rect 33182 28018 33234 28030
rect 38894 28018 38946 28030
rect 39454 28082 39506 28094
rect 48862 28082 48914 28094
rect 56702 28082 56754 28094
rect 41570 28030 41582 28082
rect 41634 28030 41646 28082
rect 47730 28030 47742 28082
rect 47794 28030 47806 28082
rect 53106 28030 53118 28082
rect 53170 28030 53182 28082
rect 39454 28018 39506 28030
rect 48862 28018 48914 28030
rect 56702 28018 56754 28030
rect 8318 27970 8370 27982
rect 12686 27970 12738 27982
rect 10546 27918 10558 27970
rect 10610 27918 10622 27970
rect 8318 27906 8370 27918
rect 12686 27906 12738 27918
rect 24222 27970 24274 27982
rect 24222 27906 24274 27918
rect 31502 27970 31554 27982
rect 40238 27970 40290 27982
rect 55246 27970 55298 27982
rect 56030 27970 56082 27982
rect 33618 27918 33630 27970
rect 33682 27918 33694 27970
rect 38098 27918 38110 27970
rect 38162 27918 38174 27970
rect 39890 27918 39902 27970
rect 39954 27918 39966 27970
rect 54562 27918 54574 27970
rect 54626 27918 54638 27970
rect 54898 27918 54910 27970
rect 54962 27918 54974 27970
rect 55682 27918 55694 27970
rect 55746 27918 55758 27970
rect 58930 27918 58942 27970
rect 58994 27918 59006 27970
rect 61394 27918 61406 27970
rect 61458 27918 61470 27970
rect 31502 27906 31554 27918
rect 40238 27906 40290 27918
rect 55246 27906 55298 27918
rect 56030 27906 56082 27918
rect 1822 27858 1874 27870
rect 5406 27858 5458 27870
rect 9886 27858 9938 27870
rect 2258 27806 2270 27858
rect 2322 27806 2334 27858
rect 5954 27806 5966 27858
rect 6018 27806 6030 27858
rect 1822 27794 1874 27806
rect 5406 27794 5458 27806
rect 9886 27794 9938 27806
rect 10894 27858 10946 27870
rect 15598 27858 15650 27870
rect 23662 27858 23714 27870
rect 31166 27858 31218 27870
rect 34414 27858 34466 27870
rect 44270 27858 44322 27870
rect 11442 27806 11454 27858
rect 11506 27806 11518 27858
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 18162 27806 18174 27858
rect 18226 27806 18238 27858
rect 22978 27806 22990 27858
rect 23042 27806 23054 27858
rect 25218 27806 25230 27858
rect 25282 27806 25294 27858
rect 30594 27806 30606 27858
rect 30658 27806 30670 27858
rect 32386 27806 32398 27858
rect 32450 27806 32462 27858
rect 33842 27806 33854 27858
rect 33906 27806 33918 27858
rect 34738 27806 34750 27858
rect 34802 27806 34814 27858
rect 38322 27806 38334 27858
rect 38386 27806 38398 27858
rect 43922 27806 43934 27858
rect 43986 27806 43998 27858
rect 10894 27794 10946 27806
rect 15598 27794 15650 27806
rect 23662 27794 23714 27806
rect 31166 27794 31218 27806
rect 34414 27794 34466 27806
rect 44270 27794 44322 27806
rect 44830 27858 44882 27870
rect 49982 27858 50034 27870
rect 45266 27806 45278 27858
rect 45330 27806 45342 27858
rect 50642 27806 50654 27858
rect 50706 27806 50718 27858
rect 54338 27806 54350 27858
rect 54402 27806 54414 27858
rect 44830 27794 44882 27806
rect 49982 27794 50034 27806
rect 15934 27746 15986 27758
rect 9538 27694 9550 27746
rect 9602 27694 9614 27746
rect 11666 27694 11678 27746
rect 11730 27694 11742 27746
rect 15934 27682 15986 27694
rect 16382 27746 16434 27758
rect 16382 27682 16434 27694
rect 17614 27746 17666 27758
rect 17614 27682 17666 27694
rect 19742 27746 19794 27758
rect 24670 27746 24722 27758
rect 39566 27746 39618 27758
rect 49534 27746 49586 27758
rect 23874 27694 23886 27746
rect 23938 27694 23950 27746
rect 31826 27694 31838 27746
rect 31890 27694 31902 27746
rect 32162 27694 32174 27746
rect 32226 27694 32238 27746
rect 49186 27694 49198 27746
rect 49250 27694 49262 27746
rect 57586 27694 57598 27746
rect 57650 27694 57662 27746
rect 60386 27694 60398 27746
rect 60450 27694 60462 27746
rect 19742 27682 19794 27694
rect 24670 27682 24722 27694
rect 39566 27682 39618 27694
rect 49534 27682 49586 27694
rect 5294 27634 5346 27646
rect 5294 27570 5346 27582
rect 9102 27634 9154 27646
rect 9102 27570 9154 27582
rect 11902 27634 11954 27646
rect 19966 27634 20018 27646
rect 27470 27634 27522 27646
rect 15922 27582 15934 27634
rect 15986 27631 15998 27634
rect 16706 27631 16718 27634
rect 15986 27585 16718 27631
rect 15986 27582 15998 27585
rect 16706 27582 16718 27585
rect 16770 27582 16782 27634
rect 25778 27582 25790 27634
rect 25842 27582 25854 27634
rect 26226 27582 26238 27634
rect 26290 27631 26302 27634
rect 27010 27631 27022 27634
rect 26290 27585 27022 27631
rect 26290 27582 26302 27585
rect 27010 27582 27022 27585
rect 27074 27582 27086 27634
rect 11902 27570 11954 27582
rect 19966 27570 20018 27582
rect 27470 27570 27522 27582
rect 37886 27634 37938 27646
rect 37886 27570 37938 27582
rect 40798 27634 40850 27646
rect 40798 27570 40850 27582
rect 48302 27634 48354 27646
rect 48302 27570 48354 27582
rect 53678 27634 53730 27646
rect 53678 27570 53730 27582
rect 1344 27466 66640 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 66640 27466
rect 1344 27380 66640 27414
rect 56254 27298 56306 27310
rect 21298 27246 21310 27298
rect 21362 27246 21374 27298
rect 56254 27234 56306 27246
rect 12798 27186 12850 27198
rect 15374 27186 15426 27198
rect 3938 27134 3950 27186
rect 4002 27134 4014 27186
rect 13682 27134 13694 27186
rect 13746 27134 13758 27186
rect 12798 27122 12850 27134
rect 15374 27122 15426 27134
rect 27022 27186 27074 27198
rect 28590 27186 28642 27198
rect 35758 27186 35810 27198
rect 51886 27186 51938 27198
rect 28242 27134 28254 27186
rect 28306 27134 28318 27186
rect 33954 27134 33966 27186
rect 34018 27134 34030 27186
rect 49746 27134 49758 27186
rect 49810 27134 49822 27186
rect 51538 27134 51550 27186
rect 51602 27134 51614 27186
rect 57474 27134 57486 27186
rect 57538 27134 57550 27186
rect 59266 27134 59278 27186
rect 59330 27134 59342 27186
rect 61506 27134 61518 27186
rect 61570 27134 61582 27186
rect 27022 27122 27074 27134
rect 28590 27122 28642 27134
rect 35758 27122 35810 27134
rect 51886 27122 51938 27134
rect 17390 27074 17442 27086
rect 23214 27074 23266 27086
rect 29262 27074 29314 27086
rect 37102 27074 37154 27086
rect 40686 27074 40738 27086
rect 44718 27074 44770 27086
rect 52782 27074 52834 27086
rect 11666 27022 11678 27074
rect 11730 27022 11742 27074
rect 13906 27022 13918 27074
rect 13970 27022 13982 27074
rect 14802 27022 14814 27074
rect 14866 27022 14878 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 21522 27022 21534 27074
rect 21586 27022 21598 27074
rect 22418 27022 22430 27074
rect 22482 27022 22494 27074
rect 23650 27022 23662 27074
rect 23714 27022 23726 27074
rect 29698 27022 29710 27074
rect 29762 27022 29774 27074
rect 37538 27022 37550 27074
rect 37602 27022 37614 27074
rect 41346 27022 41358 27074
rect 41410 27022 41422 27074
rect 45378 27022 45390 27074
rect 45442 27022 45454 27074
rect 50754 27022 50766 27074
rect 50818 27022 50830 27074
rect 53218 27022 53230 27074
rect 53282 27022 53294 27074
rect 59490 27022 59502 27074
rect 59554 27022 59566 27074
rect 17390 27010 17442 27022
rect 23214 27010 23266 27022
rect 29262 27010 29314 27022
rect 37102 27010 37154 27022
rect 40686 27010 40738 27022
rect 44718 27010 44770 27022
rect 52782 27010 52834 27022
rect 5742 26962 5794 26974
rect 20078 26962 20130 26974
rect 3042 26910 3054 26962
rect 3106 26910 3118 26962
rect 7186 26910 7198 26962
rect 7250 26910 7262 26962
rect 5742 26898 5794 26910
rect 20078 26898 20130 26910
rect 25902 26962 25954 26974
rect 25902 26898 25954 26910
rect 27470 26962 27522 26974
rect 27470 26898 27522 26910
rect 27918 26962 27970 26974
rect 27918 26898 27970 26910
rect 31950 26962 32002 26974
rect 39790 26962 39842 26974
rect 34962 26910 34974 26962
rect 35026 26910 35038 26962
rect 36082 26910 36094 26962
rect 36146 26910 36158 26962
rect 58482 26910 58494 26962
rect 58546 26910 58558 26962
rect 62514 26910 62526 26962
rect 62578 26910 62590 26962
rect 31950 26898 32002 26910
rect 39790 26898 39842 26910
rect 20862 26850 20914 26862
rect 26686 26850 26738 26862
rect 22194 26798 22206 26850
rect 22258 26798 22270 26850
rect 20862 26786 20914 26798
rect 26686 26786 26738 26798
rect 32734 26850 32786 26862
rect 32734 26786 32786 26798
rect 40574 26850 40626 26862
rect 44382 26850 44434 26862
rect 48414 26850 48466 26862
rect 43810 26798 43822 26850
rect 43874 26798 43886 26850
rect 47842 26798 47854 26850
rect 47906 26798 47918 26850
rect 55458 26798 55470 26850
rect 55522 26798 55534 26850
rect 40574 26786 40626 26798
rect 44382 26786 44434 26798
rect 48414 26786 48466 26798
rect 1344 26682 66640 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 66640 26682
rect 1344 26596 66640 26630
rect 41022 26514 41074 26526
rect 45054 26514 45106 26526
rect 52782 26514 52834 26526
rect 7410 26462 7422 26514
rect 7474 26462 7486 26514
rect 15026 26462 15038 26514
rect 15090 26462 15102 26514
rect 28242 26462 28254 26514
rect 28306 26462 28318 26514
rect 32050 26462 32062 26514
rect 32114 26462 32126 26514
rect 33730 26462 33742 26514
rect 33794 26462 33806 26514
rect 44482 26462 44494 26514
rect 44546 26462 44558 26514
rect 51762 26462 51774 26514
rect 51826 26462 51838 26514
rect 41022 26450 41074 26462
rect 45054 26450 45106 26462
rect 52782 26450 52834 26462
rect 53118 26514 53170 26526
rect 53118 26450 53170 26462
rect 55470 26514 55522 26526
rect 55470 26450 55522 26462
rect 8766 26402 8818 26414
rect 2034 26350 2046 26402
rect 2098 26350 2110 26402
rect 8418 26350 8430 26402
rect 8482 26350 8494 26402
rect 8766 26338 8818 26350
rect 18062 26402 18114 26414
rect 18062 26338 18114 26350
rect 23998 26402 24050 26414
rect 23998 26338 24050 26350
rect 39678 26402 39730 26414
rect 54562 26350 54574 26402
rect 54626 26350 54638 26402
rect 58818 26350 58830 26402
rect 58882 26350 58894 26402
rect 61394 26350 61406 26402
rect 61458 26350 61470 26402
rect 39678 26338 39730 26350
rect 4510 26290 4562 26302
rect 12126 26290 12178 26302
rect 21086 26290 21138 26302
rect 25118 26290 25170 26302
rect 29150 26290 29202 26302
rect 36430 26290 36482 26302
rect 5058 26238 5070 26290
rect 5122 26238 5134 26290
rect 9762 26238 9774 26290
rect 9826 26238 9838 26290
rect 10882 26238 10894 26290
rect 10946 26238 10958 26290
rect 12674 26238 12686 26290
rect 12738 26238 12750 26290
rect 20402 26238 20414 26290
rect 20466 26238 20478 26290
rect 20850 26238 20862 26290
rect 20914 26238 20926 26290
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 25666 26238 25678 26290
rect 25730 26238 25742 26290
rect 29586 26238 29598 26290
rect 29650 26238 29662 26290
rect 36082 26238 36094 26290
rect 36146 26238 36158 26290
rect 4510 26226 4562 26238
rect 12126 26226 12178 26238
rect 21086 26226 21138 26238
rect 25118 26226 25170 26238
rect 29150 26226 29202 26238
rect 36430 26226 36482 26238
rect 36766 26290 36818 26302
rect 41358 26290 41410 26302
rect 48862 26290 48914 26302
rect 37426 26238 37438 26290
rect 37490 26238 37502 26290
rect 42018 26238 42030 26290
rect 42082 26238 42094 26290
rect 45378 26238 45390 26290
rect 45442 26238 45454 26290
rect 49298 26238 49310 26290
rect 49362 26238 49374 26290
rect 36766 26226 36818 26238
rect 41358 26226 41410 26238
rect 48862 26226 48914 26238
rect 10334 26178 10386 26190
rect 11454 26178 11506 26190
rect 3266 26126 3278 26178
rect 3330 26126 3342 26178
rect 9538 26126 9550 26178
rect 9602 26126 9614 26178
rect 10658 26126 10670 26178
rect 10722 26126 10734 26178
rect 10334 26114 10386 26126
rect 11454 26114 11506 26126
rect 11902 26178 11954 26190
rect 11902 26114 11954 26126
rect 16382 26178 16434 26190
rect 16382 26114 16434 26126
rect 16830 26178 16882 26190
rect 55358 26178 55410 26190
rect 46946 26126 46958 26178
rect 47010 26126 47022 26178
rect 53554 26126 53566 26178
rect 53618 26126 53630 26178
rect 57586 26126 57598 26178
rect 57650 26126 57662 26178
rect 60386 26126 60398 26178
rect 60450 26126 60462 26178
rect 16830 26114 16882 26126
rect 55358 26114 55410 26126
rect 8206 26066 8258 26078
rect 8206 26002 8258 26014
rect 15822 26066 15874 26078
rect 15822 26002 15874 26014
rect 17278 26066 17330 26078
rect 17278 26002 17330 26014
rect 24782 26066 24834 26078
rect 24782 26002 24834 26014
rect 28814 26066 28866 26078
rect 28814 26002 28866 26014
rect 32622 26066 32674 26078
rect 32622 26002 32674 26014
rect 32958 26066 33010 26078
rect 32958 26002 33010 26014
rect 40462 26066 40514 26078
rect 40462 26002 40514 26014
rect 52334 26066 52386 26078
rect 52334 26002 52386 26014
rect 1344 25898 66640 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 66640 25898
rect 1344 25812 66640 25846
rect 19394 25678 19406 25730
rect 19458 25678 19470 25730
rect 5966 25618 6018 25630
rect 8318 25618 8370 25630
rect 4050 25566 4062 25618
rect 4114 25566 4126 25618
rect 7746 25566 7758 25618
rect 7810 25566 7822 25618
rect 5966 25554 6018 25566
rect 8318 25554 8370 25566
rect 8766 25618 8818 25630
rect 8766 25554 8818 25566
rect 13582 25618 13634 25630
rect 13582 25554 13634 25566
rect 14702 25618 14754 25630
rect 24110 25618 24162 25630
rect 21746 25566 21758 25618
rect 21810 25566 21822 25618
rect 23538 25566 23550 25618
rect 23602 25566 23614 25618
rect 14702 25554 14754 25566
rect 24110 25554 24162 25566
rect 29486 25618 29538 25630
rect 29486 25554 29538 25566
rect 30494 25618 30546 25630
rect 30494 25554 30546 25566
rect 42702 25618 42754 25630
rect 44046 25618 44098 25630
rect 43362 25566 43374 25618
rect 43426 25566 43438 25618
rect 43810 25566 43822 25618
rect 43874 25566 43886 25618
rect 42702 25554 42754 25566
rect 44046 25554 44098 25566
rect 44942 25618 44994 25630
rect 44942 25554 44994 25566
rect 51550 25618 51602 25630
rect 59502 25618 59554 25630
rect 57698 25566 57710 25618
rect 57762 25566 57774 25618
rect 51550 25554 51602 25566
rect 59502 25554 59554 25566
rect 8990 25506 9042 25518
rect 15710 25506 15762 25518
rect 24782 25506 24834 25518
rect 31390 25506 31442 25518
rect 38446 25506 38498 25518
rect 45278 25506 45330 25518
rect 48974 25506 49026 25518
rect 9538 25454 9550 25506
rect 9602 25454 9614 25506
rect 16146 25454 16158 25506
rect 16210 25454 16222 25506
rect 19618 25454 19630 25506
rect 19682 25454 19694 25506
rect 20626 25454 20638 25506
rect 20690 25454 20702 25506
rect 25330 25454 25342 25506
rect 25394 25454 25406 25506
rect 32050 25454 32062 25506
rect 32114 25454 32126 25506
rect 38098 25454 38110 25506
rect 38162 25454 38174 25506
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 43138 25454 43150 25506
rect 43202 25454 43214 25506
rect 45938 25454 45950 25506
rect 46002 25454 46014 25506
rect 49186 25454 49198 25506
rect 49250 25454 49262 25506
rect 52882 25454 52894 25506
rect 52946 25454 52958 25506
rect 53442 25454 53454 25506
rect 53506 25454 53518 25506
rect 8990 25442 9042 25454
rect 15710 25442 15762 25454
rect 24782 25442 24834 25454
rect 31390 25442 31442 25454
rect 38446 25442 38498 25454
rect 45278 25442 45330 25454
rect 48974 25442 49026 25454
rect 1710 25394 1762 25406
rect 15262 25394 15314 25406
rect 2930 25342 2942 25394
rect 2994 25342 3006 25394
rect 6626 25342 6638 25394
rect 6690 25342 6702 25394
rect 14914 25342 14926 25394
rect 14978 25342 14990 25394
rect 1710 25330 1762 25342
rect 15262 25330 15314 25342
rect 19182 25394 19234 25406
rect 19182 25330 19234 25342
rect 21422 25394 21474 25406
rect 48190 25394 48242 25406
rect 22530 25342 22542 25394
rect 22594 25342 22606 25394
rect 37874 25342 37886 25394
rect 37938 25342 37950 25394
rect 42354 25342 42366 25394
rect 42418 25342 42430 25394
rect 58818 25342 58830 25394
rect 58882 25342 58894 25394
rect 21422 25330 21474 25342
rect 48190 25330 48242 25342
rect 2046 25282 2098 25294
rect 2046 25218 2098 25230
rect 5854 25282 5906 25294
rect 12686 25282 12738 25294
rect 20638 25282 20690 25294
rect 12002 25230 12014 25282
rect 12066 25230 12078 25282
rect 18386 25230 18398 25282
rect 18450 25230 18462 25282
rect 5854 25218 5906 25230
rect 12686 25218 12738 25230
rect 20638 25218 20690 25230
rect 24558 25282 24610 25294
rect 28478 25282 28530 25294
rect 27906 25230 27918 25282
rect 27970 25230 27982 25282
rect 24558 25218 24610 25230
rect 28478 25218 28530 25230
rect 29374 25282 29426 25294
rect 29374 25218 29426 25230
rect 30382 25282 30434 25294
rect 30382 25218 30434 25230
rect 30942 25282 30994 25294
rect 35086 25282 35138 25294
rect 42142 25282 42194 25294
rect 56478 25282 56530 25294
rect 34514 25230 34526 25282
rect 34578 25230 34590 25282
rect 41570 25230 41582 25282
rect 41634 25230 41646 25282
rect 55906 25230 55918 25282
rect 55970 25230 55982 25282
rect 30942 25218 30994 25230
rect 35086 25218 35138 25230
rect 42142 25218 42194 25230
rect 56478 25218 56530 25230
rect 59614 25282 59666 25294
rect 59614 25218 59666 25230
rect 1344 25114 66640 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 66640 25114
rect 1344 25028 66640 25062
rect 19182 24946 19234 24958
rect 39678 24946 39730 24958
rect 50206 24946 50258 24958
rect 4722 24894 4734 24946
rect 4786 24894 4798 24946
rect 8306 24894 8318 24946
rect 8370 24894 8382 24946
rect 16370 24894 16382 24946
rect 16434 24894 16446 24946
rect 20626 24894 20638 24946
rect 20690 24894 20702 24946
rect 43922 24894 43934 24946
rect 43986 24894 43998 24946
rect 47730 24894 47742 24946
rect 47794 24894 47806 24946
rect 54338 24894 54350 24946
rect 54402 24894 54414 24946
rect 19182 24882 19234 24894
rect 39678 24882 39730 24894
rect 50206 24882 50258 24894
rect 12350 24834 12402 24846
rect 12350 24770 12402 24782
rect 19630 24834 19682 24846
rect 39566 24834 39618 24846
rect 30034 24782 30046 24834
rect 30098 24782 30110 24834
rect 34066 24782 34078 24834
rect 34130 24782 34142 24834
rect 19630 24770 19682 24782
rect 39566 24770 39618 24782
rect 48750 24834 48802 24846
rect 49758 24834 49810 24846
rect 49074 24782 49086 24834
rect 49138 24782 49150 24834
rect 48750 24770 48802 24782
rect 49758 24770 49810 24782
rect 50094 24834 50146 24846
rect 50094 24770 50146 24782
rect 50878 24834 50930 24846
rect 55122 24782 55134 24834
rect 55186 24782 55198 24834
rect 58818 24782 58830 24834
rect 58882 24782 58894 24834
rect 61394 24782 61406 24834
rect 61458 24782 61470 24834
rect 50878 24770 50930 24782
rect 1822 24722 1874 24734
rect 5406 24722 5458 24734
rect 9438 24722 9490 24734
rect 17614 24722 17666 24734
rect 23326 24722 23378 24734
rect 30942 24722 30994 24734
rect 41022 24722 41074 24734
rect 44830 24722 44882 24734
rect 51214 24722 51266 24734
rect 2146 24670 2158 24722
rect 2210 24670 2222 24722
rect 5954 24670 5966 24722
rect 6018 24670 6030 24722
rect 10098 24670 10110 24722
rect 10162 24670 10174 24722
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 13794 24670 13806 24722
rect 13858 24670 13870 24722
rect 17938 24670 17950 24722
rect 18002 24670 18014 24722
rect 22866 24670 22878 24722
rect 22930 24670 22942 24722
rect 24658 24670 24670 24722
rect 24722 24670 24734 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 39106 24670 39118 24722
rect 39170 24670 39182 24722
rect 41346 24670 41358 24722
rect 41410 24670 41422 24722
rect 45266 24670 45278 24722
rect 45330 24670 45342 24722
rect 51874 24670 51886 24722
rect 51938 24670 51950 24722
rect 1822 24658 1874 24670
rect 5406 24658 5458 24670
rect 9438 24658 9490 24670
rect 17614 24658 17666 24670
rect 23326 24658 23378 24670
rect 30942 24658 30994 24670
rect 41022 24658 41074 24670
rect 44830 24658 44882 24670
rect 51214 24658 51266 24670
rect 40350 24610 40402 24622
rect 55470 24610 55522 24622
rect 18386 24558 18398 24610
rect 18450 24558 18462 24610
rect 49410 24558 49422 24610
rect 49474 24558 49486 24610
rect 57586 24558 57598 24610
rect 57650 24558 57662 24610
rect 60386 24558 60398 24610
rect 60450 24558 60462 24610
rect 40350 24546 40402 24558
rect 55470 24546 55522 24558
rect 5294 24498 5346 24510
rect 5294 24434 5346 24446
rect 9102 24498 9154 24510
rect 9102 24434 9154 24446
rect 13134 24498 13186 24510
rect 13134 24434 13186 24446
rect 16942 24498 16994 24510
rect 16942 24434 16994 24446
rect 19854 24498 19906 24510
rect 44494 24498 44546 24510
rect 24098 24446 24110 24498
rect 24162 24446 24174 24498
rect 19854 24434 19906 24446
rect 44494 24434 44546 24446
rect 48302 24498 48354 24510
rect 48302 24434 48354 24446
rect 54910 24498 54962 24510
rect 54910 24434 54962 24446
rect 1344 24330 66640 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 66640 24330
rect 1344 24244 66640 24278
rect 1822 24050 1874 24062
rect 5070 24050 5122 24062
rect 3826 23998 3838 24050
rect 3890 23998 3902 24050
rect 1822 23986 1874 23998
rect 5070 23986 5122 23998
rect 5854 24050 5906 24062
rect 6526 24050 6578 24062
rect 6178 23998 6190 24050
rect 6242 23998 6254 24050
rect 5854 23986 5906 23998
rect 6526 23986 6578 23998
rect 11454 24050 11506 24062
rect 19966 24050 20018 24062
rect 12226 23998 12238 24050
rect 12290 23998 12302 24050
rect 19058 23998 19070 24050
rect 19122 23998 19134 24050
rect 11454 23986 11506 23998
rect 19966 23986 20018 23998
rect 20302 24050 20354 24062
rect 20302 23986 20354 23998
rect 20750 24050 20802 24062
rect 29486 24050 29538 24062
rect 29138 23998 29150 24050
rect 29202 23998 29214 24050
rect 20750 23986 20802 23998
rect 29486 23986 29538 23998
rect 45054 24050 45106 24062
rect 45054 23986 45106 23998
rect 49310 24050 49362 24062
rect 49310 23986 49362 23998
rect 49646 24050 49698 24062
rect 51998 24050 52050 24062
rect 58606 24050 58658 24062
rect 50082 23998 50094 24050
rect 50146 23998 50158 24050
rect 52882 23998 52894 24050
rect 52946 23998 52958 24050
rect 49646 23986 49698 23998
rect 51998 23986 52050 23998
rect 58606 23986 58658 23998
rect 10222 23938 10274 23950
rect 11902 23938 11954 23950
rect 9762 23886 9774 23938
rect 9826 23886 9838 23938
rect 10882 23886 10894 23938
rect 10946 23886 10958 23938
rect 10222 23874 10274 23886
rect 11902 23874 11954 23886
rect 12910 23938 12962 23950
rect 21198 23938 21250 23950
rect 25006 23938 25058 23950
rect 35086 23938 35138 23950
rect 37102 23938 37154 23950
rect 40686 23938 40738 23950
rect 17266 23886 17278 23938
rect 17330 23886 17342 23938
rect 19282 23886 19294 23938
rect 19346 23886 19358 23938
rect 21746 23886 21758 23938
rect 21810 23886 21822 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 34626 23886 34638 23938
rect 34690 23886 34702 23938
rect 35746 23886 35758 23938
rect 35810 23886 35822 23938
rect 37426 23886 37438 23938
rect 37490 23886 37502 23938
rect 41234 23886 41246 23938
rect 41298 23886 41310 23938
rect 45266 23886 45278 23938
rect 45330 23886 45342 23938
rect 45826 23886 45838 23938
rect 45890 23886 45902 23938
rect 56466 23886 56478 23938
rect 56530 23886 56542 23938
rect 12910 23874 12962 23886
rect 21198 23874 21250 23886
rect 25006 23874 25058 23886
rect 35086 23874 35138 23886
rect 37102 23874 37154 23886
rect 40686 23874 40738 23886
rect 6750 23826 6802 23838
rect 3042 23774 3054 23826
rect 3106 23774 3118 23826
rect 6750 23762 6802 23774
rect 7534 23826 7586 23838
rect 24110 23826 24162 23838
rect 10658 23774 10670 23826
rect 10722 23774 10734 23826
rect 12562 23774 12574 23826
rect 12626 23774 12638 23826
rect 13682 23774 13694 23826
rect 13746 23774 13758 23826
rect 7534 23762 7586 23774
rect 24110 23762 24162 23774
rect 30606 23826 30658 23838
rect 35522 23774 35534 23826
rect 35586 23774 35598 23826
rect 51090 23774 51102 23826
rect 51154 23774 51166 23826
rect 58258 23774 58270 23826
rect 58322 23774 58334 23826
rect 30606 23762 30658 23774
rect 24894 23714 24946 23726
rect 28702 23714 28754 23726
rect 28130 23662 28142 23714
rect 28194 23662 28206 23714
rect 24894 23650 24946 23662
rect 28702 23650 28754 23662
rect 29934 23714 29986 23726
rect 29934 23650 29986 23662
rect 30718 23714 30770 23726
rect 30718 23650 30770 23662
rect 31614 23714 31666 23726
rect 40574 23714 40626 23726
rect 44382 23714 44434 23726
rect 48862 23714 48914 23726
rect 32386 23662 32398 23714
rect 32450 23662 32462 23714
rect 39778 23662 39790 23714
rect 39842 23662 39854 23714
rect 43810 23662 43822 23714
rect 43874 23662 43886 23714
rect 48066 23662 48078 23714
rect 48130 23662 48142 23714
rect 31614 23650 31666 23662
rect 40574 23650 40626 23662
rect 44382 23650 44434 23662
rect 48862 23650 48914 23662
rect 1344 23546 66640 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 66640 23546
rect 1344 23460 66640 23494
rect 40350 23378 40402 23390
rect 8306 23326 8318 23378
rect 8370 23326 8382 23378
rect 10210 23326 10222 23378
rect 10274 23326 10286 23378
rect 14018 23326 14030 23378
rect 14082 23326 14094 23378
rect 21858 23326 21870 23378
rect 21922 23326 21934 23378
rect 28242 23326 28254 23378
rect 28306 23326 28318 23378
rect 32050 23326 32062 23378
rect 32114 23326 32126 23378
rect 37426 23326 37438 23378
rect 37490 23326 37502 23378
rect 40350 23314 40402 23326
rect 47854 23378 47906 23390
rect 51650 23326 51662 23378
rect 51714 23326 51726 23378
rect 47854 23314 47906 23326
rect 18062 23266 18114 23278
rect 47966 23266 48018 23278
rect 2818 23214 2830 23266
rect 2882 23214 2894 23266
rect 33058 23214 33070 23266
rect 33122 23214 33134 23266
rect 33730 23214 33742 23266
rect 33794 23214 33806 23266
rect 39218 23214 39230 23266
rect 39282 23214 39294 23266
rect 18062 23202 18114 23214
rect 47966 23202 48018 23214
rect 55358 23266 55410 23278
rect 58818 23214 58830 23266
rect 58882 23214 58894 23266
rect 55358 23202 55410 23214
rect 5406 23154 5458 23166
rect 12910 23154 12962 23166
rect 20750 23154 20802 23166
rect 24782 23154 24834 23166
rect 5954 23102 5966 23154
rect 6018 23102 6030 23154
rect 12562 23102 12574 23154
rect 12626 23102 12638 23154
rect 16258 23102 16270 23154
rect 16322 23102 16334 23154
rect 16818 23102 16830 23154
rect 16882 23102 16894 23154
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 5406 23090 5458 23102
rect 12910 23090 12962 23102
rect 20750 23090 20802 23102
rect 24782 23090 24834 23102
rect 25118 23154 25170 23166
rect 29150 23154 29202 23166
rect 34302 23154 34354 23166
rect 38894 23154 38946 23166
rect 25666 23102 25678 23154
rect 25730 23102 25742 23154
rect 29586 23102 29598 23154
rect 29650 23102 29662 23154
rect 33282 23102 33294 23154
rect 33346 23102 33358 23154
rect 33954 23102 33966 23154
rect 34018 23102 34030 23154
rect 34962 23102 34974 23154
rect 35026 23102 35038 23154
rect 38434 23102 38446 23154
rect 38498 23102 38510 23154
rect 25118 23090 25170 23102
rect 29150 23090 29202 23102
rect 34302 23090 34354 23102
rect 38894 23090 38946 23102
rect 39566 23154 39618 23166
rect 39566 23090 39618 23102
rect 41694 23154 41746 23166
rect 48862 23154 48914 23166
rect 52446 23154 52498 23166
rect 42018 23102 42030 23154
rect 42082 23102 42094 23154
rect 49298 23102 49310 23154
rect 49362 23102 49374 23154
rect 52994 23102 53006 23154
rect 53058 23102 53070 23154
rect 59490 23102 59502 23154
rect 59554 23102 59566 23154
rect 41694 23090 41746 23102
rect 48862 23090 48914 23102
rect 52446 23090 52498 23102
rect 41022 23042 41074 23054
rect 3938 22990 3950 23042
rect 4002 22990 4014 23042
rect 38210 22990 38222 23042
rect 38274 22990 38286 23042
rect 39778 22990 39790 23042
rect 39842 22990 39854 23042
rect 46946 22990 46958 23042
rect 47010 22990 47022 23042
rect 57586 22990 57598 23042
rect 57650 22990 57662 23042
rect 59602 22990 59614 23042
rect 59666 22990 59678 23042
rect 41022 22978 41074 22990
rect 9102 22930 9154 22942
rect 9102 22866 9154 22878
rect 9438 22930 9490 22942
rect 9438 22866 9490 22878
rect 13246 22930 13298 22942
rect 13246 22866 13298 22878
rect 17278 22930 17330 22942
rect 17278 22866 17330 22878
rect 21086 22930 21138 22942
rect 21086 22866 21138 22878
rect 28814 22930 28866 22942
rect 28814 22866 28866 22878
rect 32622 22930 32674 22942
rect 32622 22866 32674 22878
rect 37998 22930 38050 22942
rect 37998 22866 38050 22878
rect 52334 22930 52386 22942
rect 52334 22866 52386 22878
rect 56142 22930 56194 22942
rect 56142 22866 56194 22878
rect 1344 22762 66640 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 66640 22762
rect 1344 22676 66640 22710
rect 56254 22594 56306 22606
rect 27010 22542 27022 22594
rect 27074 22591 27086 22594
rect 27346 22591 27358 22594
rect 27074 22545 27358 22591
rect 27074 22542 27086 22545
rect 27346 22542 27358 22545
rect 27410 22542 27422 22594
rect 56254 22530 56306 22542
rect 27022 22482 27074 22494
rect 4050 22430 4062 22482
rect 4114 22430 4126 22482
rect 27022 22418 27074 22430
rect 27470 22482 27522 22494
rect 27470 22418 27522 22430
rect 27918 22482 27970 22494
rect 28242 22430 28254 22482
rect 28306 22430 28318 22482
rect 57474 22430 57486 22482
rect 57538 22430 57550 22482
rect 27918 22418 27970 22430
rect 5518 22370 5570 22382
rect 9326 22370 9378 22382
rect 13582 22370 13634 22382
rect 17166 22370 17218 22382
rect 33070 22370 33122 22382
rect 40350 22370 40402 22382
rect 6178 22318 6190 22370
rect 6242 22318 6254 22370
rect 9986 22318 9998 22370
rect 10050 22318 10062 22370
rect 13906 22318 13918 22370
rect 13970 22318 13982 22370
rect 17826 22318 17838 22370
rect 17890 22318 17902 22370
rect 22754 22318 22766 22370
rect 22818 22318 22830 22370
rect 29138 22318 29150 22370
rect 29202 22318 29214 22370
rect 33394 22318 33406 22370
rect 33458 22318 33470 22370
rect 40002 22318 40014 22370
rect 40066 22318 40078 22370
rect 5518 22306 5570 22318
rect 9326 22306 9378 22318
rect 13582 22306 13634 22318
rect 17166 22306 17218 22318
rect 33070 22306 33122 22318
rect 40350 22306 40402 22318
rect 40910 22370 40962 22382
rect 52558 22370 52610 22382
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 44818 22318 44830 22370
rect 44882 22318 44894 22370
rect 45378 22318 45390 22370
rect 45442 22318 45454 22370
rect 48626 22318 48638 22370
rect 48690 22318 48702 22370
rect 49074 22318 49086 22370
rect 49138 22318 49150 22370
rect 53218 22318 53230 22370
rect 53282 22318 53294 22370
rect 40910 22306 40962 22318
rect 52558 22306 52610 22318
rect 28590 22258 28642 22270
rect 2706 22206 2718 22258
rect 2770 22206 2782 22258
rect 23538 22206 23550 22258
rect 23602 22206 23614 22258
rect 28590 22194 28642 22206
rect 37662 22258 37714 22270
rect 37662 22194 37714 22206
rect 48414 22258 48466 22270
rect 58482 22206 58494 22258
rect 58546 22206 58558 22258
rect 48414 22194 48466 22206
rect 9214 22146 9266 22158
rect 13022 22146 13074 22158
rect 17054 22146 17106 22158
rect 20862 22146 20914 22158
rect 8642 22094 8654 22146
rect 8706 22094 8718 22146
rect 12450 22094 12462 22146
rect 12514 22094 12526 22146
rect 16482 22094 16494 22146
rect 16546 22094 16558 22146
rect 20178 22094 20190 22146
rect 20242 22094 20254 22146
rect 9214 22082 9266 22094
rect 13022 22082 13074 22094
rect 17054 22082 17106 22094
rect 20862 22082 20914 22094
rect 30158 22146 30210 22158
rect 36542 22146 36594 22158
rect 35970 22094 35982 22146
rect 36034 22094 36046 22146
rect 30158 22082 30210 22094
rect 36542 22082 36594 22094
rect 36878 22146 36930 22158
rect 44382 22146 44434 22158
rect 52222 22146 52274 22158
rect 43586 22094 43598 22146
rect 43650 22094 43662 22146
rect 47618 22094 47630 22146
rect 47682 22094 47694 22146
rect 51426 22094 51438 22146
rect 51490 22094 51502 22146
rect 55682 22094 55694 22146
rect 55746 22094 55758 22146
rect 36878 22082 36930 22094
rect 44382 22082 44434 22094
rect 52222 22082 52274 22094
rect 1344 21978 66640 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 66640 21978
rect 1344 21892 66640 21926
rect 25342 21810 25394 21822
rect 10210 21758 10222 21810
rect 10274 21758 10286 21810
rect 20962 21758 20974 21810
rect 21026 21758 21038 21810
rect 25342 21746 25394 21758
rect 26910 21810 26962 21822
rect 45614 21810 45666 21822
rect 30706 21758 30718 21810
rect 30770 21758 30782 21810
rect 36530 21758 36542 21810
rect 36594 21758 36606 21810
rect 42354 21758 42366 21810
rect 42418 21758 42430 21810
rect 26910 21746 26962 21758
rect 45614 21746 45666 21758
rect 46062 21810 46114 21822
rect 53006 21810 53058 21822
rect 51762 21758 51774 21810
rect 51826 21758 51838 21810
rect 46062 21746 46114 21758
rect 53006 21746 53058 21758
rect 8318 21698 8370 21710
rect 3154 21646 3166 21698
rect 3218 21646 3230 21698
rect 8318 21634 8370 21646
rect 16158 21698 16210 21710
rect 55918 21698 55970 21710
rect 35186 21646 35198 21698
rect 35250 21646 35262 21698
rect 47730 21646 47742 21698
rect 47794 21646 47806 21698
rect 54786 21646 54798 21698
rect 54850 21646 54862 21698
rect 55570 21646 55582 21698
rect 55634 21646 55646 21698
rect 58818 21646 58830 21698
rect 58882 21646 58894 21698
rect 16158 21634 16210 21646
rect 55918 21634 55970 21646
rect 5630 21586 5682 21598
rect 12910 21586 12962 21598
rect 5954 21534 5966 21586
rect 6018 21534 6030 21586
rect 12450 21534 12462 21586
rect 12514 21534 12526 21586
rect 5630 21522 5682 21534
rect 12910 21522 12962 21534
rect 13246 21586 13298 21598
rect 23886 21586 23938 21598
rect 27582 21586 27634 21598
rect 13906 21534 13918 21586
rect 13970 21534 13982 21586
rect 17378 21534 17390 21586
rect 17442 21534 17454 21586
rect 23426 21534 23438 21586
rect 23490 21534 23502 21586
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 13246 21522 13298 21534
rect 23886 21522 23938 21534
rect 27582 21522 27634 21534
rect 27806 21586 27858 21598
rect 39454 21586 39506 21598
rect 28466 21534 28478 21586
rect 28530 21534 28542 21586
rect 38882 21534 38894 21586
rect 38946 21534 38958 21586
rect 27806 21522 27858 21534
rect 39454 21522 39506 21534
rect 39790 21586 39842 21598
rect 45278 21586 45330 21598
rect 44706 21534 44718 21586
rect 44770 21534 44782 21586
rect 39790 21522 39842 21534
rect 45278 21522 45330 21534
rect 48862 21586 48914 21598
rect 49522 21534 49534 21586
rect 49586 21534 49598 21586
rect 48862 21522 48914 21534
rect 24446 21474 24498 21486
rect 41022 21474 41074 21486
rect 4162 21422 4174 21474
rect 4226 21422 4238 21474
rect 25890 21422 25902 21474
rect 25954 21422 25966 21474
rect 34066 21422 34078 21474
rect 34130 21422 34142 21474
rect 46498 21422 46510 21474
rect 46562 21422 46574 21474
rect 53778 21422 53790 21474
rect 53842 21422 53854 21474
rect 57586 21422 57598 21474
rect 57650 21422 57662 21474
rect 24446 21410 24498 21422
rect 41022 21410 41074 21422
rect 9102 21362 9154 21374
rect 9102 21298 9154 21310
rect 9438 21362 9490 21374
rect 9438 21298 9490 21310
rect 16942 21362 16994 21374
rect 20414 21362 20466 21374
rect 31502 21362 31554 21374
rect 19282 21310 19294 21362
rect 19346 21310 19358 21362
rect 24434 21310 24446 21362
rect 24498 21359 24510 21362
rect 24658 21359 24670 21362
rect 24498 21313 24670 21359
rect 24498 21310 24510 21313
rect 24658 21310 24670 21313
rect 24722 21310 24734 21362
rect 16942 21298 16994 21310
rect 20414 21298 20466 21310
rect 31502 21298 31554 21310
rect 35758 21362 35810 21374
rect 35758 21298 35810 21310
rect 41582 21362 41634 21374
rect 41582 21298 41634 21310
rect 52558 21362 52610 21374
rect 52558 21298 52610 21310
rect 1344 21194 66640 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 66640 21194
rect 1344 21108 66640 21142
rect 48414 21026 48466 21038
rect 48414 20962 48466 20974
rect 13470 20914 13522 20926
rect 15262 20914 15314 20926
rect 19742 20914 19794 20926
rect 20414 20914 20466 20926
rect 23886 20914 23938 20926
rect 4050 20862 4062 20914
rect 4114 20862 4126 20914
rect 8642 20862 8654 20914
rect 8706 20862 8718 20914
rect 11778 20862 11790 20914
rect 11842 20862 11854 20914
rect 13794 20862 13806 20914
rect 13858 20862 13870 20914
rect 15586 20862 15598 20914
rect 15650 20862 15662 20914
rect 20066 20862 20078 20914
rect 20130 20862 20142 20914
rect 20626 20862 20638 20914
rect 20690 20862 20702 20914
rect 22642 20862 22654 20914
rect 22706 20862 22718 20914
rect 13470 20850 13522 20862
rect 15262 20850 15314 20862
rect 19742 20850 19794 20862
rect 20414 20850 20466 20862
rect 23886 20850 23938 20862
rect 28142 20914 28194 20926
rect 37326 20914 37378 20926
rect 49198 20914 49250 20926
rect 36978 20862 36990 20914
rect 37042 20862 37054 20914
rect 38882 20862 38894 20914
rect 38946 20862 38958 20914
rect 42130 20862 42142 20914
rect 42194 20862 42206 20914
rect 43922 20862 43934 20914
rect 43986 20862 43998 20914
rect 49634 20862 49646 20914
rect 49698 20862 49710 20914
rect 51650 20862 51662 20914
rect 51714 20862 51726 20914
rect 53666 20862 53678 20914
rect 53730 20862 53742 20914
rect 28142 20850 28194 20862
rect 37326 20850 37378 20862
rect 49198 20850 49250 20862
rect 7982 20802 8034 20814
rect 7982 20738 8034 20750
rect 8430 20802 8482 20814
rect 8430 20738 8482 20750
rect 15822 20802 15874 20814
rect 27470 20802 27522 20814
rect 34974 20802 35026 20814
rect 16370 20750 16382 20802
rect 16434 20750 16446 20802
rect 27010 20750 27022 20802
rect 27074 20750 27086 20802
rect 34626 20750 34638 20802
rect 34690 20750 34702 20802
rect 15822 20738 15874 20750
rect 27470 20738 27522 20750
rect 34974 20738 35026 20750
rect 44942 20802 44994 20814
rect 45378 20750 45390 20802
rect 45442 20750 45454 20802
rect 51538 20750 51550 20802
rect 51602 20750 51614 20802
rect 44942 20738 44994 20750
rect 24782 20690 24834 20702
rect 3042 20638 3054 20690
rect 3106 20638 3118 20690
rect 9650 20638 9662 20690
rect 9714 20638 9726 20690
rect 10882 20638 10894 20690
rect 10946 20638 10958 20690
rect 21634 20638 21646 20690
rect 21698 20638 21710 20690
rect 24782 20626 24834 20638
rect 32286 20690 32338 20702
rect 44270 20690 44322 20702
rect 39890 20638 39902 20690
rect 39954 20638 39966 20690
rect 43138 20638 43150 20690
rect 43202 20638 43214 20690
rect 50642 20638 50654 20690
rect 50706 20638 50718 20690
rect 54674 20638 54686 20690
rect 54738 20638 54750 20690
rect 32286 20626 32338 20638
rect 44270 20626 44322 20638
rect 19518 20578 19570 20590
rect 18722 20526 18734 20578
rect 18786 20526 18798 20578
rect 19518 20514 19570 20526
rect 23214 20578 23266 20590
rect 23214 20514 23266 20526
rect 23998 20578 24050 20590
rect 23998 20514 24050 20526
rect 31502 20578 31554 20590
rect 47730 20526 47742 20578
rect 47794 20526 47806 20578
rect 31502 20514 31554 20526
rect 1344 20410 66640 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 66640 20410
rect 1344 20324 66640 20358
rect 24222 20242 24274 20254
rect 4834 20190 4846 20242
rect 4898 20190 4910 20242
rect 24222 20178 24274 20190
rect 24670 20242 24722 20254
rect 24670 20178 24722 20190
rect 46286 20242 46338 20254
rect 46286 20178 46338 20190
rect 16830 20130 16882 20142
rect 8306 20078 8318 20130
rect 8370 20078 8382 20130
rect 9874 20078 9886 20130
rect 9938 20078 9950 20130
rect 13458 20078 13470 20130
rect 13522 20078 13534 20130
rect 16482 20078 16494 20130
rect 16546 20078 16558 20130
rect 16830 20066 16882 20078
rect 17502 20130 17554 20142
rect 21982 20130 22034 20142
rect 45054 20130 45106 20142
rect 47070 20130 47122 20142
rect 48190 20130 48242 20142
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 18498 20078 18510 20130
rect 18562 20078 18574 20130
rect 26002 20078 26014 20130
rect 26066 20078 26078 20130
rect 29698 20078 29710 20130
rect 29762 20078 29774 20130
rect 33170 20078 33182 20130
rect 33234 20078 33246 20130
rect 37874 20078 37886 20130
rect 37938 20078 37950 20130
rect 46722 20078 46734 20130
rect 46786 20078 46798 20130
rect 47730 20078 47742 20130
rect 47794 20078 47806 20130
rect 17502 20066 17554 20078
rect 21982 20066 22034 20078
rect 45054 20066 45106 20078
rect 47070 20066 47122 20078
rect 48190 20066 48242 20078
rect 48862 20130 48914 20142
rect 50754 20078 50766 20130
rect 50818 20078 50830 20130
rect 53890 20078 53902 20130
rect 53954 20078 53966 20130
rect 54674 20078 54686 20130
rect 54738 20078 54750 20130
rect 48862 20066 48914 20078
rect 7758 20018 7810 20030
rect 17838 20018 17890 20030
rect 7186 19966 7198 20018
rect 7250 19966 7262 20018
rect 14914 19966 14926 20018
rect 14978 19966 14990 20018
rect 7758 19954 7810 19966
rect 17838 19954 17890 19966
rect 18846 20018 18898 20030
rect 18846 19954 18898 19966
rect 19070 20018 19122 20030
rect 42366 20018 42418 20030
rect 19618 19966 19630 20018
rect 19682 19966 19694 20018
rect 23538 19966 23550 20018
rect 23602 19966 23614 20018
rect 42802 19966 42814 20018
rect 42866 19966 42878 20018
rect 47506 19966 47518 20018
rect 47570 19966 47582 20018
rect 54450 19966 54462 20018
rect 54514 19966 54526 20018
rect 19070 19954 19122 19966
rect 42366 19954 42418 19966
rect 7982 19906 8034 19918
rect 8990 19906 9042 19918
rect 15486 19906 15538 19918
rect 8754 19854 8766 19906
rect 8818 19854 8830 19906
rect 10994 19854 11006 19906
rect 11058 19854 11070 19906
rect 7982 19842 8034 19854
rect 8990 19842 9042 19854
rect 15486 19842 15538 19854
rect 25454 19906 25506 19918
rect 46398 19906 46450 19918
rect 27122 19854 27134 19906
rect 27186 19854 27198 19906
rect 30594 19854 30606 19906
rect 30658 19854 30670 19906
rect 34290 19854 34302 19906
rect 34354 19854 34366 19906
rect 36866 19854 36878 19906
rect 36930 19854 36942 19906
rect 49746 19854 49758 19906
rect 49810 19854 49822 19906
rect 52546 19854 52558 19906
rect 52610 19854 52622 19906
rect 25454 19842 25506 19854
rect 46398 19842 46450 19854
rect 4062 19794 4114 19806
rect 4062 19730 4114 19742
rect 22766 19794 22818 19806
rect 45838 19794 45890 19806
rect 23762 19742 23774 19794
rect 23826 19742 23838 19794
rect 22766 19730 22818 19742
rect 45838 19730 45890 19742
rect 1344 19626 66640 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 66640 19626
rect 1344 19540 66640 19574
rect 20638 19346 20690 19358
rect 8306 19294 8318 19346
rect 8370 19294 8382 19346
rect 11778 19294 11790 19346
rect 11842 19294 11854 19346
rect 16818 19294 16830 19346
rect 16882 19294 16894 19346
rect 19730 19294 19742 19346
rect 19794 19294 19806 19346
rect 20638 19282 20690 19294
rect 21422 19346 21474 19358
rect 21422 19282 21474 19294
rect 21870 19346 21922 19358
rect 21870 19282 21922 19294
rect 26574 19346 26626 19358
rect 43710 19346 43762 19358
rect 31042 19294 31054 19346
rect 31106 19294 31118 19346
rect 33506 19294 33518 19346
rect 33570 19294 33582 19346
rect 38322 19294 38334 19346
rect 38386 19294 38398 19346
rect 41570 19294 41582 19346
rect 41634 19294 41646 19346
rect 26574 19282 26626 19294
rect 43710 19282 43762 19294
rect 44382 19346 44434 19358
rect 44382 19282 44434 19294
rect 45054 19346 45106 19358
rect 45054 19282 45106 19294
rect 45502 19346 45554 19358
rect 51102 19346 51154 19358
rect 46050 19294 46062 19346
rect 46114 19294 46126 19346
rect 48626 19294 48638 19346
rect 48690 19294 48702 19346
rect 50866 19294 50878 19346
rect 50930 19294 50942 19346
rect 54002 19294 54014 19346
rect 54066 19294 54078 19346
rect 45502 19282 45554 19294
rect 51102 19282 51154 19294
rect 22542 19234 22594 19246
rect 23090 19182 23102 19234
rect 23154 19182 23166 19234
rect 22542 19170 22594 19182
rect 25454 19122 25506 19134
rect 9538 19070 9550 19122
rect 9602 19070 9614 19122
rect 10546 19070 10558 19122
rect 10610 19070 10622 19122
rect 15586 19070 15598 19122
rect 15650 19070 15662 19122
rect 18722 19070 18734 19122
rect 18786 19070 18798 19122
rect 30034 19070 30046 19122
rect 30098 19070 30110 19122
rect 34514 19070 34526 19122
rect 34578 19070 34590 19122
rect 39330 19070 39342 19122
rect 39394 19070 39406 19122
rect 42578 19070 42590 19122
rect 42642 19070 42654 19122
rect 47058 19070 47070 19122
rect 47122 19070 47134 19122
rect 49634 19070 49646 19122
rect 49698 19070 49710 19122
rect 55010 19070 55022 19122
rect 55074 19070 55086 19122
rect 25454 19058 25506 19070
rect 20302 19010 20354 19022
rect 20302 18946 20354 18958
rect 21982 19010 22034 19022
rect 21982 18946 22034 18958
rect 26238 19010 26290 19022
rect 26238 18946 26290 18958
rect 43598 19010 43650 19022
rect 43598 18946 43650 18958
rect 1344 18842 66640 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 66640 18842
rect 1344 18756 66640 18790
rect 23886 18674 23938 18686
rect 23886 18610 23938 18622
rect 46846 18562 46898 18574
rect 4050 18510 4062 18562
rect 4114 18510 4126 18562
rect 6626 18510 6638 18562
rect 6690 18510 6702 18562
rect 9874 18510 9886 18562
rect 9938 18510 9950 18562
rect 13346 18510 13358 18562
rect 13410 18510 13422 18562
rect 18274 18510 18286 18562
rect 18338 18510 18350 18562
rect 22978 18510 22990 18562
rect 23042 18510 23054 18562
rect 28914 18510 28926 18562
rect 28978 18510 28990 18562
rect 29474 18510 29486 18562
rect 29538 18510 29550 18562
rect 33618 18510 33630 18562
rect 33682 18510 33694 18562
rect 38434 18510 38446 18562
rect 38498 18510 38510 18562
rect 42914 18510 42926 18562
rect 42978 18510 42990 18562
rect 45714 18510 45726 18562
rect 45778 18510 45790 18562
rect 46846 18498 46898 18510
rect 47854 18562 47906 18574
rect 51538 18510 51550 18562
rect 51602 18510 51614 18562
rect 47854 18498 47906 18510
rect 47170 18398 47182 18450
rect 47234 18398 47246 18450
rect 5170 18286 5182 18338
rect 5234 18286 5246 18338
rect 7858 18286 7870 18338
rect 7922 18286 7934 18338
rect 11106 18286 11118 18338
rect 11170 18286 11182 18338
rect 14466 18286 14478 18338
rect 14530 18286 14542 18338
rect 19506 18286 19518 18338
rect 19570 18286 19582 18338
rect 21858 18286 21870 18338
rect 21922 18286 21934 18338
rect 27794 18286 27806 18338
rect 27858 18286 27870 18338
rect 30818 18286 30830 18338
rect 30882 18286 30894 18338
rect 34738 18286 34750 18338
rect 34802 18286 34814 18338
rect 37314 18286 37326 18338
rect 37378 18286 37390 18338
rect 41906 18286 41918 18338
rect 41970 18286 41982 18338
rect 44706 18286 44718 18338
rect 44770 18286 44782 18338
rect 48066 18286 48078 18338
rect 48130 18286 48142 18338
rect 50194 18286 50206 18338
rect 50258 18286 50270 18338
rect 1344 18058 66640 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 66640 18058
rect 1344 17972 66640 18006
rect 8642 17726 8654 17778
rect 8706 17726 8718 17778
rect 11890 17726 11902 17778
rect 11954 17726 11966 17778
rect 16594 17726 16606 17778
rect 16658 17726 16670 17778
rect 19730 17726 19742 17778
rect 19794 17726 19806 17778
rect 24770 17726 24782 17778
rect 24834 17726 24846 17778
rect 27122 17726 27134 17778
rect 27186 17726 27198 17778
rect 32386 17726 32398 17778
rect 32450 17726 32462 17778
rect 35410 17726 35422 17778
rect 35474 17726 35486 17778
rect 40114 17726 40126 17778
rect 40178 17726 40190 17778
rect 45826 17726 45838 17778
rect 45890 17726 45902 17778
rect 48626 17726 48638 17778
rect 48690 17726 48702 17778
rect 9650 17502 9662 17554
rect 9714 17502 9726 17554
rect 10770 17502 10782 17554
rect 10834 17502 10846 17554
rect 17490 17502 17502 17554
rect 17554 17502 17566 17554
rect 18722 17502 18734 17554
rect 18786 17502 18798 17554
rect 23762 17502 23774 17554
rect 23826 17502 23838 17554
rect 28354 17502 28366 17554
rect 28418 17502 28430 17554
rect 31490 17502 31502 17554
rect 31554 17502 31566 17554
rect 34402 17502 34414 17554
rect 34466 17502 34478 17554
rect 41122 17502 41134 17554
rect 41186 17502 41198 17554
rect 47058 17502 47070 17554
rect 47122 17502 47134 17554
rect 49634 17502 49646 17554
rect 49698 17502 49710 17554
rect 1344 17274 66640 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 66640 17274
rect 1344 17188 66640 17222
rect 12674 16942 12686 16994
rect 12738 16942 12750 16994
rect 16706 16942 16718 16994
rect 16770 16942 16782 16994
rect 18386 16942 18398 16994
rect 18450 16942 18462 16994
rect 20962 16942 20974 16994
rect 21026 16942 21038 16994
rect 28690 16942 28702 16994
rect 28754 16942 28766 16994
rect 29362 16942 29374 16994
rect 29426 16942 29438 16994
rect 35298 16942 35310 16994
rect 35362 16942 35374 16994
rect 38882 16942 38894 16994
rect 38946 16942 38958 16994
rect 43026 16942 43038 16994
rect 43090 16942 43102 16994
rect 46050 16942 46062 16994
rect 46114 16942 46126 16994
rect 11330 16718 11342 16770
rect 11394 16718 11406 16770
rect 15586 16718 15598 16770
rect 15650 16718 15662 16770
rect 19394 16718 19406 16770
rect 19458 16718 19470 16770
rect 22306 16718 22318 16770
rect 22370 16718 22382 16770
rect 27458 16718 27470 16770
rect 27522 16718 27534 16770
rect 30706 16718 30718 16770
rect 30770 16718 30782 16770
rect 34178 16718 34190 16770
rect 34242 16718 34254 16770
rect 38098 16718 38110 16770
rect 38162 16718 38174 16770
rect 41906 16718 41918 16770
rect 41970 16718 41982 16770
rect 44706 16718 44718 16770
rect 44770 16718 44782 16770
rect 1344 16490 66640 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 66640 16490
rect 1344 16404 66640 16438
rect 9986 16158 9998 16210
rect 10050 16158 10062 16210
rect 14802 16158 14814 16210
rect 14866 16158 14878 16210
rect 18722 16158 18734 16210
rect 18786 16158 18798 16210
rect 22642 16158 22654 16210
rect 22706 16158 22718 16210
rect 26450 16158 26462 16210
rect 26514 16158 26526 16210
rect 31938 16158 31950 16210
rect 32002 16158 32014 16210
rect 35298 16158 35310 16210
rect 35362 16158 35374 16210
rect 39106 16158 39118 16210
rect 39170 16158 39182 16210
rect 42578 16158 42590 16210
rect 42642 16158 42654 16210
rect 10882 15934 10894 15986
rect 10946 15934 10958 15986
rect 16146 15934 16158 15986
rect 16210 15934 16222 15986
rect 19730 15934 19742 15986
rect 19794 15934 19806 15986
rect 23650 15934 23662 15986
rect 23714 15934 23726 15986
rect 27234 15934 27246 15986
rect 27298 15934 27310 15986
rect 33282 15934 33294 15986
rect 33346 15934 33358 15986
rect 33954 15934 33966 15986
rect 34018 15934 34030 15986
rect 37986 15934 37998 15986
rect 38050 15934 38062 15986
rect 43698 15934 43710 15986
rect 43762 15934 43774 15986
rect 1344 15706 66640 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 66640 15706
rect 1344 15620 66640 15654
rect 21298 15374 21310 15426
rect 21362 15374 21374 15426
rect 22530 15374 22542 15426
rect 22594 15374 22606 15426
rect 29586 15374 29598 15426
rect 29650 15374 29662 15426
rect 32050 15374 32062 15426
rect 32114 15374 32126 15426
rect 36754 15374 36766 15426
rect 36818 15374 36830 15426
rect 20290 15150 20302 15202
rect 20354 15150 20366 15202
rect 23538 15150 23550 15202
rect 23602 15150 23614 15202
rect 28242 15150 28254 15202
rect 28306 15150 28318 15202
rect 31154 15150 31166 15202
rect 31218 15150 31230 15202
rect 35746 15150 35758 15202
rect 35810 15150 35822 15202
rect 1344 14922 66640 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 66640 14922
rect 1344 14836 66640 14870
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 23314 14590 23326 14642
rect 23378 14590 23390 14642
rect 27346 14590 27358 14642
rect 27410 14590 27422 14642
rect 30146 14590 30158 14642
rect 30210 14590 30222 14642
rect 19170 14366 19182 14418
rect 19234 14366 19246 14418
rect 24322 14366 24334 14418
rect 24386 14366 24398 14418
rect 26338 14366 26350 14418
rect 26402 14366 26414 14418
rect 31266 14366 31278 14418
rect 31330 14366 31342 14418
rect 1344 14138 66640 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 66640 14138
rect 1344 14052 66640 14086
rect 1344 13354 66640 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 66640 13354
rect 1344 13268 66640 13302
rect 1344 12570 66640 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 66640 12570
rect 1344 12484 66640 12518
rect 1344 11786 66640 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 66640 11786
rect 1344 11700 66640 11734
rect 1344 11002 66640 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 66640 11002
rect 1344 10916 66640 10950
rect 1344 10218 66640 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 66640 10218
rect 1344 10132 66640 10166
rect 1344 9434 66640 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 66640 9434
rect 1344 9348 66640 9382
rect 1344 8650 66640 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 66640 8650
rect 1344 8564 66640 8598
rect 1344 7866 66640 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 66640 7866
rect 1344 7780 66640 7814
rect 1344 7082 66640 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 66640 7082
rect 1344 6996 66640 7030
rect 1344 6298 66640 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 66640 6298
rect 1344 6212 66640 6246
rect 1344 5514 66640 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 66640 5514
rect 1344 5428 66640 5462
rect 1344 4730 66640 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 66640 4730
rect 1344 4644 66640 4678
rect 1344 3946 66640 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 66640 3946
rect 1344 3860 66640 3894
rect 40574 3330 40626 3342
rect 40574 3266 40626 3278
rect 41246 3330 41298 3342
rect 41246 3266 41298 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 44606 3330 44658 3342
rect 44606 3266 44658 3278
rect 48638 3330 48690 3342
rect 48638 3266 48690 3278
rect 55022 3330 55074 3342
rect 55022 3266 55074 3278
rect 1344 3162 66640 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 66640 3162
rect 1344 3076 66640 3110
<< via1 >>
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 56702 64094 56754 64146
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 66222 62862 66274 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 43710 54574 43762 54626
rect 42702 54350 42754 54402
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 30382 53790 30434 53842
rect 33630 53790 33682 53842
rect 38558 53790 38610 53842
rect 41358 53790 41410 53842
rect 45838 53790 45890 53842
rect 31390 53566 31442 53618
rect 34638 53566 34690 53618
rect 39566 53566 39618 53618
rect 42366 53566 42418 53618
rect 47070 53566 47122 53618
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 32062 53006 32114 53058
rect 35870 53006 35922 53058
rect 38670 53006 38722 53058
rect 41246 53006 41298 53058
rect 45950 53006 46002 53058
rect 51102 53006 51154 53058
rect 31054 52782 31106 52834
rect 34862 52782 34914 52834
rect 37662 52782 37714 52834
rect 42590 52782 42642 52834
rect 44942 52782 44994 52834
rect 50094 52782 50146 52834
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 27246 52222 27298 52274
rect 32062 52222 32114 52274
rect 34414 52222 34466 52274
rect 37998 52222 38050 52274
rect 40798 52222 40850 52274
rect 46062 52222 46114 52274
rect 48638 52222 48690 52274
rect 28142 51998 28194 52050
rect 30718 51998 30770 52050
rect 35422 51998 35474 52050
rect 39118 51998 39170 52050
rect 41806 51998 41858 52050
rect 47182 51998 47234 52050
rect 49870 51998 49922 52050
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 23662 51438 23714 51490
rect 28478 51438 28530 51490
rect 29038 51438 29090 51490
rect 37774 51438 37826 51490
rect 43150 51438 43202 51490
rect 45726 51438 45778 51490
rect 50766 51438 50818 51490
rect 53790 51438 53842 51490
rect 22318 51214 22370 51266
rect 27134 51214 27186 51266
rect 30158 51214 30210 51266
rect 36766 51214 36818 51266
rect 41918 51214 41970 51266
rect 44718 51214 44770 51266
rect 49758 51214 49810 51266
rect 52558 51214 52610 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 24558 50654 24610 50706
rect 27582 50654 27634 50706
rect 32622 50654 32674 50706
rect 40014 50654 40066 50706
rect 42590 50654 42642 50706
rect 45838 50654 45890 50706
rect 48638 50654 48690 50706
rect 54014 50654 54066 50706
rect 56814 50654 56866 50706
rect 25342 50430 25394 50482
rect 26574 50430 26626 50482
rect 33966 50430 34018 50482
rect 38894 50430 38946 50482
rect 43934 50430 43986 50482
rect 47070 50430 47122 50482
rect 49646 50430 49698 50482
rect 55134 50430 55186 50482
rect 57822 50430 57874 50482
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 45390 49982 45442 50034
rect 45950 49982 46002 50034
rect 53342 49982 53394 50034
rect 53902 49982 53954 50034
rect 23886 49870 23938 49922
rect 29374 49870 29426 49922
rect 32062 49870 32114 49922
rect 35310 49870 35362 49922
rect 36990 49870 37042 49922
rect 46846 49870 46898 49922
rect 54126 49870 54178 49922
rect 58830 49870 58882 49922
rect 25454 49758 25506 49810
rect 42254 49758 42306 49810
rect 42926 49758 42978 49810
rect 46398 49758 46450 49810
rect 47070 49758 47122 49810
rect 50318 49758 50370 49810
rect 50878 49758 50930 49810
rect 54350 49758 54402 49810
rect 22542 49646 22594 49698
rect 25230 49646 25282 49698
rect 26126 49646 26178 49698
rect 27918 49646 27970 49698
rect 28254 49646 28306 49698
rect 31054 49646 31106 49698
rect 34078 49646 34130 49698
rect 38110 49646 38162 49698
rect 46174 49646 46226 49698
rect 47518 49646 47570 49698
rect 47854 49646 47906 49698
rect 49422 49646 49474 49698
rect 49646 49646 49698 49698
rect 49982 49646 50034 49698
rect 55022 49646 55074 49698
rect 55470 49646 55522 49698
rect 57598 49646 57650 49698
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 27918 49198 27970 49250
rect 35198 49198 35250 49250
rect 41694 49198 41746 49250
rect 48638 49198 48690 49250
rect 55358 49198 55410 49250
rect 55582 49198 55634 49250
rect 19630 49086 19682 49138
rect 22878 49086 22930 49138
rect 28142 49086 28194 49138
rect 49870 49086 49922 49138
rect 53678 49086 53730 49138
rect 55582 49086 55634 49138
rect 56478 49086 56530 49138
rect 24334 48974 24386 49026
rect 24782 48974 24834 49026
rect 31726 48974 31778 49026
rect 32062 48974 32114 49026
rect 36094 48974 36146 49026
rect 37998 48974 38050 49026
rect 38670 48974 38722 49026
rect 43374 48974 43426 49026
rect 44942 48974 44994 49026
rect 45614 48974 45666 49026
rect 51886 48974 51938 49026
rect 52782 48974 52834 49026
rect 18510 48862 18562 48914
rect 21534 48862 21586 48914
rect 29262 48862 29314 48914
rect 29598 48862 29650 48914
rect 30270 48862 30322 48914
rect 42254 48862 42306 48914
rect 42926 48862 42978 48914
rect 43598 48862 43650 48914
rect 47854 48862 47906 48914
rect 50878 48862 50930 48914
rect 51662 48862 51714 48914
rect 54686 48862 54738 48914
rect 57486 48862 57538 48914
rect 27358 48750 27410 48802
rect 28254 48750 28306 48802
rect 30158 48750 30210 48802
rect 34414 48750 34466 48802
rect 36094 48750 36146 48802
rect 41134 48750 41186 48802
rect 42142 48750 42194 48802
rect 42814 48750 42866 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 29262 48414 29314 48466
rect 29934 48414 29986 48466
rect 36094 48414 36146 48466
rect 39902 48414 39954 48466
rect 40462 48414 40514 48466
rect 44830 48414 44882 48466
rect 45390 48414 45442 48466
rect 48638 48414 48690 48466
rect 49422 48414 49474 48466
rect 19518 48302 19570 48354
rect 22654 48302 22706 48354
rect 41246 48302 41298 48354
rect 54574 48302 54626 48354
rect 55358 48302 55410 48354
rect 58830 48302 58882 48354
rect 25902 48190 25954 48242
rect 26462 48190 26514 48242
rect 26910 48190 26962 48242
rect 30830 48190 30882 48242
rect 31950 48190 32002 48242
rect 33070 48190 33122 48242
rect 36094 48190 36146 48242
rect 36766 48190 36818 48242
rect 37438 48190 37490 48242
rect 41918 48190 41970 48242
rect 42254 48190 42306 48242
rect 45614 48190 45666 48242
rect 51774 48190 51826 48242
rect 52334 48190 52386 48242
rect 53118 48190 53170 48242
rect 20862 48078 20914 48130
rect 23662 48078 23714 48130
rect 25342 48078 25394 48130
rect 25678 48078 25730 48130
rect 30942 48078 30994 48130
rect 31614 48078 31666 48130
rect 32622 48078 32674 48130
rect 35422 48078 35474 48130
rect 40910 48078 40962 48130
rect 47966 48078 48018 48130
rect 52670 48078 52722 48130
rect 53566 48078 53618 48130
rect 55582 48078 55634 48130
rect 57598 48078 57650 48130
rect 52670 47966 52722 48018
rect 53118 47966 53170 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 28702 47630 28754 47682
rect 32734 47630 32786 47682
rect 36542 47630 36594 47682
rect 48414 47630 48466 47682
rect 52222 47630 52274 47682
rect 56254 47630 56306 47682
rect 19518 47518 19570 47570
rect 23438 47518 23490 47570
rect 40462 47518 40514 47570
rect 44270 47518 44322 47570
rect 57486 47518 57538 47570
rect 25118 47406 25170 47458
rect 25566 47406 25618 47458
rect 29038 47406 29090 47458
rect 29710 47406 29762 47458
rect 32846 47406 32898 47458
rect 33518 47406 33570 47458
rect 42254 47406 42306 47458
rect 44942 47406 44994 47458
rect 45390 47406 45442 47458
rect 48526 47406 48578 47458
rect 49198 47406 49250 47458
rect 52670 47406 52722 47458
rect 53118 47406 53170 47458
rect 18622 47294 18674 47346
rect 21646 47294 21698 47346
rect 21982 47294 22034 47346
rect 22430 47294 22482 47346
rect 24670 47294 24722 47346
rect 58494 47294 58546 47346
rect 28142 47182 28194 47234
rect 32062 47182 32114 47234
rect 35870 47182 35922 47234
rect 42926 47182 42978 47234
rect 47630 47182 47682 47234
rect 51550 47182 51602 47234
rect 55582 47182 55634 47234
rect 56590 47182 56642 47234
rect 59390 47182 59442 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 23886 46846 23938 46898
rect 30942 46846 30994 46898
rect 31614 46846 31666 46898
rect 38894 46846 38946 46898
rect 39454 46846 39506 46898
rect 43710 46846 43762 46898
rect 44494 46846 44546 46898
rect 44606 46846 44658 46898
rect 52446 46846 52498 46898
rect 17726 46734 17778 46786
rect 25678 46734 25730 46786
rect 35422 46734 35474 46786
rect 40014 46734 40066 46786
rect 40350 46734 40402 46786
rect 45390 46734 45442 46786
rect 51550 46734 51602 46786
rect 53230 46734 53282 46786
rect 58830 46734 58882 46786
rect 59390 46734 59442 46786
rect 20862 46622 20914 46674
rect 21310 46622 21362 46674
rect 28142 46622 28194 46674
rect 28590 46622 28642 46674
rect 32286 46622 32338 46674
rect 35982 46622 36034 46674
rect 36430 46622 36482 46674
rect 40798 46622 40850 46674
rect 41470 46622 41522 46674
rect 47742 46622 47794 46674
rect 48078 46622 48130 46674
rect 48638 46622 48690 46674
rect 49310 46622 49362 46674
rect 55582 46622 55634 46674
rect 56142 46622 56194 46674
rect 59614 46622 59666 46674
rect 18846 46510 18898 46562
rect 26574 46510 26626 46562
rect 32510 46510 32562 46562
rect 34302 46510 34354 46562
rect 56702 46510 56754 46562
rect 57150 46510 57202 46562
rect 57598 46510 57650 46562
rect 24446 46398 24498 46450
rect 52334 46398 52386 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 17166 46062 17218 46114
rect 24894 46062 24946 46114
rect 28702 46062 28754 46114
rect 29038 46062 29090 46114
rect 36542 46062 36594 46114
rect 37438 46062 37490 46114
rect 56254 46062 56306 46114
rect 43598 45950 43650 46002
rect 44942 45950 44994 46002
rect 57486 45950 57538 46002
rect 20302 45838 20354 45890
rect 20862 45838 20914 45890
rect 21422 45838 21474 45890
rect 21758 45838 21810 45890
rect 25118 45838 25170 45890
rect 25566 45838 25618 45890
rect 32062 45838 32114 45890
rect 32734 45838 32786 45890
rect 32846 45838 32898 45890
rect 33406 45838 33458 45890
rect 40462 45838 40514 45890
rect 40910 45838 40962 45890
rect 41806 45838 41858 45890
rect 50430 45838 50482 45890
rect 52670 45838 52722 45890
rect 53118 45838 53170 45890
rect 59278 45838 59330 45890
rect 59502 45838 59554 45890
rect 27918 45726 27970 45778
rect 29822 45726 29874 45778
rect 35758 45726 35810 45778
rect 38222 45726 38274 45778
rect 46286 45726 46338 45778
rect 58494 45726 58546 45778
rect 17726 45614 17778 45666
rect 24222 45614 24274 45666
rect 45726 45614 45778 45666
rect 51886 45614 51938 45666
rect 55694 45614 55746 45666
rect 56590 45614 56642 45666
rect 57038 45614 57090 45666
rect 60622 45614 60674 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 23662 45278 23714 45330
rect 24446 45278 24498 45330
rect 32958 45278 33010 45330
rect 33742 45278 33794 45330
rect 39902 45278 39954 45330
rect 40462 45278 40514 45330
rect 41022 45278 41074 45330
rect 42366 45278 42418 45330
rect 47294 45278 47346 45330
rect 48190 45278 48242 45330
rect 52334 45278 52386 45330
rect 56142 45278 56194 45330
rect 17726 45166 17778 45218
rect 18398 45166 18450 45218
rect 28590 45166 28642 45218
rect 32174 45166 32226 45218
rect 41470 45166 41522 45218
rect 43150 45166 43202 45218
rect 46846 45166 46898 45218
rect 51550 45166 51602 45218
rect 55358 45166 55410 45218
rect 58830 45166 58882 45218
rect 61406 45166 61458 45218
rect 17502 45054 17554 45106
rect 20862 45054 20914 45106
rect 21310 45054 21362 45106
rect 26686 45054 26738 45106
rect 30942 45054 30994 45106
rect 32398 45054 32450 45106
rect 35982 45054 36034 45106
rect 36430 45054 36482 45106
rect 36766 45054 36818 45106
rect 37438 45054 37490 45106
rect 41694 45054 41746 45106
rect 45502 45054 45554 45106
rect 45950 45054 46002 45106
rect 48862 45054 48914 45106
rect 49310 45054 49362 45106
rect 52558 45054 52610 45106
rect 53006 45054 53058 45106
rect 16942 44942 16994 44994
rect 19518 44942 19570 44994
rect 46510 44942 46562 44994
rect 47182 44942 47234 44994
rect 56702 44942 56754 44994
rect 57150 44942 57202 44994
rect 57598 44942 57650 44994
rect 59502 44942 59554 44994
rect 60398 44942 60450 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 17166 44494 17218 44546
rect 28030 44494 28082 44546
rect 35198 44494 35250 44546
rect 40574 44494 40626 44546
rect 49646 44494 49698 44546
rect 14814 44382 14866 44434
rect 23102 44382 23154 44434
rect 24110 44382 24162 44434
rect 29486 44382 29538 44434
rect 29822 44382 29874 44434
rect 41806 44382 41858 44434
rect 45166 44382 45218 44434
rect 49870 44382 49922 44434
rect 50206 44382 50258 44434
rect 51102 44382 51154 44434
rect 51438 44382 51490 44434
rect 57150 44382 57202 44434
rect 58942 44382 58994 44434
rect 61518 44382 61570 44434
rect 20190 44270 20242 44322
rect 20862 44270 20914 44322
rect 24558 44270 24610 44322
rect 24894 44270 24946 44322
rect 30494 44270 30546 44322
rect 31502 44270 31554 44322
rect 32062 44270 32114 44322
rect 36990 44270 37042 44322
rect 37438 44270 37490 44322
rect 45390 44270 45442 44322
rect 45950 44270 46002 44322
rect 46622 44270 46674 44322
rect 52670 44270 52722 44322
rect 58494 44270 58546 44322
rect 16158 44158 16210 44210
rect 22094 44158 22146 44210
rect 28254 44158 28306 44210
rect 30270 44158 30322 44210
rect 35982 44158 36034 44210
rect 36318 44158 36370 44210
rect 42814 44158 42866 44210
rect 43598 44158 43650 44210
rect 58270 44158 58322 44210
rect 59278 44158 59330 44210
rect 62526 44158 62578 44210
rect 17726 44046 17778 44098
rect 27470 44046 27522 44098
rect 28366 44046 28418 44098
rect 34638 44046 34690 44098
rect 39902 44046 39954 44098
rect 40910 44046 40962 44098
rect 43710 44046 43762 44098
rect 49086 44046 49138 44098
rect 50654 44046 50706 44098
rect 51550 44046 51602 44098
rect 59726 44046 59778 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 43710 43710 43762 43762
rect 59502 43710 59554 43762
rect 14814 43598 14866 43650
rect 17726 43598 17778 43650
rect 19406 43598 19458 43650
rect 20750 43598 20802 43650
rect 21534 43598 21586 43650
rect 25678 43598 25730 43650
rect 27918 43598 27970 43650
rect 28702 43598 28754 43650
rect 33070 43598 33122 43650
rect 34190 43598 34242 43650
rect 44494 43598 44546 43650
rect 47742 43598 47794 43650
rect 48190 43598 48242 43650
rect 49198 43598 49250 43650
rect 49534 43598 49586 43650
rect 50766 43598 50818 43650
rect 51774 43598 51826 43650
rect 54910 43598 54962 43650
rect 58830 43598 58882 43650
rect 61406 43598 61458 43650
rect 17502 43486 17554 43538
rect 23774 43486 23826 43538
rect 24446 43486 24498 43538
rect 31054 43486 31106 43538
rect 31390 43486 31442 43538
rect 32398 43486 32450 43538
rect 33294 43486 33346 43538
rect 36542 43486 36594 43538
rect 40910 43486 40962 43538
rect 41470 43486 41522 43538
rect 45166 43486 45218 43538
rect 49982 43486 50034 43538
rect 50990 43486 51042 43538
rect 54126 43486 54178 43538
rect 54686 43486 54738 43538
rect 55134 43486 55186 43538
rect 55918 43486 55970 43538
rect 15822 43374 15874 43426
rect 18062 43374 18114 43426
rect 26686 43374 26738 43426
rect 27694 43374 27746 43426
rect 32174 43374 32226 43426
rect 33854 43374 33906 43426
rect 39006 43374 39058 43426
rect 45726 43374 45778 43426
rect 48862 43374 48914 43426
rect 50206 43374 50258 43426
rect 55694 43374 55746 43426
rect 56702 43374 56754 43426
rect 57150 43374 57202 43426
rect 57598 43374 57650 43426
rect 60398 43374 60450 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 17614 42926 17666 42978
rect 17950 42926 18002 42978
rect 21198 42926 21250 42978
rect 32734 42926 32786 42978
rect 40574 42926 40626 42978
rect 44382 42926 44434 42978
rect 52222 42926 52274 42978
rect 60062 42926 60114 42978
rect 16830 42814 16882 42866
rect 17950 42814 18002 42866
rect 19518 42814 19570 42866
rect 61518 42814 61570 42866
rect 24222 42702 24274 42754
rect 24894 42702 24946 42754
rect 28030 42702 28082 42754
rect 28590 42702 28642 42754
rect 29262 42702 29314 42754
rect 29710 42702 29762 42754
rect 32846 42702 32898 42754
rect 35982 42702 36034 42754
rect 36430 42702 36482 42754
rect 36878 42702 36930 42754
rect 37438 42702 37490 42754
rect 40910 42702 40962 42754
rect 41246 42702 41298 42754
rect 44942 42702 44994 42754
rect 45390 42702 45442 42754
rect 48638 42702 48690 42754
rect 49086 42702 49138 42754
rect 52782 42702 52834 42754
rect 53118 42702 53170 42754
rect 56590 42702 56642 42754
rect 57038 42702 57090 42754
rect 15934 42590 15986 42642
rect 18734 42590 18786 42642
rect 25790 42590 25842 42642
rect 33630 42590 33682 42642
rect 48414 42590 48466 42642
rect 55470 42590 55522 42642
rect 56254 42590 56306 42642
rect 62526 42590 62578 42642
rect 21982 42478 22034 42530
rect 25006 42478 25058 42530
rect 32174 42478 32226 42530
rect 40014 42478 40066 42530
rect 43598 42478 43650 42530
rect 47630 42478 47682 42530
rect 51662 42478 51714 42530
rect 59390 42478 59442 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 23102 42142 23154 42194
rect 43934 42142 43986 42194
rect 51550 42142 51602 42194
rect 55358 42142 55410 42194
rect 12014 42030 12066 42082
rect 16718 42030 16770 42082
rect 17838 42030 17890 42082
rect 30606 42030 30658 42082
rect 36654 42030 36706 42082
rect 47518 42030 47570 42082
rect 58830 42030 58882 42082
rect 61406 42030 61458 42082
rect 20302 41918 20354 41970
rect 20638 41918 20690 41970
rect 23774 41918 23826 41970
rect 23998 41918 24050 41970
rect 27134 41918 27186 41970
rect 27470 41918 27522 41970
rect 27918 41918 27970 41970
rect 28254 41918 28306 41970
rect 31390 41918 31442 41970
rect 31726 41918 31778 41970
rect 32510 41918 32562 41970
rect 33294 41918 33346 41970
rect 35870 41918 35922 41970
rect 38894 41918 38946 41970
rect 39566 41918 39618 41970
rect 40798 41918 40850 41970
rect 41470 41918 41522 41970
rect 44494 41918 44546 41970
rect 44830 41918 44882 41970
rect 45278 41918 45330 41970
rect 48302 41918 48354 41970
rect 48638 41918 48690 41970
rect 49310 41918 49362 41970
rect 52334 41918 52386 41970
rect 52446 41918 52498 41970
rect 53006 41918 53058 41970
rect 56142 41918 56194 41970
rect 56702 41918 56754 41970
rect 59502 41918 59554 41970
rect 62414 41918 62466 41970
rect 13022 41806 13074 41858
rect 15374 41806 15426 41858
rect 18846 41806 18898 41858
rect 24334 41806 24386 41858
rect 25454 41806 25506 41858
rect 25790 41806 25842 41858
rect 26126 41806 26178 41858
rect 26462 41806 26514 41858
rect 26798 41806 26850 41858
rect 31838 41806 31890 41858
rect 39902 41806 39954 41858
rect 40126 41806 40178 41858
rect 57150 41806 57202 41858
rect 57598 41806 57650 41858
rect 60398 41806 60450 41858
rect 62190 41806 62242 41858
rect 62974 41806 63026 41858
rect 34078 41694 34130 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 25006 41358 25058 41410
rect 35870 41358 35922 41410
rect 56254 41358 56306 41410
rect 11902 41246 11954 41298
rect 16830 41246 16882 41298
rect 19742 41246 19794 41298
rect 24446 41246 24498 41298
rect 24782 41246 24834 41298
rect 30942 41246 30994 41298
rect 36094 41246 36146 41298
rect 36990 41246 37042 41298
rect 38222 41246 38274 41298
rect 43374 41246 43426 41298
rect 45502 41246 45554 41298
rect 46174 41246 46226 41298
rect 46510 41246 46562 41298
rect 46846 41246 46898 41298
rect 47182 41246 47234 41298
rect 51662 41246 51714 41298
rect 52110 41246 52162 41298
rect 56702 41246 56754 41298
rect 57038 41246 57090 41298
rect 57486 41246 57538 41298
rect 59278 41246 59330 41298
rect 59614 41246 59666 41298
rect 61742 41246 61794 41298
rect 23550 41134 23602 41186
rect 28030 41134 28082 41186
rect 28590 41134 28642 41186
rect 32174 41134 32226 41186
rect 32734 41134 32786 41186
rect 39006 41134 39058 41186
rect 39454 41134 39506 41186
rect 42478 41134 42530 41186
rect 45726 41134 45778 41186
rect 47630 41134 47682 41186
rect 48078 41134 48130 41186
rect 51438 41134 51490 41186
rect 52558 41134 52610 41186
rect 53230 41134 53282 41186
rect 10782 41022 10834 41074
rect 15934 41022 15986 41074
rect 18734 41022 18786 41074
rect 25790 41022 25842 41074
rect 29934 41022 29986 41074
rect 36430 41022 36482 41074
rect 38558 41022 38610 41074
rect 42702 41022 42754 41074
rect 43038 41022 43090 41074
rect 43710 41022 43762 41074
rect 44830 41022 44882 41074
rect 45166 41022 45218 41074
rect 58494 41022 58546 41074
rect 62526 41022 62578 41074
rect 20750 40910 20802 40962
rect 22878 40910 22930 40962
rect 35198 40910 35250 40962
rect 37102 40910 37154 40962
rect 41694 40910 41746 40962
rect 50318 40910 50370 40962
rect 51102 40910 51154 40962
rect 55694 40910 55746 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 11678 40574 11730 40626
rect 12238 40574 12290 40626
rect 16382 40574 16434 40626
rect 21086 40574 21138 40626
rect 28142 40574 28194 40626
rect 31838 40574 31890 40626
rect 32622 40574 32674 40626
rect 36430 40574 36482 40626
rect 37214 40574 37266 40626
rect 47406 40574 47458 40626
rect 47966 40574 48018 40626
rect 56142 40574 56194 40626
rect 56702 40574 56754 40626
rect 57150 40574 57202 40626
rect 59502 40574 59554 40626
rect 17838 40462 17890 40514
rect 18846 40462 18898 40514
rect 21870 40462 21922 40514
rect 25566 40462 25618 40514
rect 26462 40462 26514 40514
rect 39454 40462 39506 40514
rect 42926 40462 42978 40514
rect 43710 40462 43762 40514
rect 44046 40462 44098 40514
rect 55358 40462 55410 40514
rect 58830 40462 58882 40514
rect 61406 40462 61458 40514
rect 14702 40350 14754 40402
rect 15150 40350 15202 40402
rect 16494 40350 16546 40402
rect 17502 40350 17554 40402
rect 20302 40350 20354 40402
rect 24110 40350 24162 40402
rect 24670 40350 24722 40402
rect 25790 40350 25842 40402
rect 28926 40350 28978 40402
rect 29486 40350 29538 40402
rect 33518 40350 33570 40402
rect 34190 40350 34242 40402
rect 44494 40350 44546 40402
rect 44942 40350 44994 40402
rect 49198 40350 49250 40402
rect 51998 40350 52050 40402
rect 52446 40350 52498 40402
rect 53118 40350 53170 40402
rect 19854 40238 19906 40290
rect 27694 40238 27746 40290
rect 38446 40238 38498 40290
rect 41918 40238 41970 40290
rect 51102 40238 51154 40290
rect 52222 40238 52274 40290
rect 57598 40238 57650 40290
rect 60398 40238 60450 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 17054 39790 17106 39842
rect 20862 39790 20914 39842
rect 27470 39790 27522 39842
rect 37774 39790 37826 39842
rect 48414 39790 48466 39842
rect 9102 39678 9154 39730
rect 11902 39678 11954 39730
rect 22206 39678 22258 39730
rect 23102 39678 23154 39730
rect 27918 39678 27970 39730
rect 28590 39678 28642 39730
rect 31166 39678 31218 39730
rect 34750 39678 34802 39730
rect 42702 39678 42754 39730
rect 49198 39678 49250 39730
rect 49646 39678 49698 39730
rect 51438 39678 51490 39730
rect 51774 39678 51826 39730
rect 57038 39678 57090 39730
rect 57934 39678 57986 39730
rect 61518 39678 61570 39730
rect 13470 39566 13522 39618
rect 14030 39566 14082 39618
rect 17166 39566 17218 39618
rect 17726 39566 17778 39618
rect 22430 39566 22482 39618
rect 23998 39566 24050 39618
rect 24334 39566 24386 39618
rect 29150 39566 29202 39618
rect 34974 39566 35026 39618
rect 40910 39566 40962 39618
rect 41246 39566 41298 39618
rect 44942 39566 44994 39618
rect 45390 39566 45442 39618
rect 53006 39566 53058 39618
rect 53678 39566 53730 39618
rect 8094 39454 8146 39506
rect 10782 39454 10834 39506
rect 16270 39454 16322 39506
rect 21310 39454 21362 39506
rect 21646 39454 21698 39506
rect 22878 39454 22930 39506
rect 26686 39454 26738 39506
rect 38558 39454 38610 39506
rect 44046 39454 44098 39506
rect 50878 39454 50930 39506
rect 58942 39454 58994 39506
rect 62526 39454 62578 39506
rect 20190 39342 20242 39394
rect 28478 39342 28530 39394
rect 37438 39342 37490 39394
rect 41806 39342 41858 39394
rect 47854 39342 47906 39394
rect 48750 39342 48802 39394
rect 52782 39342 52834 39394
rect 55918 39342 55970 39394
rect 56702 39342 56754 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 16270 39006 16322 39058
rect 16942 39006 16994 39058
rect 20974 39006 21026 39058
rect 21086 39006 21138 39058
rect 21870 39006 21922 39058
rect 28030 39006 28082 39058
rect 36878 39006 36930 39058
rect 37550 39006 37602 39058
rect 43934 39006 43986 39058
rect 44606 39006 44658 39058
rect 45390 39006 45442 39058
rect 52446 39006 52498 39058
rect 53790 39006 53842 39058
rect 56702 39006 56754 39058
rect 6974 38894 7026 38946
rect 11006 38894 11058 38946
rect 20190 38894 20242 38946
rect 28814 38894 28866 38946
rect 31950 38894 32002 38946
rect 32286 38894 32338 38946
rect 47070 38894 47122 38946
rect 53230 38894 53282 38946
rect 55470 38894 55522 38946
rect 58830 38894 58882 38946
rect 61406 38894 61458 38946
rect 13470 38782 13522 38834
rect 13806 38782 13858 38834
rect 17278 38782 17330 38834
rect 17838 38782 17890 38834
rect 24222 38782 24274 38834
rect 24670 38782 24722 38834
rect 27806 38782 27858 38834
rect 31166 38782 31218 38834
rect 31502 38782 31554 38834
rect 33854 38782 33906 38834
rect 34526 38782 34578 38834
rect 40238 38782 40290 38834
rect 40910 38782 40962 38834
rect 41582 38782 41634 38834
rect 49534 38782 49586 38834
rect 50206 38782 50258 38834
rect 7982 38670 8034 38722
rect 9998 38670 10050 38722
rect 10222 38670 10274 38722
rect 12014 38670 12066 38722
rect 25454 38670 25506 38722
rect 44942 38670 44994 38722
rect 45838 38670 45890 38722
rect 47742 38670 47794 38722
rect 47966 38670 48018 38722
rect 48750 38670 48802 38722
rect 48974 38670 49026 38722
rect 54462 38670 54514 38722
rect 57598 38670 57650 38722
rect 60398 38670 60450 38722
rect 37998 38558 38050 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 27694 38222 27746 38274
rect 35086 38222 35138 38274
rect 42702 38222 42754 38274
rect 7870 38110 7922 38162
rect 15822 38110 15874 38162
rect 22654 38110 22706 38162
rect 28030 38110 28082 38162
rect 37438 38110 37490 38162
rect 37662 38110 37714 38162
rect 38110 38110 38162 38162
rect 43710 38110 43762 38162
rect 56702 38110 56754 38162
rect 61518 38110 61570 38162
rect 9326 37998 9378 38050
rect 9886 37998 9938 38050
rect 15038 37998 15090 38050
rect 20638 37998 20690 38050
rect 23998 37998 24050 38050
rect 24558 37998 24610 38050
rect 31390 37998 31442 38050
rect 31950 37998 32002 38050
rect 39230 37998 39282 38050
rect 39678 37998 39730 38050
rect 43150 37998 43202 38050
rect 43822 37998 43874 38050
rect 44830 37998 44882 38050
rect 45390 37998 45442 38050
rect 48750 37998 48802 38050
rect 49198 37998 49250 38050
rect 52782 37998 52834 38050
rect 7086 37886 7138 37938
rect 19742 37886 19794 37938
rect 20078 37886 20130 37938
rect 20414 37886 20466 37938
rect 21534 37886 21586 37938
rect 26910 37886 26962 37938
rect 30830 37886 30882 37938
rect 31166 37886 31218 37938
rect 38446 37886 38498 37938
rect 42926 37886 42978 37938
rect 62526 37886 62578 37938
rect 12462 37774 12514 37826
rect 13022 37774 13074 37826
rect 23326 37774 23378 37826
rect 34302 37774 34354 37826
rect 42142 37774 42194 37826
rect 47630 37774 47682 37826
rect 48414 37774 48466 37826
rect 51438 37774 51490 37826
rect 52222 37774 52274 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 16382 37438 16434 37490
rect 16942 37438 16994 37490
rect 20190 37438 20242 37490
rect 20974 37438 21026 37490
rect 24222 37438 24274 37490
rect 24782 37438 24834 37490
rect 32622 37438 32674 37490
rect 34302 37438 34354 37490
rect 38558 37438 38610 37490
rect 48190 37438 48242 37490
rect 53118 37438 53170 37490
rect 4174 37326 4226 37378
rect 6974 37326 7026 37378
rect 11006 37326 11058 37378
rect 25230 37326 25282 37378
rect 25566 37326 25618 37378
rect 31838 37326 31890 37378
rect 33406 37326 33458 37378
rect 34190 37326 34242 37378
rect 47294 37326 47346 37378
rect 47630 37326 47682 37378
rect 48750 37326 48802 37378
rect 49534 37326 49586 37378
rect 53902 37326 53954 37378
rect 54910 37326 54962 37378
rect 55806 37326 55858 37378
rect 56702 37326 56754 37378
rect 58830 37326 58882 37378
rect 61406 37326 61458 37378
rect 13246 37214 13298 37266
rect 13918 37214 13970 37266
rect 17278 37214 17330 37266
rect 17950 37214 18002 37266
rect 21310 37214 21362 37266
rect 21646 37214 21698 37266
rect 26126 37214 26178 37266
rect 28926 37214 28978 37266
rect 29486 37214 29538 37266
rect 35646 37214 35698 37266
rect 36318 37214 36370 37266
rect 41806 37214 41858 37266
rect 49982 37214 50034 37266
rect 50654 37214 50706 37266
rect 54238 37214 54290 37266
rect 54686 37214 54738 37266
rect 5182 37102 5234 37154
rect 7982 37102 8034 37154
rect 12014 37102 12066 37154
rect 28030 37102 28082 37154
rect 33070 37102 33122 37154
rect 39678 37102 39730 37154
rect 40126 37102 40178 37154
rect 40350 37102 40402 37154
rect 41358 37102 41410 37154
rect 46734 37102 46786 37154
rect 48974 37102 49026 37154
rect 55470 37102 55522 37154
rect 57598 37102 57650 37154
rect 60398 37102 60450 37154
rect 39342 36990 39394 37042
rect 53678 36990 53730 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 13022 36654 13074 36706
rect 27694 36654 27746 36706
rect 36542 36654 36594 36706
rect 41694 36654 41746 36706
rect 45502 36654 45554 36706
rect 56254 36654 56306 36706
rect 3950 36542 4002 36594
rect 8094 36542 8146 36594
rect 14030 36542 14082 36594
rect 19742 36542 19794 36594
rect 20078 36542 20130 36594
rect 22654 36542 22706 36594
rect 37326 36542 37378 36594
rect 42030 36542 42082 36594
rect 42814 36542 42866 36594
rect 43150 36542 43202 36594
rect 44382 36542 44434 36594
rect 50318 36542 50370 36594
rect 51438 36542 51490 36594
rect 57710 36542 57762 36594
rect 61518 36542 61570 36594
rect 9326 36430 9378 36482
rect 9886 36430 9938 36482
rect 14814 36430 14866 36482
rect 18174 36430 18226 36482
rect 18622 36430 18674 36482
rect 24222 36430 24274 36482
rect 24558 36430 24610 36482
rect 29038 36430 29090 36482
rect 29598 36430 29650 36482
rect 32734 36430 32786 36482
rect 33070 36430 33122 36482
rect 33518 36430 33570 36482
rect 37774 36430 37826 36482
rect 37998 36430 38050 36482
rect 38670 36430 38722 36482
rect 47070 36430 47122 36482
rect 48078 36430 48130 36482
rect 48302 36430 48354 36482
rect 51326 36430 51378 36482
rect 52558 36430 52610 36482
rect 53230 36430 53282 36482
rect 56590 36430 56642 36482
rect 1710 36318 1762 36370
rect 3054 36318 3106 36370
rect 7086 36318 7138 36370
rect 13694 36318 13746 36370
rect 14590 36318 14642 36370
rect 19518 36318 19570 36370
rect 20414 36318 20466 36370
rect 20750 36318 20802 36370
rect 21758 36318 21810 36370
rect 36990 36318 37042 36370
rect 40910 36318 40962 36370
rect 43486 36318 43538 36370
rect 58494 36318 58546 36370
rect 62526 36318 62578 36370
rect 2046 36206 2098 36258
rect 12462 36206 12514 36258
rect 15150 36206 15202 36258
rect 15934 36206 15986 36258
rect 23214 36206 23266 36258
rect 23662 36206 23714 36258
rect 27022 36206 27074 36258
rect 28030 36206 28082 36258
rect 32174 36206 32226 36258
rect 35982 36206 36034 36258
rect 55470 36206 55522 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 1822 35870 1874 35922
rect 11454 35870 11506 35922
rect 11902 35870 11954 35922
rect 12686 35870 12738 35922
rect 19182 35870 19234 35922
rect 19742 35870 19794 35922
rect 28366 35870 28418 35922
rect 29150 35870 29202 35922
rect 37774 35870 37826 35922
rect 38558 35870 38610 35922
rect 38894 35870 38946 35922
rect 43710 35870 43762 35922
rect 44494 35870 44546 35922
rect 47742 35870 47794 35922
rect 48302 35870 48354 35922
rect 48862 35870 48914 35922
rect 49310 35870 49362 35922
rect 53678 35870 53730 35922
rect 56702 35870 56754 35922
rect 4174 35758 4226 35810
rect 6974 35758 7026 35810
rect 15822 35758 15874 35810
rect 16494 35758 16546 35810
rect 17390 35758 17442 35810
rect 18174 35758 18226 35810
rect 23438 35758 23490 35810
rect 33070 35758 33122 35810
rect 33406 35758 33458 35810
rect 34078 35758 34130 35810
rect 50318 35758 50370 35810
rect 55134 35758 55186 35810
rect 58830 35758 58882 35810
rect 61406 35758 61458 35810
rect 15038 35646 15090 35698
rect 15374 35646 15426 35698
rect 16046 35646 16098 35698
rect 16718 35646 16770 35698
rect 17614 35646 17666 35698
rect 22206 35646 22258 35698
rect 22878 35646 22930 35698
rect 26014 35646 26066 35698
rect 31390 35646 31442 35698
rect 31950 35646 32002 35698
rect 34862 35646 34914 35698
rect 35534 35646 35586 35698
rect 41022 35646 41074 35698
rect 41470 35646 41522 35698
rect 44830 35646 44882 35698
rect 45278 35646 45330 35698
rect 50542 35646 50594 35698
rect 51102 35646 51154 35698
rect 54910 35646 54962 35698
rect 55582 35646 55634 35698
rect 5182 35534 5234 35586
rect 7982 35534 8034 35586
rect 11342 35534 11394 35586
rect 18398 35534 18450 35586
rect 18958 35534 19010 35586
rect 24446 35534 24498 35586
rect 27806 35534 27858 35586
rect 32622 35534 32674 35586
rect 33742 35534 33794 35586
rect 49982 35534 50034 35586
rect 55694 35534 55746 35586
rect 57598 35534 57650 35586
rect 60398 35534 60450 35586
rect 54238 35422 54290 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 17054 35086 17106 35138
rect 56366 35086 56418 35138
rect 3838 34974 3890 35026
rect 7310 34974 7362 35026
rect 12910 34974 12962 35026
rect 26350 34974 26402 35026
rect 27022 34974 27074 35026
rect 29934 34974 29986 35026
rect 37102 34974 37154 35026
rect 37326 34974 37378 35026
rect 44270 34974 44322 35026
rect 46734 34974 46786 35026
rect 52110 34974 52162 35026
rect 56814 34974 56866 35026
rect 57598 34974 57650 35026
rect 59390 34974 59442 35026
rect 61518 34974 61570 35026
rect 8766 34862 8818 34914
rect 9102 34862 9154 34914
rect 12238 34862 12290 34914
rect 13470 34862 13522 34914
rect 13918 34862 13970 34914
rect 17166 34862 17218 34914
rect 17726 34862 17778 34914
rect 22766 34862 22818 34914
rect 30158 34862 30210 34914
rect 37886 34862 37938 34914
rect 46062 34862 46114 34914
rect 46958 34862 47010 34914
rect 47630 34862 47682 34914
rect 50990 34862 51042 34914
rect 52670 34862 52722 34914
rect 53342 34862 53394 34914
rect 3054 34750 3106 34802
rect 6302 34750 6354 34802
rect 12574 34750 12626 34802
rect 27246 34750 27298 34802
rect 27582 34750 27634 34802
rect 35198 34750 35250 34802
rect 42926 34750 42978 34802
rect 45166 34750 45218 34802
rect 45502 34750 45554 34802
rect 46286 34750 46338 34802
rect 51214 34750 51266 34802
rect 51774 34750 51826 34802
rect 58830 34750 58882 34802
rect 62526 34750 62578 34802
rect 11678 34638 11730 34690
rect 16494 34638 16546 34690
rect 20190 34638 20242 34690
rect 20862 34638 20914 34690
rect 27694 34638 27746 34690
rect 28366 34638 28418 34690
rect 29262 34638 29314 34690
rect 36542 34638 36594 34690
rect 43598 34638 43650 34690
rect 49982 34638 50034 34690
rect 50654 34638 50706 34690
rect 55694 34638 55746 34690
rect 59502 34638 59554 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 11118 34302 11170 34354
rect 11902 34302 11954 34354
rect 15262 34302 15314 34354
rect 20414 34302 20466 34354
rect 20974 34302 21026 34354
rect 24222 34302 24274 34354
rect 24782 34302 24834 34354
rect 31278 34302 31330 34354
rect 31838 34302 31890 34354
rect 39902 34302 39954 34354
rect 51550 34302 51602 34354
rect 52334 34302 52386 34354
rect 55358 34302 55410 34354
rect 56142 34302 56194 34354
rect 4174 34190 4226 34242
rect 6974 34190 7026 34242
rect 27134 34190 27186 34242
rect 32062 34190 32114 34242
rect 32398 34190 32450 34242
rect 33742 34190 33794 34242
rect 43710 34190 43762 34242
rect 58830 34190 58882 34242
rect 61406 34190 61458 34242
rect 14142 34078 14194 34130
rect 14702 34078 14754 34130
rect 17278 34078 17330 34130
rect 17838 34078 17890 34130
rect 21086 34078 21138 34130
rect 21646 34078 21698 34130
rect 25342 34078 25394 34130
rect 28366 34078 28418 34130
rect 28702 34078 28754 34130
rect 36094 34078 36146 34130
rect 36430 34078 36482 34130
rect 36766 34078 36818 34130
rect 37438 34078 37490 34130
rect 41022 34078 41074 34130
rect 41470 34078 41522 34130
rect 45614 34078 45666 34130
rect 48862 34078 48914 34130
rect 49310 34078 49362 34130
rect 52446 34078 52498 34130
rect 53118 34078 53170 34130
rect 5182 33966 5234 34018
rect 7982 33966 8034 34018
rect 9998 33966 10050 34018
rect 10222 33966 10274 34018
rect 10558 33966 10610 34018
rect 15822 33966 15874 34018
rect 16270 33966 16322 34018
rect 16494 33966 16546 34018
rect 16830 33966 16882 34018
rect 44494 33966 44546 34018
rect 44718 33966 44770 34018
rect 45054 33966 45106 34018
rect 56814 33966 56866 34018
rect 57598 33966 57650 34018
rect 60398 33966 60450 34018
rect 32958 33854 33010 33906
rect 40462 33854 40514 33906
rect 47966 33854 48018 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 9102 33518 9154 33570
rect 15934 33518 15986 33570
rect 4062 33406 4114 33458
rect 7870 33406 7922 33458
rect 13470 33406 13522 33458
rect 13806 33406 13858 33458
rect 21422 33406 21474 33458
rect 22206 33406 22258 33458
rect 34302 33406 34354 33458
rect 35086 33406 35138 33458
rect 35646 33406 35698 33458
rect 42926 33406 42978 33458
rect 43262 33406 43314 33458
rect 43934 33406 43986 33458
rect 52782 33406 52834 33458
rect 53678 33406 53730 33458
rect 56478 33406 56530 33458
rect 61518 33406 61570 33458
rect 12126 33294 12178 33346
rect 12574 33294 12626 33346
rect 16718 33294 16770 33346
rect 17166 33294 17218 33346
rect 17726 33294 17778 33346
rect 22542 33294 22594 33346
rect 22766 33294 22818 33346
rect 28478 33294 28530 33346
rect 30606 33294 30658 33346
rect 30942 33294 30994 33346
rect 34526 33294 34578 33346
rect 36094 33294 36146 33346
rect 38558 33294 38610 33346
rect 44718 33294 44770 33346
rect 45390 33294 45442 33346
rect 48526 33294 48578 33346
rect 49198 33294 49250 33346
rect 3054 33182 3106 33234
rect 6638 33182 6690 33234
rect 9886 33182 9938 33234
rect 21646 33182 21698 33234
rect 23550 33182 23602 33234
rect 29822 33182 29874 33234
rect 30158 33182 30210 33234
rect 35870 33182 35922 33234
rect 40350 33182 40402 33234
rect 47630 33182 47682 33234
rect 54686 33182 54738 33234
rect 57486 33182 57538 33234
rect 62526 33182 62578 33234
rect 8878 33070 8930 33122
rect 20302 33070 20354 33122
rect 20862 33070 20914 33122
rect 33518 33070 33570 33122
rect 34078 33070 34130 33122
rect 43822 33070 43874 33122
rect 48414 33070 48466 33122
rect 51662 33070 51714 33122
rect 52222 33070 52274 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 16158 32734 16210 32786
rect 29486 32734 29538 32786
rect 39902 32734 39954 32786
rect 41134 32734 41186 32786
rect 44382 32734 44434 32786
rect 44942 32734 44994 32786
rect 4174 32622 4226 32674
rect 6974 32622 7026 32674
rect 15374 32622 15426 32674
rect 24334 32622 24386 32674
rect 27246 32622 27298 32674
rect 33742 32622 33794 32674
rect 47182 32622 47234 32674
rect 50766 32622 50818 32674
rect 53790 32622 53842 32674
rect 58830 32622 58882 32674
rect 61406 32622 61458 32674
rect 9102 32510 9154 32562
rect 9886 32510 9938 32562
rect 12574 32510 12626 32562
rect 13022 32510 13074 32562
rect 18398 32510 18450 32562
rect 23774 32510 23826 32562
rect 25902 32510 25954 32562
rect 28478 32510 28530 32562
rect 31838 32510 31890 32562
rect 32398 32510 32450 32562
rect 36094 32510 36146 32562
rect 36542 32510 36594 32562
rect 36766 32510 36818 32562
rect 37438 32510 37490 32562
rect 41246 32510 41298 32562
rect 41918 32510 41970 32562
rect 45390 32510 45442 32562
rect 48078 32510 48130 32562
rect 54574 32510 54626 32562
rect 5182 32398 5234 32450
rect 7982 32398 8034 32450
rect 16494 32398 16546 32450
rect 16830 32398 16882 32450
rect 19518 32398 19570 32450
rect 22990 32398 23042 32450
rect 23326 32398 23378 32450
rect 23886 32398 23938 32450
rect 24670 32398 24722 32450
rect 45726 32398 45778 32450
rect 46174 32398 46226 32450
rect 48862 32398 48914 32450
rect 49310 32398 49362 32450
rect 49758 32398 49810 32450
rect 52222 32398 52274 32450
rect 52558 32398 52610 32450
rect 54462 32398 54514 32450
rect 57598 32398 57650 32450
rect 60398 32398 60450 32450
rect 10670 32286 10722 32338
rect 28702 32286 28754 32338
rect 32958 32286 33010 32338
rect 40462 32286 40514 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 4062 31838 4114 31890
rect 7870 31838 7922 31890
rect 9102 31838 9154 31890
rect 13022 31838 13074 31890
rect 17054 31838 17106 31890
rect 21198 31838 21250 31890
rect 36990 31838 37042 31890
rect 42926 31838 42978 31890
rect 43262 31838 43314 31890
rect 49646 31838 49698 31890
rect 51438 31838 51490 31890
rect 57486 31838 57538 31890
rect 61518 31838 61570 31890
rect 64318 31838 64370 31890
rect 9438 31726 9490 31778
rect 9886 31726 9938 31778
rect 13358 31726 13410 31778
rect 13918 31726 13970 31778
rect 17166 31726 17218 31778
rect 17726 31726 17778 31778
rect 24222 31726 24274 31778
rect 24670 31726 24722 31778
rect 28142 31726 28194 31778
rect 28590 31726 28642 31778
rect 29262 31726 29314 31778
rect 29710 31726 29762 31778
rect 32958 31726 33010 31778
rect 33406 31726 33458 31778
rect 36542 31726 36594 31778
rect 38222 31726 38274 31778
rect 38670 31726 38722 31778
rect 42254 31726 42306 31778
rect 42702 31726 42754 31778
rect 44158 31726 44210 31778
rect 44718 31726 44770 31778
rect 45390 31726 45442 31778
rect 52782 31726 52834 31778
rect 53230 31726 53282 31778
rect 3054 31614 3106 31666
rect 7086 31614 7138 31666
rect 20078 31614 20130 31666
rect 20862 31614 20914 31666
rect 21982 31614 22034 31666
rect 25790 31614 25842 31666
rect 37326 31614 37378 31666
rect 41694 31614 41746 31666
rect 41918 31614 41970 31666
rect 43934 31614 43986 31666
rect 50878 31614 50930 31666
rect 58494 31614 58546 31666
rect 62526 31614 62578 31666
rect 65550 31614 65602 31666
rect 8654 31502 8706 31554
rect 12350 31502 12402 31554
rect 16494 31502 16546 31554
rect 25006 31502 25058 31554
rect 32062 31502 32114 31554
rect 32734 31502 32786 31554
rect 35870 31502 35922 31554
rect 37774 31502 37826 31554
rect 41134 31502 41186 31554
rect 43374 31502 43426 31554
rect 47854 31502 47906 31554
rect 48414 31502 48466 31554
rect 48750 31502 48802 31554
rect 49198 31502 49250 31554
rect 51550 31502 51602 31554
rect 55694 31502 55746 31554
rect 56254 31502 56306 31554
rect 56590 31502 56642 31554
rect 57038 31502 57090 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 8878 31166 8930 31218
rect 12462 31166 12514 31218
rect 13134 31166 13186 31218
rect 16382 31166 16434 31218
rect 17838 31166 17890 31218
rect 22542 31166 22594 31218
rect 23998 31166 24050 31218
rect 25454 31166 25506 31218
rect 36094 31166 36146 31218
rect 39902 31166 39954 31218
rect 43710 31166 43762 31218
rect 47742 31166 47794 31218
rect 48302 31166 48354 31218
rect 56142 31166 56194 31218
rect 59502 31166 59554 31218
rect 60510 31166 60562 31218
rect 2158 31054 2210 31106
rect 5182 31054 5234 31106
rect 8990 31054 9042 31106
rect 16942 31054 16994 31106
rect 17726 31054 17778 31106
rect 26686 31054 26738 31106
rect 51550 31054 51602 31106
rect 55358 31054 55410 31106
rect 62414 31054 62466 31106
rect 7534 30942 7586 30994
rect 7982 30942 8034 30994
rect 9438 30942 9490 30994
rect 10110 30942 10162 30994
rect 13246 30942 13298 30994
rect 13806 30942 13858 30994
rect 19518 30942 19570 30994
rect 20190 30942 20242 30994
rect 27134 30942 27186 30994
rect 32958 30942 33010 30994
rect 33630 30942 33682 30994
rect 37326 30942 37378 30994
rect 39790 30942 39842 30994
rect 41022 30942 41074 30994
rect 41470 30942 41522 30994
rect 44718 30942 44770 30994
rect 45166 30942 45218 30994
rect 48750 30942 48802 30994
rect 49310 30942 49362 30994
rect 52670 30942 52722 30994
rect 53118 30942 53170 30994
rect 56478 30942 56530 30994
rect 57150 30942 57202 30994
rect 60174 30942 60226 30994
rect 64990 30942 65042 30994
rect 66110 30942 66162 30994
rect 3166 30830 3218 30882
rect 18510 30830 18562 30882
rect 19294 30830 19346 30882
rect 23550 30830 23602 30882
rect 26014 30830 26066 30882
rect 26350 30830 26402 30882
rect 32174 30830 32226 30882
rect 61406 30830 61458 30882
rect 4398 30718 4450 30770
rect 23214 30718 23266 30770
rect 36654 30718 36706 30770
rect 38334 30718 38386 30770
rect 44494 30718 44546 30770
rect 52334 30718 52386 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 4062 30270 4114 30322
rect 7086 30270 7138 30322
rect 12462 30270 12514 30322
rect 14702 30270 14754 30322
rect 15038 30270 15090 30322
rect 19630 30270 19682 30322
rect 21422 30270 21474 30322
rect 22542 30270 22594 30322
rect 50766 30270 50818 30322
rect 55470 30270 55522 30322
rect 61518 30270 61570 30322
rect 4510 30158 4562 30210
rect 8318 30158 8370 30210
rect 11342 30158 11394 30210
rect 12014 30158 12066 30210
rect 13694 30158 13746 30210
rect 14030 30158 14082 30210
rect 15374 30158 15426 30210
rect 18622 30158 18674 30210
rect 19070 30158 19122 30210
rect 20302 30158 20354 30210
rect 20750 30158 20802 30210
rect 21646 30158 21698 30210
rect 22318 30158 22370 30210
rect 26686 30158 26738 30210
rect 27246 30158 27298 30210
rect 27470 30158 27522 30210
rect 28254 30158 28306 30210
rect 29262 30158 29314 30210
rect 29598 30158 29650 30210
rect 32958 30158 33010 30210
rect 33518 30158 33570 30210
rect 37102 30158 37154 30210
rect 37550 30158 37602 30210
rect 40686 30158 40738 30210
rect 41246 30158 41298 30210
rect 46286 30158 46338 30210
rect 53902 30158 53954 30210
rect 3054 30046 3106 30098
rect 6078 30046 6130 30098
rect 12238 30046 12290 30098
rect 16382 30046 16434 30098
rect 24334 30046 24386 30098
rect 46846 30046 46898 30098
rect 50430 30046 50482 30098
rect 51662 30046 51714 30098
rect 51998 30046 52050 30098
rect 52782 30046 52834 30098
rect 53118 30046 53170 30098
rect 62526 30046 62578 30098
rect 7646 29934 7698 29986
rect 8094 29934 8146 29986
rect 8878 29934 8930 29986
rect 15598 29934 15650 29986
rect 23550 29934 23602 29986
rect 27582 29934 27634 29986
rect 32174 29934 32226 29986
rect 32734 29934 32786 29986
rect 35982 29934 36034 29986
rect 36542 29934 36594 29986
rect 40014 29934 40066 29986
rect 40574 29934 40626 29986
rect 43598 29934 43650 29986
rect 44382 29934 44434 29986
rect 51214 29934 51266 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 12574 29598 12626 29650
rect 13246 29598 13298 29650
rect 17502 29598 17554 29650
rect 17950 29598 18002 29650
rect 20302 29598 20354 29650
rect 20862 29598 20914 29650
rect 23998 29598 24050 29650
rect 28142 29598 28194 29650
rect 45278 29598 45330 29650
rect 46286 29598 46338 29650
rect 46734 29598 46786 29650
rect 47182 29598 47234 29650
rect 51662 29598 51714 29650
rect 53118 29598 53170 29650
rect 56702 29598 56754 29650
rect 57150 29598 57202 29650
rect 3166 29486 3218 29538
rect 6190 29486 6242 29538
rect 14030 29486 14082 29538
rect 18846 29486 18898 29538
rect 29710 29486 29762 29538
rect 33070 29486 33122 29538
rect 33742 29486 33794 29538
rect 40910 29486 40962 29538
rect 41246 29486 41298 29538
rect 41918 29486 41970 29538
rect 58830 29486 58882 29538
rect 61406 29486 61458 29538
rect 8430 29374 8482 29426
rect 9102 29374 9154 29426
rect 9662 29374 9714 29426
rect 10110 29374 10162 29426
rect 16382 29374 16434 29426
rect 16830 29374 16882 29426
rect 21310 29374 21362 29426
rect 21646 29374 21698 29426
rect 25342 29374 25394 29426
rect 25790 29374 25842 29426
rect 32062 29374 32114 29426
rect 32622 29374 32674 29426
rect 33966 29374 34018 29426
rect 36206 29374 36258 29426
rect 42254 29374 42306 29426
rect 42926 29374 42978 29426
rect 48862 29374 48914 29426
rect 49310 29374 49362 29426
rect 55582 29374 55634 29426
rect 55918 29374 55970 29426
rect 4174 29262 4226 29314
rect 19854 29262 19906 29314
rect 33406 29262 33458 29314
rect 38558 29262 38610 29314
rect 41582 29262 41634 29314
rect 47966 29262 48018 29314
rect 48190 29262 48242 29314
rect 57598 29262 57650 29314
rect 60398 29262 60450 29314
rect 5406 29150 5458 29202
rect 13134 29150 13186 29202
rect 24782 29150 24834 29202
rect 28814 29150 28866 29202
rect 28926 29150 28978 29202
rect 45950 29150 46002 29202
rect 52334 29150 52386 29202
rect 52446 29150 52498 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 25790 28814 25842 28866
rect 48526 28814 48578 28866
rect 4062 28702 4114 28754
rect 4510 28702 4562 28754
rect 6862 28702 6914 28754
rect 7870 28702 7922 28754
rect 12238 28702 12290 28754
rect 12686 28702 12738 28754
rect 12910 28702 12962 28754
rect 15710 28702 15762 28754
rect 16382 28702 16434 28754
rect 28366 28702 28418 28754
rect 29262 28702 29314 28754
rect 30494 28702 30546 28754
rect 30718 28702 30770 28754
rect 36094 28702 36146 28754
rect 51102 28702 51154 28754
rect 51662 28702 51714 28754
rect 51998 28702 52050 28754
rect 56590 28702 56642 28754
rect 57486 28702 57538 28754
rect 59502 28702 59554 28754
rect 61518 28702 61570 28754
rect 6526 28590 6578 28642
rect 7198 28590 7250 28642
rect 7646 28590 7698 28642
rect 11118 28590 11170 28642
rect 11566 28590 11618 28642
rect 13806 28590 13858 28642
rect 17166 28590 17218 28642
rect 17726 28590 17778 28642
rect 21534 28590 21586 28642
rect 22318 28590 22370 28642
rect 22654 28590 22706 28642
rect 26014 28590 26066 28642
rect 29710 28590 29762 28642
rect 29934 28590 29986 28642
rect 34078 28590 34130 28642
rect 34638 28590 34690 28642
rect 35086 28590 35138 28642
rect 36318 28590 36370 28642
rect 36878 28590 36930 28642
rect 40014 28590 40066 28642
rect 40574 28590 40626 28642
rect 43710 28590 43762 28642
rect 44158 28590 44210 28642
rect 44830 28590 44882 28642
rect 45502 28590 45554 28642
rect 48750 28590 48802 28642
rect 52670 28590 52722 28642
rect 53230 28590 53282 28642
rect 59278 28590 59330 28642
rect 3054 28478 3106 28530
rect 8878 28478 8930 28530
rect 34862 28478 34914 28530
rect 41470 28478 41522 28530
rect 58494 28478 58546 28530
rect 62526 28478 62578 28530
rect 6414 28366 6466 28418
rect 8094 28366 8146 28418
rect 16494 28366 16546 28418
rect 20302 28366 20354 28418
rect 20862 28366 20914 28418
rect 21310 28366 21362 28418
rect 25118 28366 25170 28418
rect 30942 28366 30994 28418
rect 31726 28366 31778 28418
rect 37662 28366 37714 28418
rect 40686 28366 40738 28418
rect 47854 28366 47906 28418
rect 55582 28366 55634 28418
rect 56254 28366 56306 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 4734 28030 4786 28082
rect 16830 28030 16882 28082
rect 17950 28030 18002 28082
rect 19294 28030 19346 28082
rect 20750 28030 20802 28082
rect 26238 28030 26290 28082
rect 26686 28030 26738 28082
rect 27246 28030 27298 28082
rect 28254 28030 28306 28082
rect 33182 28030 33234 28082
rect 37326 28030 37378 28082
rect 38894 28030 38946 28082
rect 39454 28030 39506 28082
rect 41582 28030 41634 28082
rect 47742 28030 47794 28082
rect 48862 28030 48914 28082
rect 53118 28030 53170 28082
rect 56702 28030 56754 28082
rect 8318 27918 8370 27970
rect 10558 27918 10610 27970
rect 12686 27918 12738 27970
rect 24222 27918 24274 27970
rect 31502 27918 31554 27970
rect 33630 27918 33682 27970
rect 38110 27918 38162 27970
rect 39902 27918 39954 27970
rect 40238 27918 40290 27970
rect 54574 27918 54626 27970
rect 54910 27918 54962 27970
rect 55246 27918 55298 27970
rect 55694 27918 55746 27970
rect 56030 27918 56082 27970
rect 58942 27918 58994 27970
rect 61406 27918 61458 27970
rect 1822 27806 1874 27858
rect 2270 27806 2322 27858
rect 5406 27806 5458 27858
rect 5966 27806 6018 27858
rect 9886 27806 9938 27858
rect 10894 27806 10946 27858
rect 11454 27806 11506 27858
rect 14926 27806 14978 27858
rect 15598 27806 15650 27858
rect 18174 27806 18226 27858
rect 22990 27806 23042 27858
rect 23662 27806 23714 27858
rect 25230 27806 25282 27858
rect 30606 27806 30658 27858
rect 31166 27806 31218 27858
rect 32398 27806 32450 27858
rect 33854 27806 33906 27858
rect 34414 27806 34466 27858
rect 34750 27806 34802 27858
rect 38334 27806 38386 27858
rect 43934 27806 43986 27858
rect 44270 27806 44322 27858
rect 44830 27806 44882 27858
rect 45278 27806 45330 27858
rect 49982 27806 50034 27858
rect 50654 27806 50706 27858
rect 54350 27806 54402 27858
rect 9550 27694 9602 27746
rect 11678 27694 11730 27746
rect 15934 27694 15986 27746
rect 16382 27694 16434 27746
rect 17614 27694 17666 27746
rect 19742 27694 19794 27746
rect 23886 27694 23938 27746
rect 24670 27694 24722 27746
rect 31838 27694 31890 27746
rect 32174 27694 32226 27746
rect 39566 27694 39618 27746
rect 49198 27694 49250 27746
rect 49534 27694 49586 27746
rect 57598 27694 57650 27746
rect 60398 27694 60450 27746
rect 5294 27582 5346 27634
rect 9102 27582 9154 27634
rect 11902 27582 11954 27634
rect 15934 27582 15986 27634
rect 16718 27582 16770 27634
rect 19966 27582 20018 27634
rect 25790 27582 25842 27634
rect 26238 27582 26290 27634
rect 27022 27582 27074 27634
rect 27470 27582 27522 27634
rect 37886 27582 37938 27634
rect 40798 27582 40850 27634
rect 48302 27582 48354 27634
rect 53678 27582 53730 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 21310 27246 21362 27298
rect 56254 27246 56306 27298
rect 3950 27134 4002 27186
rect 12798 27134 12850 27186
rect 13694 27134 13746 27186
rect 15374 27134 15426 27186
rect 27022 27134 27074 27186
rect 28254 27134 28306 27186
rect 28590 27134 28642 27186
rect 33966 27134 34018 27186
rect 35758 27134 35810 27186
rect 49758 27134 49810 27186
rect 51550 27134 51602 27186
rect 51886 27134 51938 27186
rect 57486 27134 57538 27186
rect 59278 27134 59330 27186
rect 61518 27134 61570 27186
rect 11678 27022 11730 27074
rect 13918 27022 13970 27074
rect 14814 27022 14866 27074
rect 17390 27022 17442 27074
rect 17726 27022 17778 27074
rect 21534 27022 21586 27074
rect 22430 27022 22482 27074
rect 23214 27022 23266 27074
rect 23662 27022 23714 27074
rect 29262 27022 29314 27074
rect 29710 27022 29762 27074
rect 37102 27022 37154 27074
rect 37550 27022 37602 27074
rect 40686 27022 40738 27074
rect 41358 27022 41410 27074
rect 44718 27022 44770 27074
rect 45390 27022 45442 27074
rect 50766 27022 50818 27074
rect 52782 27022 52834 27074
rect 53230 27022 53282 27074
rect 59502 27022 59554 27074
rect 3054 26910 3106 26962
rect 5742 26910 5794 26962
rect 7198 26910 7250 26962
rect 20078 26910 20130 26962
rect 25902 26910 25954 26962
rect 27470 26910 27522 26962
rect 27918 26910 27970 26962
rect 31950 26910 32002 26962
rect 34974 26910 35026 26962
rect 36094 26910 36146 26962
rect 39790 26910 39842 26962
rect 58494 26910 58546 26962
rect 62526 26910 62578 26962
rect 20862 26798 20914 26850
rect 22206 26798 22258 26850
rect 26686 26798 26738 26850
rect 32734 26798 32786 26850
rect 40574 26798 40626 26850
rect 43822 26798 43874 26850
rect 44382 26798 44434 26850
rect 47854 26798 47906 26850
rect 48414 26798 48466 26850
rect 55470 26798 55522 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 7422 26462 7474 26514
rect 15038 26462 15090 26514
rect 28254 26462 28306 26514
rect 32062 26462 32114 26514
rect 33742 26462 33794 26514
rect 41022 26462 41074 26514
rect 44494 26462 44546 26514
rect 45054 26462 45106 26514
rect 51774 26462 51826 26514
rect 52782 26462 52834 26514
rect 53118 26462 53170 26514
rect 55470 26462 55522 26514
rect 2046 26350 2098 26402
rect 8430 26350 8482 26402
rect 8766 26350 8818 26402
rect 18062 26350 18114 26402
rect 23998 26350 24050 26402
rect 39678 26350 39730 26402
rect 54574 26350 54626 26402
rect 58830 26350 58882 26402
rect 61406 26350 61458 26402
rect 4510 26238 4562 26290
rect 5070 26238 5122 26290
rect 9774 26238 9826 26290
rect 10894 26238 10946 26290
rect 12126 26238 12178 26290
rect 12686 26238 12738 26290
rect 20414 26238 20466 26290
rect 20862 26238 20914 26290
rect 21086 26238 21138 26290
rect 21646 26238 21698 26290
rect 25118 26238 25170 26290
rect 25678 26238 25730 26290
rect 29150 26238 29202 26290
rect 29598 26238 29650 26290
rect 36094 26238 36146 26290
rect 36430 26238 36482 26290
rect 36766 26238 36818 26290
rect 37438 26238 37490 26290
rect 41358 26238 41410 26290
rect 42030 26238 42082 26290
rect 45390 26238 45442 26290
rect 48862 26238 48914 26290
rect 49310 26238 49362 26290
rect 3278 26126 3330 26178
rect 9550 26126 9602 26178
rect 10334 26126 10386 26178
rect 10670 26126 10722 26178
rect 11454 26126 11506 26178
rect 11902 26126 11954 26178
rect 16382 26126 16434 26178
rect 16830 26126 16882 26178
rect 46958 26126 47010 26178
rect 53566 26126 53618 26178
rect 55358 26126 55410 26178
rect 57598 26126 57650 26178
rect 60398 26126 60450 26178
rect 8206 26014 8258 26066
rect 15822 26014 15874 26066
rect 17278 26014 17330 26066
rect 24782 26014 24834 26066
rect 28814 26014 28866 26066
rect 32622 26014 32674 26066
rect 32958 26014 33010 26066
rect 40462 26014 40514 26066
rect 52334 26014 52386 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 19406 25678 19458 25730
rect 4062 25566 4114 25618
rect 5966 25566 6018 25618
rect 7758 25566 7810 25618
rect 8318 25566 8370 25618
rect 8766 25566 8818 25618
rect 13582 25566 13634 25618
rect 14702 25566 14754 25618
rect 21758 25566 21810 25618
rect 23550 25566 23602 25618
rect 24110 25566 24162 25618
rect 29486 25566 29538 25618
rect 30494 25566 30546 25618
rect 42702 25566 42754 25618
rect 43374 25566 43426 25618
rect 43822 25566 43874 25618
rect 44046 25566 44098 25618
rect 44942 25566 44994 25618
rect 51550 25566 51602 25618
rect 57710 25566 57762 25618
rect 59502 25566 59554 25618
rect 8990 25454 9042 25506
rect 9550 25454 9602 25506
rect 15710 25454 15762 25506
rect 16158 25454 16210 25506
rect 19630 25454 19682 25506
rect 20638 25454 20690 25506
rect 24782 25454 24834 25506
rect 25342 25454 25394 25506
rect 31390 25454 31442 25506
rect 32062 25454 32114 25506
rect 38110 25454 38162 25506
rect 38446 25454 38498 25506
rect 39006 25454 39058 25506
rect 43150 25454 43202 25506
rect 45278 25454 45330 25506
rect 45950 25454 46002 25506
rect 48974 25454 49026 25506
rect 49198 25454 49250 25506
rect 52894 25454 52946 25506
rect 53454 25454 53506 25506
rect 1710 25342 1762 25394
rect 2942 25342 2994 25394
rect 6638 25342 6690 25394
rect 14926 25342 14978 25394
rect 15262 25342 15314 25394
rect 19182 25342 19234 25394
rect 21422 25342 21474 25394
rect 22542 25342 22594 25394
rect 37886 25342 37938 25394
rect 42366 25342 42418 25394
rect 48190 25342 48242 25394
rect 58830 25342 58882 25394
rect 2046 25230 2098 25282
rect 5854 25230 5906 25282
rect 12014 25230 12066 25282
rect 12686 25230 12738 25282
rect 18398 25230 18450 25282
rect 20638 25230 20690 25282
rect 24558 25230 24610 25282
rect 27918 25230 27970 25282
rect 28478 25230 28530 25282
rect 29374 25230 29426 25282
rect 30382 25230 30434 25282
rect 30942 25230 30994 25282
rect 34526 25230 34578 25282
rect 35086 25230 35138 25282
rect 41582 25230 41634 25282
rect 42142 25230 42194 25282
rect 55918 25230 55970 25282
rect 56478 25230 56530 25282
rect 59614 25230 59666 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4734 24894 4786 24946
rect 8318 24894 8370 24946
rect 16382 24894 16434 24946
rect 19182 24894 19234 24946
rect 20638 24894 20690 24946
rect 39678 24894 39730 24946
rect 43934 24894 43986 24946
rect 47742 24894 47794 24946
rect 50206 24894 50258 24946
rect 54350 24894 54402 24946
rect 12350 24782 12402 24834
rect 19630 24782 19682 24834
rect 30046 24782 30098 24834
rect 34078 24782 34130 24834
rect 39566 24782 39618 24834
rect 48750 24782 48802 24834
rect 49086 24782 49138 24834
rect 49758 24782 49810 24834
rect 50094 24782 50146 24834
rect 50878 24782 50930 24834
rect 55134 24782 55186 24834
rect 58830 24782 58882 24834
rect 61406 24782 61458 24834
rect 1822 24670 1874 24722
rect 2158 24670 2210 24722
rect 5406 24670 5458 24722
rect 5966 24670 6018 24722
rect 9438 24670 9490 24722
rect 10110 24670 10162 24722
rect 13358 24670 13410 24722
rect 13806 24670 13858 24722
rect 17614 24670 17666 24722
rect 17950 24670 18002 24722
rect 22878 24670 22930 24722
rect 23326 24670 23378 24722
rect 24670 24670 24722 24722
rect 25230 24670 25282 24722
rect 30942 24670 30994 24722
rect 39118 24670 39170 24722
rect 41022 24670 41074 24722
rect 41358 24670 41410 24722
rect 44830 24670 44882 24722
rect 45278 24670 45330 24722
rect 51214 24670 51266 24722
rect 51886 24670 51938 24722
rect 18398 24558 18450 24610
rect 40350 24558 40402 24610
rect 49422 24558 49474 24610
rect 55470 24558 55522 24610
rect 57598 24558 57650 24610
rect 60398 24558 60450 24610
rect 5294 24446 5346 24498
rect 9102 24446 9154 24498
rect 13134 24446 13186 24498
rect 16942 24446 16994 24498
rect 19854 24446 19906 24498
rect 24110 24446 24162 24498
rect 44494 24446 44546 24498
rect 48302 24446 48354 24498
rect 54910 24446 54962 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 1822 23998 1874 24050
rect 3838 23998 3890 24050
rect 5070 23998 5122 24050
rect 5854 23998 5906 24050
rect 6190 23998 6242 24050
rect 6526 23998 6578 24050
rect 11454 23998 11506 24050
rect 12238 23998 12290 24050
rect 19070 23998 19122 24050
rect 19966 23998 20018 24050
rect 20302 23998 20354 24050
rect 20750 23998 20802 24050
rect 29150 23998 29202 24050
rect 29486 23998 29538 24050
rect 45054 23998 45106 24050
rect 49310 23998 49362 24050
rect 49646 23998 49698 24050
rect 50094 23998 50146 24050
rect 51998 23998 52050 24050
rect 52894 23998 52946 24050
rect 58606 23998 58658 24050
rect 9774 23886 9826 23938
rect 10222 23886 10274 23938
rect 10894 23886 10946 23938
rect 11902 23886 11954 23938
rect 12910 23886 12962 23938
rect 17278 23886 17330 23938
rect 19294 23886 19346 23938
rect 21198 23886 21250 23938
rect 21758 23886 21810 23938
rect 25006 23886 25058 23938
rect 25678 23886 25730 23938
rect 34638 23886 34690 23938
rect 35086 23886 35138 23938
rect 35758 23886 35810 23938
rect 37102 23886 37154 23938
rect 37438 23886 37490 23938
rect 40686 23886 40738 23938
rect 41246 23886 41298 23938
rect 45278 23886 45330 23938
rect 45838 23886 45890 23938
rect 56478 23886 56530 23938
rect 3054 23774 3106 23826
rect 6750 23774 6802 23826
rect 7534 23774 7586 23826
rect 10670 23774 10722 23826
rect 12574 23774 12626 23826
rect 13694 23774 13746 23826
rect 24110 23774 24162 23826
rect 30606 23774 30658 23826
rect 35534 23774 35586 23826
rect 51102 23774 51154 23826
rect 58270 23774 58322 23826
rect 24894 23662 24946 23714
rect 28142 23662 28194 23714
rect 28702 23662 28754 23714
rect 29934 23662 29986 23714
rect 30718 23662 30770 23714
rect 31614 23662 31666 23714
rect 32398 23662 32450 23714
rect 39790 23662 39842 23714
rect 40574 23662 40626 23714
rect 43822 23662 43874 23714
rect 44382 23662 44434 23714
rect 48078 23662 48130 23714
rect 48862 23662 48914 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 8318 23326 8370 23378
rect 10222 23326 10274 23378
rect 14030 23326 14082 23378
rect 21870 23326 21922 23378
rect 28254 23326 28306 23378
rect 32062 23326 32114 23378
rect 37438 23326 37490 23378
rect 40350 23326 40402 23378
rect 47854 23326 47906 23378
rect 51662 23326 51714 23378
rect 2830 23214 2882 23266
rect 18062 23214 18114 23266
rect 33070 23214 33122 23266
rect 33742 23214 33794 23266
rect 39230 23214 39282 23266
rect 47966 23214 48018 23266
rect 55358 23214 55410 23266
rect 58830 23214 58882 23266
rect 5406 23102 5458 23154
rect 5966 23102 6018 23154
rect 12574 23102 12626 23154
rect 12910 23102 12962 23154
rect 16270 23102 16322 23154
rect 16830 23102 16882 23154
rect 20302 23102 20354 23154
rect 20750 23102 20802 23154
rect 24222 23102 24274 23154
rect 24782 23102 24834 23154
rect 25118 23102 25170 23154
rect 25678 23102 25730 23154
rect 29150 23102 29202 23154
rect 29598 23102 29650 23154
rect 33294 23102 33346 23154
rect 33966 23102 34018 23154
rect 34302 23102 34354 23154
rect 34974 23102 35026 23154
rect 38446 23102 38498 23154
rect 38894 23102 38946 23154
rect 39566 23102 39618 23154
rect 41694 23102 41746 23154
rect 42030 23102 42082 23154
rect 48862 23102 48914 23154
rect 49310 23102 49362 23154
rect 52446 23102 52498 23154
rect 53006 23102 53058 23154
rect 59502 23102 59554 23154
rect 3950 22990 4002 23042
rect 38222 22990 38274 23042
rect 39790 22990 39842 23042
rect 41022 22990 41074 23042
rect 46958 22990 47010 23042
rect 57598 22990 57650 23042
rect 59614 22990 59666 23042
rect 9102 22878 9154 22930
rect 9438 22878 9490 22930
rect 13246 22878 13298 22930
rect 17278 22878 17330 22930
rect 21086 22878 21138 22930
rect 28814 22878 28866 22930
rect 32622 22878 32674 22930
rect 37998 22878 38050 22930
rect 52334 22878 52386 22930
rect 56142 22878 56194 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 27022 22542 27074 22594
rect 27358 22542 27410 22594
rect 56254 22542 56306 22594
rect 4062 22430 4114 22482
rect 27022 22430 27074 22482
rect 27470 22430 27522 22482
rect 27918 22430 27970 22482
rect 28254 22430 28306 22482
rect 57486 22430 57538 22482
rect 5518 22318 5570 22370
rect 6190 22318 6242 22370
rect 9326 22318 9378 22370
rect 9998 22318 10050 22370
rect 13582 22318 13634 22370
rect 13918 22318 13970 22370
rect 17166 22318 17218 22370
rect 17838 22318 17890 22370
rect 22766 22318 22818 22370
rect 29150 22318 29202 22370
rect 33070 22318 33122 22370
rect 33406 22318 33458 22370
rect 40014 22318 40066 22370
rect 40350 22318 40402 22370
rect 40910 22318 40962 22370
rect 41358 22318 41410 22370
rect 44830 22318 44882 22370
rect 45390 22318 45442 22370
rect 48638 22318 48690 22370
rect 49086 22318 49138 22370
rect 52558 22318 52610 22370
rect 53230 22318 53282 22370
rect 2718 22206 2770 22258
rect 23550 22206 23602 22258
rect 28590 22206 28642 22258
rect 37662 22206 37714 22258
rect 48414 22206 48466 22258
rect 58494 22206 58546 22258
rect 8654 22094 8706 22146
rect 9214 22094 9266 22146
rect 12462 22094 12514 22146
rect 13022 22094 13074 22146
rect 16494 22094 16546 22146
rect 17054 22094 17106 22146
rect 20190 22094 20242 22146
rect 20862 22094 20914 22146
rect 30158 22094 30210 22146
rect 35982 22094 36034 22146
rect 36542 22094 36594 22146
rect 36878 22094 36930 22146
rect 43598 22094 43650 22146
rect 44382 22094 44434 22146
rect 47630 22094 47682 22146
rect 51438 22094 51490 22146
rect 52222 22094 52274 22146
rect 55694 22094 55746 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 10222 21758 10274 21810
rect 20974 21758 21026 21810
rect 25342 21758 25394 21810
rect 26910 21758 26962 21810
rect 30718 21758 30770 21810
rect 36542 21758 36594 21810
rect 42366 21758 42418 21810
rect 45614 21758 45666 21810
rect 46062 21758 46114 21810
rect 51774 21758 51826 21810
rect 53006 21758 53058 21810
rect 3166 21646 3218 21698
rect 8318 21646 8370 21698
rect 16158 21646 16210 21698
rect 35198 21646 35250 21698
rect 47742 21646 47794 21698
rect 54798 21646 54850 21698
rect 55582 21646 55634 21698
rect 55918 21646 55970 21698
rect 58830 21646 58882 21698
rect 5630 21534 5682 21586
rect 5966 21534 6018 21586
rect 12462 21534 12514 21586
rect 12910 21534 12962 21586
rect 13246 21534 13298 21586
rect 13918 21534 13970 21586
rect 17390 21534 17442 21586
rect 23438 21534 23490 21586
rect 23886 21534 23938 21586
rect 25790 21534 25842 21586
rect 27582 21534 27634 21586
rect 27806 21534 27858 21586
rect 28478 21534 28530 21586
rect 38894 21534 38946 21586
rect 39454 21534 39506 21586
rect 39790 21534 39842 21586
rect 44718 21534 44770 21586
rect 45278 21534 45330 21586
rect 48862 21534 48914 21586
rect 49534 21534 49586 21586
rect 4174 21422 4226 21474
rect 24446 21422 24498 21474
rect 25902 21422 25954 21474
rect 34078 21422 34130 21474
rect 41022 21422 41074 21474
rect 46510 21422 46562 21474
rect 53790 21422 53842 21474
rect 57598 21422 57650 21474
rect 9102 21310 9154 21362
rect 9438 21310 9490 21362
rect 16942 21310 16994 21362
rect 19294 21310 19346 21362
rect 20414 21310 20466 21362
rect 24446 21310 24498 21362
rect 24670 21310 24722 21362
rect 31502 21310 31554 21362
rect 35758 21310 35810 21362
rect 41582 21310 41634 21362
rect 52558 21310 52610 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 48414 20974 48466 21026
rect 4062 20862 4114 20914
rect 8654 20862 8706 20914
rect 11790 20862 11842 20914
rect 13470 20862 13522 20914
rect 13806 20862 13858 20914
rect 15262 20862 15314 20914
rect 15598 20862 15650 20914
rect 19742 20862 19794 20914
rect 20078 20862 20130 20914
rect 20414 20862 20466 20914
rect 20638 20862 20690 20914
rect 22654 20862 22706 20914
rect 23886 20862 23938 20914
rect 28142 20862 28194 20914
rect 36990 20862 37042 20914
rect 37326 20862 37378 20914
rect 38894 20862 38946 20914
rect 42142 20862 42194 20914
rect 43934 20862 43986 20914
rect 49198 20862 49250 20914
rect 49646 20862 49698 20914
rect 51662 20862 51714 20914
rect 53678 20862 53730 20914
rect 7982 20750 8034 20802
rect 8430 20750 8482 20802
rect 15822 20750 15874 20802
rect 16382 20750 16434 20802
rect 27022 20750 27074 20802
rect 27470 20750 27522 20802
rect 34638 20750 34690 20802
rect 34974 20750 35026 20802
rect 44942 20750 44994 20802
rect 45390 20750 45442 20802
rect 51550 20750 51602 20802
rect 3054 20638 3106 20690
rect 9662 20638 9714 20690
rect 10894 20638 10946 20690
rect 21646 20638 21698 20690
rect 24782 20638 24834 20690
rect 32286 20638 32338 20690
rect 39902 20638 39954 20690
rect 43150 20638 43202 20690
rect 44270 20638 44322 20690
rect 50654 20638 50706 20690
rect 54686 20638 54738 20690
rect 18734 20526 18786 20578
rect 19518 20526 19570 20578
rect 23214 20526 23266 20578
rect 23998 20526 24050 20578
rect 31502 20526 31554 20578
rect 47742 20526 47794 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4846 20190 4898 20242
rect 24222 20190 24274 20242
rect 24670 20190 24722 20242
rect 46286 20190 46338 20242
rect 8318 20078 8370 20130
rect 9886 20078 9938 20130
rect 13470 20078 13522 20130
rect 16494 20078 16546 20130
rect 16830 20078 16882 20130
rect 17502 20078 17554 20130
rect 18174 20078 18226 20130
rect 18510 20078 18562 20130
rect 21982 20078 22034 20130
rect 26014 20078 26066 20130
rect 29710 20078 29762 20130
rect 33182 20078 33234 20130
rect 37886 20078 37938 20130
rect 45054 20078 45106 20130
rect 46734 20078 46786 20130
rect 47070 20078 47122 20130
rect 47742 20078 47794 20130
rect 48190 20078 48242 20130
rect 48862 20078 48914 20130
rect 50766 20078 50818 20130
rect 53902 20078 53954 20130
rect 54686 20078 54738 20130
rect 7198 19966 7250 20018
rect 7758 19966 7810 20018
rect 14926 19966 14978 20018
rect 17838 19966 17890 20018
rect 18846 19966 18898 20018
rect 19070 19966 19122 20018
rect 19630 19966 19682 20018
rect 23550 19966 23602 20018
rect 42366 19966 42418 20018
rect 42814 19966 42866 20018
rect 47518 19966 47570 20018
rect 54462 19966 54514 20018
rect 7982 19854 8034 19906
rect 8766 19854 8818 19906
rect 8990 19854 9042 19906
rect 11006 19854 11058 19906
rect 15486 19854 15538 19906
rect 25454 19854 25506 19906
rect 27134 19854 27186 19906
rect 30606 19854 30658 19906
rect 34302 19854 34354 19906
rect 36878 19854 36930 19906
rect 46398 19854 46450 19906
rect 49758 19854 49810 19906
rect 52558 19854 52610 19906
rect 4062 19742 4114 19794
rect 22766 19742 22818 19794
rect 23774 19742 23826 19794
rect 45838 19742 45890 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 8318 19294 8370 19346
rect 11790 19294 11842 19346
rect 16830 19294 16882 19346
rect 19742 19294 19794 19346
rect 20638 19294 20690 19346
rect 21422 19294 21474 19346
rect 21870 19294 21922 19346
rect 26574 19294 26626 19346
rect 31054 19294 31106 19346
rect 33518 19294 33570 19346
rect 38334 19294 38386 19346
rect 41582 19294 41634 19346
rect 43710 19294 43762 19346
rect 44382 19294 44434 19346
rect 45054 19294 45106 19346
rect 45502 19294 45554 19346
rect 46062 19294 46114 19346
rect 48638 19294 48690 19346
rect 50878 19294 50930 19346
rect 51102 19294 51154 19346
rect 54014 19294 54066 19346
rect 22542 19182 22594 19234
rect 23102 19182 23154 19234
rect 9550 19070 9602 19122
rect 10558 19070 10610 19122
rect 15598 19070 15650 19122
rect 18734 19070 18786 19122
rect 25454 19070 25506 19122
rect 30046 19070 30098 19122
rect 34526 19070 34578 19122
rect 39342 19070 39394 19122
rect 42590 19070 42642 19122
rect 47070 19070 47122 19122
rect 49646 19070 49698 19122
rect 55022 19070 55074 19122
rect 20302 18958 20354 19010
rect 21982 18958 22034 19010
rect 26238 18958 26290 19010
rect 43598 18958 43650 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 23886 18622 23938 18674
rect 4062 18510 4114 18562
rect 6638 18510 6690 18562
rect 9886 18510 9938 18562
rect 13358 18510 13410 18562
rect 18286 18510 18338 18562
rect 22990 18510 23042 18562
rect 28926 18510 28978 18562
rect 29486 18510 29538 18562
rect 33630 18510 33682 18562
rect 38446 18510 38498 18562
rect 42926 18510 42978 18562
rect 45726 18510 45778 18562
rect 46846 18510 46898 18562
rect 47854 18510 47906 18562
rect 51550 18510 51602 18562
rect 47182 18398 47234 18450
rect 5182 18286 5234 18338
rect 7870 18286 7922 18338
rect 11118 18286 11170 18338
rect 14478 18286 14530 18338
rect 19518 18286 19570 18338
rect 21870 18286 21922 18338
rect 27806 18286 27858 18338
rect 30830 18286 30882 18338
rect 34750 18286 34802 18338
rect 37326 18286 37378 18338
rect 41918 18286 41970 18338
rect 44718 18286 44770 18338
rect 48078 18286 48130 18338
rect 50206 18286 50258 18338
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 8654 17726 8706 17778
rect 11902 17726 11954 17778
rect 16606 17726 16658 17778
rect 19742 17726 19794 17778
rect 24782 17726 24834 17778
rect 27134 17726 27186 17778
rect 32398 17726 32450 17778
rect 35422 17726 35474 17778
rect 40126 17726 40178 17778
rect 45838 17726 45890 17778
rect 48638 17726 48690 17778
rect 9662 17502 9714 17554
rect 10782 17502 10834 17554
rect 17502 17502 17554 17554
rect 18734 17502 18786 17554
rect 23774 17502 23826 17554
rect 28366 17502 28418 17554
rect 31502 17502 31554 17554
rect 34414 17502 34466 17554
rect 41134 17502 41186 17554
rect 47070 17502 47122 17554
rect 49646 17502 49698 17554
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 12686 16942 12738 16994
rect 16718 16942 16770 16994
rect 18398 16942 18450 16994
rect 20974 16942 21026 16994
rect 28702 16942 28754 16994
rect 29374 16942 29426 16994
rect 35310 16942 35362 16994
rect 38894 16942 38946 16994
rect 43038 16942 43090 16994
rect 46062 16942 46114 16994
rect 11342 16718 11394 16770
rect 15598 16718 15650 16770
rect 19406 16718 19458 16770
rect 22318 16718 22370 16770
rect 27470 16718 27522 16770
rect 30718 16718 30770 16770
rect 34190 16718 34242 16770
rect 38110 16718 38162 16770
rect 41918 16718 41970 16770
rect 44718 16718 44770 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 9998 16158 10050 16210
rect 14814 16158 14866 16210
rect 18734 16158 18786 16210
rect 22654 16158 22706 16210
rect 26462 16158 26514 16210
rect 31950 16158 32002 16210
rect 35310 16158 35362 16210
rect 39118 16158 39170 16210
rect 42590 16158 42642 16210
rect 10894 15934 10946 15986
rect 16158 15934 16210 15986
rect 19742 15934 19794 15986
rect 23662 15934 23714 15986
rect 27246 15934 27298 15986
rect 33294 15934 33346 15986
rect 33966 15934 34018 15986
rect 37998 15934 38050 15986
rect 43710 15934 43762 15986
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 21310 15374 21362 15426
rect 22542 15374 22594 15426
rect 29598 15374 29650 15426
rect 32062 15374 32114 15426
rect 36766 15374 36818 15426
rect 20302 15150 20354 15202
rect 23550 15150 23602 15202
rect 28254 15150 28306 15202
rect 31166 15150 31218 15202
rect 35758 15150 35810 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 18174 14590 18226 14642
rect 23326 14590 23378 14642
rect 27358 14590 27410 14642
rect 30158 14590 30210 14642
rect 19182 14366 19234 14418
rect 24334 14366 24386 14418
rect 26350 14366 26402 14418
rect 31278 14366 31330 14418
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 40574 3278 40626 3330
rect 41246 3278 41298 3330
rect 43934 3278 43986 3330
rect 44606 3278 44658 3330
rect 48638 3278 48690 3330
rect 55022 3278 55074 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 56448 67200 56560 68000
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 56476 64148 56532 67200
rect 56700 64148 56756 64158
rect 56476 64146 56756 64148
rect 56476 64094 56702 64146
rect 56754 64094 56756 64146
rect 56476 64092 56756 64094
rect 56700 64082 56756 64092
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 66220 62914 66276 62926
rect 66220 62862 66222 62914
rect 66274 62862 66276 62914
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 66220 62580 66276 62862
rect 66220 62514 66276 62524
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 43708 54626 43764 54638
rect 43708 54574 43710 54626
rect 43762 54574 43764 54626
rect 41468 54404 41524 54414
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 28588 53844 28644 53854
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 27244 52274 27300 52286
rect 27244 52222 27246 52274
rect 27298 52222 27300 52274
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 23660 51492 23716 51502
rect 23660 51490 24500 51492
rect 23660 51438 23662 51490
rect 23714 51438 24500 51490
rect 23660 51436 24500 51438
rect 23660 51426 23716 51436
rect 22316 51266 22372 51278
rect 22316 51214 22318 51266
rect 22370 51214 22372 51266
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 19628 49138 19684 49150
rect 19628 49086 19630 49138
rect 19682 49086 19684 49138
rect 18508 48914 18564 48926
rect 18508 48862 18510 48914
rect 18562 48862 18564 48914
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 10892 47684 10948 47694
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 10780 41074 10836 41086
rect 10780 41022 10782 41074
rect 10834 41022 10836 41074
rect 10780 40628 10836 41022
rect 10780 40562 10836 40572
rect 9996 40404 10052 40414
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 9100 39732 9156 39742
rect 9100 39638 9156 39676
rect 8092 39506 8148 39518
rect 8092 39454 8094 39506
rect 8146 39454 8148 39506
rect 6972 38946 7028 38958
rect 6972 38894 6974 38946
rect 7026 38894 7028 38946
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 6972 38164 7028 38894
rect 7980 38722 8036 38734
rect 7980 38670 7982 38722
rect 8034 38670 8036 38722
rect 7980 38388 8036 38670
rect 7980 38322 8036 38332
rect 6972 38098 7028 38108
rect 7868 38162 7924 38174
rect 7868 38110 7870 38162
rect 7922 38110 7924 38162
rect 7084 37938 7140 37950
rect 7084 37886 7086 37938
rect 7138 37886 7140 37938
rect 4172 37380 4228 37390
rect 6972 37380 7028 37390
rect 4172 37378 4340 37380
rect 4172 37326 4174 37378
rect 4226 37326 4340 37378
rect 4172 37324 4340 37326
rect 4172 37314 4228 37324
rect 3948 36594 4004 36606
rect 3948 36542 3950 36594
rect 4002 36542 4004 36594
rect 1708 36372 1764 36382
rect 1764 36316 1876 36372
rect 1708 36278 1764 36316
rect 1820 35922 1876 36316
rect 3052 36370 3108 36382
rect 3052 36318 3054 36370
rect 3106 36318 3108 36370
rect 1820 35870 1822 35922
rect 1874 35870 1876 35922
rect 1820 35858 1876 35870
rect 2044 36258 2100 36270
rect 2044 36206 2046 36258
rect 2098 36206 2100 36258
rect 2044 35924 2100 36206
rect 2044 35858 2100 35868
rect 3052 35700 3108 36318
rect 3052 35634 3108 35644
rect 3836 35026 3892 35038
rect 3836 34974 3838 35026
rect 3890 34974 3892 35026
rect 3052 34916 3108 34926
rect 3052 34802 3108 34860
rect 3052 34750 3054 34802
rect 3106 34750 3108 34802
rect 3052 34738 3108 34750
rect 3836 33348 3892 34974
rect 3836 33282 3892 33292
rect 3052 33234 3108 33246
rect 3052 33182 3054 33234
rect 3106 33182 3108 33234
rect 3052 33124 3108 33182
rect 3052 33058 3108 33068
rect 3052 31668 3108 31678
rect 3052 31574 3108 31612
rect 3948 31556 4004 36542
rect 4172 35812 4228 35822
rect 4172 35718 4228 35756
rect 4172 34242 4228 34254
rect 4172 34190 4174 34242
rect 4226 34190 4228 34242
rect 4172 34132 4228 34190
rect 4172 34066 4228 34076
rect 4284 33572 4340 37324
rect 6972 37286 7028 37324
rect 5180 37268 5236 37278
rect 5180 37154 5236 37212
rect 5180 37102 5182 37154
rect 5234 37102 5236 37154
rect 5180 37090 5236 37102
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 7084 36708 7140 37886
rect 7084 36642 7140 36652
rect 7868 36484 7924 38110
rect 8092 37828 8148 39454
rect 9996 38722 10052 40348
rect 10780 39506 10836 39518
rect 10780 39454 10782 39506
rect 10834 39454 10836 39506
rect 10780 39396 10836 39454
rect 10780 39330 10836 39340
rect 9996 38670 9998 38722
rect 10050 38670 10052 38722
rect 9996 38658 10052 38670
rect 10220 38722 10276 38734
rect 10220 38670 10222 38722
rect 10274 38670 10276 38722
rect 9884 38388 9940 38398
rect 8092 37762 8148 37772
rect 9324 38050 9380 38062
rect 9324 37998 9326 38050
rect 9378 37998 9380 38050
rect 8652 37268 8708 37278
rect 7980 37156 8036 37166
rect 7980 37062 8036 37100
rect 8092 36596 8148 36606
rect 8092 36502 8148 36540
rect 7980 36484 8036 36494
rect 7868 36428 7980 36484
rect 7980 36418 8036 36428
rect 7084 36370 7140 36382
rect 7084 36318 7086 36370
rect 7138 36318 7140 36370
rect 7084 36148 7140 36318
rect 7084 36082 7140 36092
rect 6972 35810 7028 35822
rect 6972 35758 6974 35810
rect 7026 35758 7028 35810
rect 5180 35586 5236 35598
rect 5180 35534 5182 35586
rect 5234 35534 5236 35586
rect 5180 35364 5236 35534
rect 6972 35476 7028 35758
rect 6972 35410 7028 35420
rect 7980 35586 8036 35598
rect 7980 35534 7982 35586
rect 8034 35534 8036 35586
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 5180 35298 5236 35308
rect 4476 35242 4740 35252
rect 7308 35028 7364 35038
rect 7308 34934 7364 34972
rect 6300 34804 6356 34814
rect 6300 34710 6356 34748
rect 7980 34356 8036 35534
rect 8652 34692 8708 37212
rect 9324 37268 9380 37998
rect 9884 38050 9940 38332
rect 9884 37998 9886 38050
rect 9938 37998 9940 38050
rect 9884 37986 9940 37998
rect 9324 36482 9380 37212
rect 10220 36820 10276 38670
rect 10220 36754 10276 36764
rect 9324 36430 9326 36482
rect 9378 36430 9380 36482
rect 9324 36372 9380 36430
rect 9884 36484 9940 36494
rect 9884 36390 9940 36428
rect 8988 36316 9380 36372
rect 8764 34916 8820 34926
rect 8988 34916 9044 36316
rect 10892 36260 10948 47628
rect 17164 47236 17220 47246
rect 17164 46114 17220 47180
rect 18508 47236 18564 48862
rect 19516 48354 19572 48366
rect 19516 48302 19518 48354
rect 19570 48302 19572 48354
rect 19516 47796 19572 48302
rect 19628 48132 19684 49086
rect 21532 48916 21588 48926
rect 20972 48914 21588 48916
rect 20972 48862 21534 48914
rect 21586 48862 21588 48914
rect 20972 48860 21588 48862
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20300 48580 20356 48590
rect 19740 48132 19796 48142
rect 19628 48076 19740 48132
rect 19740 48066 19796 48076
rect 19516 47740 19684 47796
rect 19516 47570 19572 47582
rect 19516 47518 19518 47570
rect 19570 47518 19572 47570
rect 18508 47170 18564 47180
rect 18620 47346 18676 47358
rect 18620 47294 18622 47346
rect 18674 47294 18676 47346
rect 17724 46788 17780 46798
rect 17164 46062 17166 46114
rect 17218 46062 17220 46114
rect 17164 46050 17220 46062
rect 17276 46786 17780 46788
rect 17276 46734 17726 46786
rect 17778 46734 17780 46786
rect 17276 46732 17780 46734
rect 17164 45668 17220 45678
rect 16940 44994 16996 45006
rect 16940 44942 16942 44994
rect 16994 44942 16996 44994
rect 16940 44884 16996 44942
rect 16940 44818 16996 44828
rect 17164 44546 17220 45612
rect 17164 44494 17166 44546
rect 17218 44494 17220 44546
rect 17164 44482 17220 44494
rect 14812 44436 14868 44446
rect 14028 44434 14868 44436
rect 14028 44382 14814 44434
rect 14866 44382 14868 44434
rect 14028 44380 14868 44382
rect 12012 42082 12068 42094
rect 12012 42030 12014 42082
rect 12066 42030 12068 42082
rect 11900 41298 11956 41310
rect 11900 41246 11902 41298
rect 11954 41246 11956 41298
rect 11676 40628 11732 40638
rect 11676 40534 11732 40572
rect 11900 39956 11956 41246
rect 12012 40628 12068 42030
rect 13020 41858 13076 41870
rect 13020 41806 13022 41858
rect 13074 41806 13076 41858
rect 12012 40562 12068 40572
rect 12236 40626 12292 40638
rect 12236 40574 12238 40626
rect 12290 40574 12292 40626
rect 12236 40404 12292 40574
rect 12236 40338 12292 40348
rect 11900 39890 11956 39900
rect 11900 39730 11956 39742
rect 11900 39678 11902 39730
rect 11954 39678 11956 39730
rect 11900 39620 11956 39678
rect 11900 39554 11956 39564
rect 12012 39060 12068 39070
rect 11004 38948 11060 38958
rect 11004 38854 11060 38892
rect 12012 38722 12068 39004
rect 13020 38836 13076 41806
rect 13916 39956 13972 39966
rect 13020 38770 13076 38780
rect 13468 39618 13524 39630
rect 13468 39566 13470 39618
rect 13522 39566 13524 39618
rect 13468 38834 13524 39566
rect 13468 38782 13470 38834
rect 13522 38782 13524 38834
rect 12012 38670 12014 38722
rect 12066 38670 12068 38722
rect 12012 38658 12068 38670
rect 13468 38724 13524 38782
rect 13804 38836 13860 38846
rect 13804 38742 13860 38780
rect 12908 38164 12964 38174
rect 12460 37826 12516 37838
rect 12460 37774 12462 37826
rect 12514 37774 12516 37826
rect 11004 37492 11060 37502
rect 11004 37378 11060 37436
rect 11004 37326 11006 37378
rect 11058 37326 11060 37378
rect 11004 37314 11060 37326
rect 11900 37380 11956 37390
rect 10892 36194 10948 36204
rect 11116 36708 11172 36718
rect 9884 35588 9940 35598
rect 8764 34914 9044 34916
rect 8764 34862 8766 34914
rect 8818 34862 9044 34914
rect 8764 34860 9044 34862
rect 9100 34914 9156 34926
rect 9100 34862 9102 34914
rect 9154 34862 9156 34914
rect 8764 34850 8820 34860
rect 9100 34692 9156 34862
rect 8652 34636 9156 34692
rect 7980 34290 8036 34300
rect 6972 34244 7028 34254
rect 6972 34150 7028 34188
rect 9100 34132 9156 34142
rect 5180 34018 5236 34030
rect 5180 33966 5182 34018
rect 5234 33966 5236 34018
rect 5180 33908 5236 33966
rect 7980 34020 8036 34030
rect 7980 33926 8036 33964
rect 5180 33842 5236 33852
rect 7868 33796 7924 33806
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33506 4340 33516
rect 4060 33460 4116 33470
rect 4060 33366 4116 33404
rect 7868 33458 7924 33740
rect 7868 33406 7870 33458
rect 7922 33406 7924 33458
rect 7868 33394 7924 33406
rect 8316 33572 8372 33582
rect 6636 33234 6692 33246
rect 6636 33182 6638 33234
rect 6690 33182 6692 33234
rect 4172 33012 4228 33022
rect 4172 32674 4228 32956
rect 6636 32788 6692 33182
rect 6636 32722 6692 32732
rect 4172 32622 4174 32674
rect 4226 32622 4228 32674
rect 4172 32610 4228 32622
rect 6972 32676 7028 32686
rect 6972 32582 7028 32620
rect 5180 32450 5236 32462
rect 5180 32398 5182 32450
rect 5234 32398 5236 32450
rect 5180 32228 5236 32398
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 5180 32162 5236 32172
rect 7980 32450 8036 32462
rect 7980 32398 7982 32450
rect 8034 32398 8036 32450
rect 4476 32106 4740 32116
rect 7980 31948 8036 32398
rect 4060 31892 4116 31902
rect 4060 31798 4116 31836
rect 7868 31890 7924 31902
rect 7980 31892 8260 31948
rect 7868 31838 7870 31890
rect 7922 31838 7924 31890
rect 3948 31490 4004 31500
rect 5292 31668 5348 31678
rect 2156 31108 2212 31118
rect 2156 31014 2212 31052
rect 5180 31106 5236 31118
rect 5180 31054 5182 31106
rect 5234 31054 5236 31106
rect 3164 30884 3220 30894
rect 3164 30790 3220 30828
rect 2828 30772 2884 30782
rect 2044 28644 2100 28654
rect 1820 27858 1876 27870
rect 1820 27806 1822 27858
rect 1874 27806 1876 27858
rect 1820 26292 1876 27806
rect 2044 26402 2100 28588
rect 2044 26350 2046 26402
rect 2098 26350 2100 26402
rect 2044 26338 2100 26350
rect 2268 27858 2324 27870
rect 2268 27806 2270 27858
rect 2322 27806 2324 27858
rect 1708 25394 1764 25406
rect 1708 25342 1710 25394
rect 1762 25342 1764 25394
rect 1708 24948 1764 25342
rect 1708 24052 1764 24892
rect 1820 24722 1876 26236
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 24658 1876 24670
rect 2044 25282 2100 25294
rect 2044 25230 2046 25282
rect 2098 25230 2100 25282
rect 2044 24724 2100 25230
rect 2156 24724 2212 24734
rect 2044 24722 2212 24724
rect 2044 24670 2158 24722
rect 2210 24670 2212 24722
rect 2044 24668 2212 24670
rect 2156 24658 2212 24668
rect 1820 24052 1876 24062
rect 1708 24050 1876 24052
rect 1708 23998 1822 24050
rect 1874 23998 1876 24050
rect 1708 23996 1876 23998
rect 1820 23986 1876 23996
rect 2268 19348 2324 27806
rect 2716 24836 2772 24846
rect 2716 22258 2772 24780
rect 2828 23266 2884 30716
rect 4396 30772 4452 30810
rect 4396 30706 4452 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5068 30436 5124 30446
rect 4060 30322 4116 30334
rect 4060 30270 4062 30322
rect 4114 30270 4116 30322
rect 4060 30212 4116 30270
rect 4060 30146 4116 30156
rect 4508 30212 4564 30222
rect 5068 30212 5124 30380
rect 4508 30210 5124 30212
rect 4508 30158 4510 30210
rect 4562 30158 5124 30210
rect 4508 30156 5124 30158
rect 3052 30100 3108 30110
rect 3052 30006 3108 30044
rect 4508 30100 4564 30156
rect 4508 30034 4564 30044
rect 3164 29764 3220 29774
rect 3164 29538 3220 29708
rect 3164 29486 3166 29538
rect 3218 29486 3220 29538
rect 3164 29474 3220 29486
rect 4172 29314 4228 29326
rect 4172 29262 4174 29314
rect 4226 29262 4228 29314
rect 4172 29204 4228 29262
rect 4172 29138 4228 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28868 4564 28878
rect 4060 28754 4116 28766
rect 4060 28702 4062 28754
rect 4114 28702 4116 28754
rect 3052 28532 3108 28542
rect 3052 28438 3108 28476
rect 3948 28308 4004 28318
rect 3052 27636 3108 27646
rect 3052 26962 3108 27580
rect 3500 27300 3556 27310
rect 3052 26910 3054 26962
rect 3106 26910 3108 26962
rect 3052 26898 3108 26910
rect 3388 27244 3500 27300
rect 3276 26180 3332 26190
rect 3388 26180 3444 27244
rect 3500 27234 3556 27244
rect 3948 27186 4004 28252
rect 4060 27860 4116 28702
rect 4508 28754 4564 28812
rect 4508 28702 4510 28754
rect 4562 28702 4564 28754
rect 4508 28532 4564 28702
rect 5180 28756 5236 31054
rect 5292 29316 5348 31612
rect 7084 31668 7140 31678
rect 7084 31574 7140 31612
rect 7868 31220 7924 31838
rect 7868 31164 8148 31220
rect 7532 30994 7588 31006
rect 7532 30942 7534 30994
rect 7586 30942 7588 30994
rect 7084 30660 7140 30670
rect 7084 30322 7140 30604
rect 7084 30270 7086 30322
rect 7138 30270 7140 30322
rect 7084 30258 7140 30270
rect 5292 29250 5348 29260
rect 6076 30098 6132 30110
rect 6076 30046 6078 30098
rect 6130 30046 6132 30098
rect 5180 28690 5236 28700
rect 5404 29202 5460 29214
rect 5404 29150 5406 29202
rect 5458 29150 5460 29202
rect 5404 28644 5460 29150
rect 6076 29092 6132 30046
rect 6188 29540 6244 29550
rect 6188 29446 6244 29484
rect 6076 29026 6132 29036
rect 6860 28756 6916 28766
rect 6860 28662 6916 28700
rect 5404 28578 5460 28588
rect 6524 28644 6580 28654
rect 6524 28550 6580 28588
rect 7196 28644 7252 28654
rect 7196 28550 7252 28588
rect 4508 28466 4564 28476
rect 6412 28420 6468 28430
rect 6412 28326 6468 28364
rect 7420 28420 7476 28430
rect 4732 28084 4788 28094
rect 4732 27990 4788 28028
rect 4060 27794 4116 27804
rect 5404 27858 5460 27870
rect 5404 27806 5406 27858
rect 5458 27806 5460 27858
rect 5292 27634 5348 27646
rect 5292 27582 5294 27634
rect 5346 27582 5348 27634
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3948 27134 3950 27186
rect 4002 27134 4004 27186
rect 3948 27122 4004 27134
rect 4060 27188 4116 27198
rect 3276 26178 3444 26180
rect 3276 26126 3278 26178
rect 3330 26126 3444 26178
rect 3276 26124 3444 26126
rect 3948 26516 4004 26526
rect 3276 26114 3332 26124
rect 2940 26068 2996 26078
rect 2940 25394 2996 26012
rect 2940 25342 2942 25394
rect 2994 25342 2996 25394
rect 2940 25330 2996 25342
rect 3836 25284 3892 25294
rect 3836 24050 3892 25228
rect 3836 23998 3838 24050
rect 3890 23998 3892 24050
rect 3836 23986 3892 23998
rect 3052 23828 3108 23838
rect 3052 23734 3108 23772
rect 2828 23214 2830 23266
rect 2882 23214 2884 23266
rect 2828 23202 2884 23214
rect 3052 23604 3108 23614
rect 2716 22206 2718 22258
rect 2770 22206 2772 22258
rect 2716 22194 2772 22206
rect 3052 20690 3108 23548
rect 3948 23042 4004 26460
rect 4060 25618 4116 27132
rect 4508 26292 4564 26302
rect 4508 26198 4564 26236
rect 5068 26290 5124 26302
rect 5068 26238 5070 26290
rect 5122 26238 5124 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4060 25566 4062 25618
rect 4114 25566 4116 25618
rect 4060 25554 4116 25566
rect 3948 22990 3950 23042
rect 4002 22990 4004 23042
rect 3948 22978 4004 22990
rect 4060 25060 4116 25070
rect 4060 22482 4116 25004
rect 5068 25060 5124 26238
rect 5068 24994 5124 25004
rect 4732 24948 4788 24958
rect 5292 24948 5348 27582
rect 4732 24854 4788 24892
rect 5180 24892 5348 24948
rect 5404 26964 5460 27806
rect 5964 27860 6020 27870
rect 5964 27766 6020 27804
rect 6636 27524 6692 27534
rect 5740 26964 5796 26974
rect 5404 26908 5740 26964
rect 5404 26292 5460 26908
rect 5740 26870 5796 26908
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 5068 24052 5124 24062
rect 5068 23958 5124 23996
rect 4060 22430 4062 22482
rect 4114 22430 4116 22482
rect 4060 22418 4116 22430
rect 4172 23156 4228 23166
rect 4060 22260 4116 22270
rect 3164 21698 3220 21710
rect 3164 21646 3166 21698
rect 3218 21646 3220 21698
rect 3164 21476 3220 21646
rect 3164 21410 3220 21420
rect 4060 20914 4116 22204
rect 4172 21474 4228 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 21422 4174 21474
rect 4226 21422 4228 21474
rect 4172 21410 4228 21422
rect 4844 21812 4900 21822
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4060 20862 4062 20914
rect 4114 20862 4116 20914
rect 4060 20850 4116 20862
rect 3052 20638 3054 20690
rect 3106 20638 3108 20690
rect 3052 20626 3108 20638
rect 4844 20242 4900 21756
rect 4844 20190 4846 20242
rect 4898 20190 4900 20242
rect 4844 20178 4900 20190
rect 5180 20244 5236 24892
rect 5404 24722 5460 26236
rect 5964 26292 6020 26302
rect 5964 25618 6020 26236
rect 5964 25566 5966 25618
rect 6018 25566 6020 25618
rect 5964 25554 6020 25566
rect 6524 26292 6580 26302
rect 5852 25282 5908 25294
rect 5852 25230 5854 25282
rect 5906 25230 5908 25282
rect 5852 24948 5908 25230
rect 6188 24948 6244 24958
rect 5852 24892 6132 24948
rect 5404 24670 5406 24722
rect 5458 24670 5460 24722
rect 5292 24498 5348 24510
rect 5292 24446 5294 24498
rect 5346 24446 5348 24498
rect 5292 23604 5348 24446
rect 5292 23538 5348 23548
rect 5404 24052 5460 24670
rect 5964 24722 6020 24734
rect 5964 24670 5966 24722
rect 6018 24670 6020 24722
rect 5852 24052 5908 24062
rect 5460 24050 5908 24052
rect 5460 23998 5854 24050
rect 5906 23998 5908 24050
rect 5460 23996 5908 23998
rect 5404 23154 5460 23996
rect 5852 23986 5908 23996
rect 5964 23380 6020 24670
rect 5404 23102 5406 23154
rect 5458 23102 5460 23154
rect 5404 22372 5460 23102
rect 5852 23324 6020 23380
rect 5516 22372 5572 22382
rect 5404 22370 5572 22372
rect 5404 22318 5518 22370
rect 5570 22318 5572 22370
rect 5404 22316 5572 22318
rect 5516 22306 5572 22316
rect 5852 22260 5908 23324
rect 5964 23156 6020 23166
rect 5964 23062 6020 23100
rect 5852 22194 5908 22204
rect 5964 21812 6020 21822
rect 6076 21812 6132 24892
rect 6188 24050 6244 24892
rect 6188 23998 6190 24050
rect 6242 23998 6244 24050
rect 6188 23986 6244 23998
rect 6524 24050 6580 26236
rect 6636 25394 6692 27468
rect 7196 26964 7252 26974
rect 7196 26870 7252 26908
rect 7420 26514 7476 28364
rect 7420 26462 7422 26514
rect 7474 26462 7476 26514
rect 7420 26450 7476 26462
rect 7532 25956 7588 30942
rect 7980 30994 8036 31006
rect 7980 30942 7982 30994
rect 8034 30942 8036 30994
rect 7644 29988 7700 29998
rect 7980 29988 8036 30942
rect 8092 30548 8148 31164
rect 8204 30772 8260 31892
rect 8204 30706 8260 30716
rect 8092 30492 8260 30548
rect 8092 29988 8148 29998
rect 7644 29986 8148 29988
rect 7644 29934 7646 29986
rect 7698 29934 8094 29986
rect 8146 29934 8148 29986
rect 7644 29932 8148 29934
rect 7644 29922 7700 29932
rect 7868 29540 7924 29550
rect 7868 28754 7924 29484
rect 8092 29428 8148 29932
rect 8204 29652 8260 30492
rect 8316 30210 8372 33516
rect 9100 33570 9156 34076
rect 9100 33518 9102 33570
rect 9154 33518 9156 33570
rect 9100 33506 9156 33518
rect 9884 33234 9940 35532
rect 11116 34354 11172 36652
rect 11452 35922 11508 35934
rect 11452 35870 11454 35922
rect 11506 35870 11508 35922
rect 11116 34302 11118 34354
rect 11170 34302 11172 34354
rect 11116 34290 11172 34302
rect 11228 35700 11284 35710
rect 9884 33182 9886 33234
rect 9938 33182 9940 33234
rect 9884 33170 9940 33182
rect 9996 34018 10052 34030
rect 9996 33966 9998 34018
rect 10050 33966 10052 34018
rect 8876 33122 8932 33134
rect 8876 33070 8878 33122
rect 8930 33070 8932 33122
rect 8876 31948 8932 33070
rect 9100 32564 9156 32574
rect 9100 32470 9156 32508
rect 9884 32564 9940 32574
rect 9884 32470 9940 32508
rect 9212 32340 9268 32350
rect 8876 31892 9156 31948
rect 9100 31798 9156 31836
rect 8652 31556 8708 31566
rect 8652 31554 8820 31556
rect 8652 31502 8654 31554
rect 8706 31502 8820 31554
rect 8652 31500 8820 31502
rect 8652 31490 8708 31500
rect 8316 30158 8318 30210
rect 8370 30158 8372 30210
rect 8316 30146 8372 30158
rect 8204 29586 8260 29596
rect 8092 29362 8148 29372
rect 8428 29428 8484 29438
rect 8764 29428 8820 31500
rect 8876 31218 8932 31230
rect 8876 31166 8878 31218
rect 8930 31166 8932 31218
rect 8876 29986 8932 31166
rect 8988 31108 9044 31118
rect 9212 31108 9268 32284
rect 8988 31106 9268 31108
rect 8988 31054 8990 31106
rect 9042 31054 9268 31106
rect 8988 31052 9268 31054
rect 9436 31892 9492 31902
rect 9436 31778 9492 31836
rect 9996 31892 10052 33966
rect 9996 31826 10052 31836
rect 10220 34018 10276 34030
rect 10220 33966 10222 34018
rect 10274 33966 10276 34018
rect 9436 31726 9438 31778
rect 9490 31726 9492 31778
rect 8988 31042 9044 31052
rect 9436 30994 9492 31726
rect 9884 31778 9940 31790
rect 9884 31726 9886 31778
rect 9938 31726 9940 31778
rect 9884 31556 9940 31726
rect 9884 31490 9940 31500
rect 9436 30942 9438 30994
rect 9490 30942 9492 30994
rect 9436 30930 9492 30942
rect 10108 30994 10164 31006
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 9884 30884 9940 30894
rect 8876 29934 8878 29986
rect 8930 29934 8932 29986
rect 8876 29922 8932 29934
rect 8988 30324 9044 30334
rect 8988 29764 9044 30268
rect 9884 30100 9940 30828
rect 9884 30034 9940 30044
rect 8428 29426 8708 29428
rect 8428 29374 8430 29426
rect 8482 29374 8708 29426
rect 8428 29372 8708 29374
rect 8428 29362 8484 29372
rect 7868 28702 7870 28754
rect 7922 28702 7924 28754
rect 7868 28690 7924 28702
rect 7644 28644 7700 28654
rect 7644 28550 7700 28588
rect 8092 28418 8148 28430
rect 8092 28366 8094 28418
rect 8146 28366 8148 28418
rect 8092 27636 8148 28366
rect 8428 28084 8484 28094
rect 8316 27972 8372 27982
rect 8316 27878 8372 27916
rect 8092 27570 8148 27580
rect 8316 26852 8372 26862
rect 8204 26066 8260 26078
rect 8204 26014 8206 26066
rect 8258 26014 8260 26066
rect 7532 25900 7700 25956
rect 6636 25342 6638 25394
rect 6690 25342 6692 25394
rect 6636 25330 6692 25342
rect 7532 25732 7588 25742
rect 6524 23998 6526 24050
rect 6578 23998 6580 24050
rect 6524 23986 6580 23998
rect 6748 23828 6804 23838
rect 6748 23734 6804 23772
rect 7532 23826 7588 25676
rect 7532 23774 7534 23826
rect 7586 23774 7588 23826
rect 7532 23762 7588 23774
rect 6020 21756 6132 21812
rect 6188 22370 6244 22382
rect 6188 22318 6190 22370
rect 6242 22318 6244 22370
rect 5964 21746 6020 21756
rect 5628 21588 5684 21598
rect 5628 21494 5684 21532
rect 5964 21586 6020 21598
rect 5964 21534 5966 21586
rect 6018 21534 6020 21586
rect 5964 20188 6020 21534
rect 5180 20178 5236 20188
rect 5292 20132 6020 20188
rect 2268 19282 2324 19292
rect 4060 19794 4116 19806
rect 4060 19742 4062 19794
rect 4114 19742 4116 19794
rect 4060 18562 4116 19742
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4060 18510 4062 18562
rect 4114 18510 4116 18562
rect 4060 18498 4116 18510
rect 5180 18340 5236 18350
rect 5292 18340 5348 20132
rect 5180 18338 5348 18340
rect 5180 18286 5182 18338
rect 5234 18286 5348 18338
rect 5180 18284 5348 18286
rect 5180 18274 5236 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 6188 17780 6244 22318
rect 7644 21924 7700 25900
rect 7756 25620 7812 25630
rect 7756 25526 7812 25564
rect 7644 21858 7700 21868
rect 7868 22036 7924 22046
rect 7756 21700 7812 21710
rect 6636 20020 6692 20030
rect 6636 18562 6692 19964
rect 6636 18510 6638 18562
rect 6690 18510 6692 18562
rect 6636 18498 6692 18510
rect 7196 20018 7252 20030
rect 7196 19966 7198 20018
rect 7250 19966 7252 20018
rect 7196 18452 7252 19966
rect 7756 20018 7812 21644
rect 7756 19966 7758 20018
rect 7810 19966 7812 20018
rect 7756 19954 7812 19966
rect 7196 18386 7252 18396
rect 7868 18338 7924 21980
rect 8204 21476 8260 26014
rect 8316 25620 8372 26796
rect 8428 26402 8484 28028
rect 8652 26516 8708 29372
rect 8764 29362 8820 29372
rect 8876 29708 9044 29764
rect 8652 26450 8708 26460
rect 8764 28644 8820 28654
rect 8428 26350 8430 26402
rect 8482 26350 8484 26402
rect 8428 26338 8484 26350
rect 8764 26402 8820 28588
rect 8876 28530 8932 29708
rect 10108 29652 10164 30942
rect 10220 30324 10276 33966
rect 10556 34018 10612 34030
rect 10556 33966 10558 34018
rect 10610 33966 10612 34018
rect 10556 33572 10612 33966
rect 10556 32340 10612 33516
rect 10668 32340 10724 32350
rect 10556 32284 10668 32340
rect 10668 32246 10724 32284
rect 11228 31948 11284 35644
rect 11340 35586 11396 35598
rect 11340 35534 11342 35586
rect 11394 35534 11396 35586
rect 11340 33572 11396 35534
rect 11452 35588 11508 35870
rect 11900 35922 11956 37324
rect 12012 37156 12068 37166
rect 12012 37062 12068 37100
rect 12460 36708 12516 37774
rect 12460 36642 12516 36652
rect 12796 36820 12852 36830
rect 12796 36596 12852 36764
rect 12908 36708 12964 38108
rect 13020 37828 13076 37838
rect 13020 37734 13076 37772
rect 13244 37268 13300 37278
rect 13468 37268 13524 38668
rect 13300 37212 13524 37268
rect 13244 37174 13300 37212
rect 13020 36708 13076 36718
rect 12908 36706 13076 36708
rect 12908 36654 13022 36706
rect 13074 36654 13076 36706
rect 12908 36652 13076 36654
rect 13020 36642 13076 36652
rect 12796 36540 12964 36596
rect 12460 36372 12516 36382
rect 12460 36258 12516 36316
rect 12460 36206 12462 36258
rect 12514 36206 12516 36258
rect 12460 36194 12516 36206
rect 11900 35870 11902 35922
rect 11954 35870 11956 35922
rect 11900 35858 11956 35870
rect 12684 36036 12740 36046
rect 12684 35922 12740 35980
rect 12684 35870 12686 35922
rect 12738 35870 12740 35922
rect 12684 35858 12740 35870
rect 11452 35522 11508 35532
rect 12796 35812 12852 35822
rect 12236 34916 12292 34926
rect 12236 34822 12292 34860
rect 12572 34804 12628 34814
rect 12348 34802 12628 34804
rect 12348 34750 12574 34802
rect 12626 34750 12628 34802
rect 12348 34748 12628 34750
rect 11676 34692 11732 34702
rect 11676 34598 11732 34636
rect 12348 34468 12404 34748
rect 12572 34738 12628 34748
rect 11900 34412 12404 34468
rect 11900 34354 11956 34412
rect 11900 34302 11902 34354
rect 11954 34302 11956 34354
rect 11900 34290 11956 34302
rect 11340 33506 11396 33516
rect 12124 33348 12180 33358
rect 12124 33254 12180 33292
rect 12572 33346 12628 33358
rect 12572 33294 12574 33346
rect 12626 33294 12628 33346
rect 12572 32562 12628 33294
rect 12572 32510 12574 32562
rect 12626 32510 12628 32562
rect 12572 31948 12628 32510
rect 11228 31892 11396 31948
rect 11340 31220 11396 31892
rect 11340 31154 11396 31164
rect 12012 31892 12068 31902
rect 10220 30258 10276 30268
rect 12012 30996 12068 31836
rect 12460 31892 12628 31948
rect 12796 31948 12852 35756
rect 12908 35026 12964 36540
rect 12908 34974 12910 35026
rect 12962 34974 12964 35026
rect 12908 34962 12964 34974
rect 13020 35364 13076 35374
rect 13020 32562 13076 35308
rect 13468 34914 13524 37212
rect 13916 37266 13972 39900
rect 14028 39618 14084 44380
rect 14812 44370 14868 44380
rect 16156 44210 16212 44222
rect 16156 44158 16158 44210
rect 16210 44158 16212 44210
rect 14812 43652 14868 43662
rect 14812 43558 14868 43596
rect 15820 43426 15876 43438
rect 15820 43374 15822 43426
rect 15874 43374 15876 43426
rect 15820 41972 15876 43374
rect 15932 42644 15988 42654
rect 15932 42550 15988 42588
rect 16156 42084 16212 44158
rect 17276 43708 17332 46732
rect 17724 46722 17780 46732
rect 17836 46564 17892 46574
rect 17724 45666 17780 45678
rect 17724 45614 17726 45666
rect 17778 45614 17780 45666
rect 17724 45218 17780 45614
rect 17724 45166 17726 45218
rect 17778 45166 17780 45218
rect 17724 45154 17780 45166
rect 17052 43652 17332 43708
rect 17500 45106 17556 45118
rect 17500 45054 17502 45106
rect 17554 45054 17556 45106
rect 17500 44884 17556 45054
rect 16828 42866 16884 42878
rect 16828 42814 16830 42866
rect 16882 42814 16884 42866
rect 16156 42018 16212 42028
rect 16716 42082 16772 42094
rect 16716 42030 16718 42082
rect 16770 42030 16772 42082
rect 15820 41906 15876 41916
rect 15372 41860 15428 41870
rect 14924 41858 15428 41860
rect 14924 41806 15374 41858
rect 15426 41806 15428 41858
rect 14924 41804 15428 41806
rect 14700 40402 14756 40414
rect 14700 40350 14702 40402
rect 14754 40350 14756 40402
rect 14700 39732 14756 40350
rect 14700 39666 14756 39676
rect 14028 39566 14030 39618
rect 14082 39566 14084 39618
rect 14028 39554 14084 39566
rect 14924 37828 14980 41804
rect 15372 41794 15428 41804
rect 15932 41076 15988 41086
rect 15932 40982 15988 41020
rect 16380 40626 16436 40638
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 15148 40402 15204 40414
rect 15148 40350 15150 40402
rect 15202 40350 15204 40402
rect 15148 38724 15204 40350
rect 16268 40404 16324 40414
rect 16268 39506 16324 40348
rect 16268 39454 16270 39506
rect 16322 39454 16324 39506
rect 16268 39442 16324 39454
rect 16268 39058 16324 39070
rect 16268 39006 16270 39058
rect 16322 39006 16324 39058
rect 15148 38658 15204 38668
rect 15820 38724 15876 38734
rect 15036 38612 15092 38622
rect 15036 38050 15092 38556
rect 15820 38162 15876 38668
rect 15820 38110 15822 38162
rect 15874 38110 15876 38162
rect 15820 38098 15876 38110
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37986 15092 37998
rect 14924 37772 15092 37828
rect 13916 37214 13918 37266
rect 13970 37214 13972 37266
rect 13916 37202 13972 37214
rect 13916 37044 13972 37054
rect 13692 36372 13748 36382
rect 13692 36278 13748 36316
rect 13468 34862 13470 34914
rect 13522 34862 13524 34914
rect 13468 34850 13524 34862
rect 13916 34914 13972 36988
rect 14028 36820 14084 36830
rect 14028 36594 14084 36764
rect 14028 36542 14030 36594
rect 14082 36542 14084 36594
rect 14028 36530 14084 36542
rect 14812 36820 14868 36830
rect 14812 36482 14868 36764
rect 14812 36430 14814 36482
rect 14866 36430 14868 36482
rect 14588 36370 14644 36382
rect 14588 36318 14590 36370
rect 14642 36318 14644 36370
rect 14588 36036 14644 36318
rect 14588 35970 14644 35980
rect 14812 35812 14868 36430
rect 14812 35746 14868 35756
rect 15036 35698 15092 37772
rect 16268 37268 16324 39006
rect 16380 37490 16436 40574
rect 16604 40516 16660 40526
rect 16492 40404 16548 40414
rect 16604 40404 16660 40460
rect 16492 40402 16660 40404
rect 16492 40350 16494 40402
rect 16546 40350 16660 40402
rect 16492 40348 16660 40350
rect 16492 40338 16548 40348
rect 16380 37438 16382 37490
rect 16434 37438 16436 37490
rect 16380 37426 16436 37438
rect 16268 37202 16324 37212
rect 15820 36708 15876 36718
rect 15036 35646 15038 35698
rect 15090 35646 15092 35698
rect 15036 35634 15092 35646
rect 15148 36258 15204 36270
rect 15148 36206 15150 36258
rect 15202 36206 15204 36258
rect 15148 35476 15204 36206
rect 15820 35810 15876 36652
rect 15932 36260 15988 36270
rect 15932 36258 16548 36260
rect 15932 36206 15934 36258
rect 15986 36206 16548 36258
rect 15932 36204 16548 36206
rect 15932 36194 15988 36204
rect 15820 35758 15822 35810
rect 15874 35758 15876 35810
rect 15820 35746 15876 35758
rect 16044 35812 16100 35822
rect 15372 35700 15428 35710
rect 16044 35700 16100 35756
rect 16492 35810 16548 36204
rect 16492 35758 16494 35810
rect 16546 35758 16548 35810
rect 16492 35746 16548 35758
rect 16604 35812 16660 40348
rect 16716 39956 16772 42030
rect 16828 41636 16884 42814
rect 16828 41570 16884 41580
rect 16940 42084 16996 42094
rect 16716 39890 16772 39900
rect 16828 41298 16884 41310
rect 16828 41246 16830 41298
rect 16882 41246 16884 41298
rect 16828 39732 16884 41246
rect 16828 39666 16884 39676
rect 16940 39058 16996 42028
rect 17052 39842 17108 43652
rect 17500 43538 17556 44828
rect 17724 44098 17780 44110
rect 17724 44046 17726 44098
rect 17778 44046 17780 44098
rect 17724 43650 17780 44046
rect 17724 43598 17726 43650
rect 17778 43598 17780 43650
rect 17724 43586 17780 43598
rect 17500 43486 17502 43538
rect 17554 43486 17556 43538
rect 17500 42980 17556 43486
rect 17612 42980 17668 42990
rect 17500 42978 17668 42980
rect 17500 42926 17614 42978
rect 17666 42926 17668 42978
rect 17500 42924 17668 42926
rect 17612 42914 17668 42924
rect 17836 42308 17892 46508
rect 18620 45668 18676 47294
rect 18844 46564 18900 46574
rect 18844 46470 18900 46508
rect 19516 46116 19572 47518
rect 19628 46452 19684 47740
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19628 46386 19684 46396
rect 19516 46050 19572 46060
rect 20300 45890 20356 48524
rect 20860 48130 20916 48142
rect 20860 48078 20862 48130
rect 20914 48078 20916 48130
rect 20860 47012 20916 48078
rect 20860 46946 20916 46956
rect 20300 45838 20302 45890
rect 20354 45838 20356 45890
rect 20300 45826 20356 45838
rect 20860 46674 20916 46686
rect 20860 46622 20862 46674
rect 20914 46622 20916 46674
rect 20860 45892 20916 46622
rect 20300 45668 20356 45678
rect 18620 45602 18676 45612
rect 20188 45612 20300 45668
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 18396 45218 18452 45230
rect 18396 45166 18398 45218
rect 18450 45166 18452 45218
rect 18060 43426 18116 43438
rect 18060 43374 18062 43426
rect 18114 43374 18116 43426
rect 17948 42978 18004 42990
rect 17948 42926 17950 42978
rect 18002 42926 18004 42978
rect 17948 42866 18004 42926
rect 17948 42814 17950 42866
rect 18002 42814 18004 42866
rect 17948 42802 18004 42814
rect 17836 42252 18004 42308
rect 17836 42084 17892 42094
rect 17836 41990 17892 42028
rect 17724 41636 17780 41646
rect 17276 40628 17332 40638
rect 17332 40572 17444 40628
rect 17276 40562 17332 40572
rect 17052 39790 17054 39842
rect 17106 39790 17108 39842
rect 17052 39778 17108 39790
rect 16940 39006 16942 39058
rect 16994 39006 16996 39058
rect 16940 38994 16996 39006
rect 17164 39618 17220 39630
rect 17164 39566 17166 39618
rect 17218 39566 17220 39618
rect 17164 38836 17220 39566
rect 17276 38836 17332 38846
rect 17164 38834 17332 38836
rect 17164 38782 17278 38834
rect 17330 38782 17332 38834
rect 17164 38780 17332 38782
rect 17164 38724 17220 38780
rect 17276 38770 17332 38780
rect 17164 38658 17220 38668
rect 17388 38500 17444 40572
rect 17500 40404 17556 40414
rect 17500 40310 17556 40348
rect 17724 40404 17780 41580
rect 17836 40516 17892 40526
rect 17836 40422 17892 40460
rect 17724 40338 17780 40348
rect 17724 39620 17780 39630
rect 17724 39526 17780 39564
rect 17836 38836 17892 38846
rect 17948 38836 18004 42252
rect 17836 38834 18004 38836
rect 17836 38782 17838 38834
rect 17890 38782 18004 38834
rect 17836 38780 18004 38782
rect 17836 38770 17892 38780
rect 16940 38444 17444 38500
rect 16940 37490 16996 38444
rect 16940 37438 16942 37490
rect 16994 37438 16996 37490
rect 16940 37426 16996 37438
rect 17276 37268 17332 37278
rect 17164 37266 17332 37268
rect 17164 37214 17278 37266
rect 17330 37214 17332 37266
rect 17164 37212 17332 37214
rect 17052 36148 17108 36158
rect 16716 35812 16772 35822
rect 16604 35756 16716 35812
rect 15148 35410 15204 35420
rect 15260 35698 15428 35700
rect 15260 35646 15374 35698
rect 15426 35646 15428 35698
rect 15260 35644 15428 35646
rect 13916 34862 13918 34914
rect 13970 34862 13972 34914
rect 13916 34850 13972 34862
rect 15260 34916 15316 35644
rect 15372 35634 15428 35644
rect 15932 35698 16100 35700
rect 15932 35646 16046 35698
rect 16098 35646 16100 35698
rect 15932 35644 16100 35646
rect 13468 34692 13524 34702
rect 13468 33458 13524 34636
rect 15260 34354 15316 34860
rect 15260 34302 15262 34354
rect 15314 34302 15316 34354
rect 15260 34290 15316 34302
rect 14140 34132 14196 34142
rect 14140 34038 14196 34076
rect 14700 34130 14756 34142
rect 14700 34078 14702 34130
rect 14754 34078 14756 34130
rect 13468 33406 13470 33458
rect 13522 33406 13524 33458
rect 13468 33394 13524 33406
rect 13580 34020 13636 34030
rect 13020 32510 13022 32562
rect 13074 32510 13076 32562
rect 13020 32498 13076 32510
rect 12796 31892 13076 31948
rect 12460 31826 12516 31836
rect 13020 31890 13076 31892
rect 13020 31838 13022 31890
rect 13074 31838 13076 31890
rect 13020 31826 13076 31838
rect 13580 31892 13636 33964
rect 14700 34020 14756 34078
rect 13804 33572 13860 33582
rect 13580 31826 13636 31836
rect 13692 33460 13748 33470
rect 13356 31780 13412 31790
rect 13244 31778 13412 31780
rect 13244 31726 13358 31778
rect 13410 31726 13412 31778
rect 13244 31724 13412 31726
rect 11340 30212 11396 30222
rect 11340 30118 11396 30156
rect 12012 30212 12068 30940
rect 12348 31554 12404 31566
rect 12348 31502 12350 31554
rect 12402 31502 12404 31554
rect 12348 30212 12404 31502
rect 12460 31218 12516 31230
rect 12460 31166 12462 31218
rect 12514 31166 12516 31218
rect 12460 30322 12516 31166
rect 13132 31220 13188 31230
rect 13132 31126 13188 31164
rect 13244 30996 13300 31724
rect 13356 31714 13412 31724
rect 13692 30996 13748 33404
rect 13804 33458 13860 33516
rect 13804 33406 13806 33458
rect 13858 33406 13860 33458
rect 13804 33394 13860 33406
rect 13916 31778 13972 31790
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 13804 30996 13860 31006
rect 13692 30994 13860 30996
rect 13692 30942 13806 30994
rect 13858 30942 13860 30994
rect 13692 30940 13860 30942
rect 13244 30902 13300 30940
rect 13804 30930 13860 30940
rect 13916 30660 13972 31726
rect 13916 30594 13972 30604
rect 14700 30996 14756 33964
rect 15820 34020 15876 34030
rect 15820 33926 15876 33964
rect 12460 30270 12462 30322
rect 12514 30270 12516 30322
rect 12460 30258 12516 30270
rect 14700 30324 14756 30940
rect 14700 30230 14756 30268
rect 15036 33572 15092 33582
rect 15036 32452 15092 33516
rect 15932 33570 15988 35644
rect 16044 35634 16100 35644
rect 16716 35698 16772 35756
rect 16716 35646 16718 35698
rect 16770 35646 16772 35698
rect 16716 35634 16772 35646
rect 16492 35364 16548 35374
rect 16492 34690 16548 35308
rect 17052 35138 17108 36092
rect 17052 35086 17054 35138
rect 17106 35086 17108 35138
rect 17052 35074 17108 35086
rect 17164 35588 17220 37212
rect 17276 37202 17332 37212
rect 17388 37268 17444 37278
rect 17388 35810 17444 37212
rect 17948 37268 18004 37278
rect 18060 37268 18116 43374
rect 18396 42980 18452 45166
rect 19516 44996 19572 45006
rect 19516 44902 19572 44940
rect 20188 44322 20244 45612
rect 20300 45602 20356 45612
rect 20860 45106 20916 45836
rect 20860 45054 20862 45106
rect 20914 45054 20916 45106
rect 20860 44324 20916 45054
rect 20188 44270 20190 44322
rect 20242 44270 20244 44322
rect 20188 44258 20244 44270
rect 20300 44322 20916 44324
rect 20300 44270 20862 44322
rect 20914 44270 20916 44322
rect 20300 44268 20916 44270
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 18396 42914 18452 42924
rect 19404 43650 19460 43662
rect 19404 43598 19406 43650
rect 19458 43598 19460 43650
rect 18732 42642 18788 42654
rect 18732 42590 18734 42642
rect 18786 42590 18788 42642
rect 18732 41860 18788 42590
rect 18732 41794 18788 41804
rect 18844 41860 18900 41870
rect 18844 41858 19012 41860
rect 18844 41806 18846 41858
rect 18898 41806 19012 41858
rect 18844 41804 19012 41806
rect 18844 41794 18900 41804
rect 18732 41636 18788 41646
rect 18732 41074 18788 41580
rect 18732 41022 18734 41074
rect 18786 41022 18788 41074
rect 18732 41010 18788 41022
rect 18844 40514 18900 40526
rect 18844 40462 18846 40514
rect 18898 40462 18900 40514
rect 17948 37266 18116 37268
rect 17948 37214 17950 37266
rect 18002 37214 18116 37266
rect 17948 37212 18116 37214
rect 18396 38724 18452 38734
rect 17948 37202 18004 37212
rect 18172 36484 18228 36494
rect 18396 36484 18452 38668
rect 18844 38276 18900 40462
rect 18844 38210 18900 38220
rect 18620 36484 18676 36494
rect 18396 36482 18676 36484
rect 18396 36430 18622 36482
rect 18674 36430 18676 36482
rect 18396 36428 18676 36430
rect 18172 36390 18228 36428
rect 18620 36418 18676 36428
rect 18956 36484 19012 41804
rect 19404 38388 19460 43598
rect 19404 38322 19460 38332
rect 19516 42866 19572 42878
rect 19516 42814 19518 42866
rect 19570 42814 19572 42866
rect 19516 38052 19572 42814
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20300 41970 20356 44268
rect 20860 44258 20916 44268
rect 20972 44100 21028 48860
rect 21532 48850 21588 48860
rect 22316 48580 22372 51214
rect 23884 49924 23940 49934
rect 23884 49922 24052 49924
rect 23884 49870 23886 49922
rect 23938 49870 24052 49922
rect 23884 49868 24052 49870
rect 23884 49858 23940 49868
rect 22316 48514 22372 48524
rect 22540 49698 22596 49710
rect 22540 49646 22542 49698
rect 22594 49646 22596 49698
rect 21308 48132 21364 48142
rect 21308 46674 21364 48076
rect 21308 46622 21310 46674
rect 21362 46622 21364 46674
rect 21308 46610 21364 46622
rect 21644 47348 21700 47358
rect 21308 46116 21364 46126
rect 21308 45106 21364 46060
rect 21420 45892 21476 45902
rect 21420 45798 21476 45836
rect 21308 45054 21310 45106
rect 21362 45054 21364 45106
rect 21308 45042 21364 45054
rect 21644 44884 21700 47292
rect 21980 47346 22036 47358
rect 21980 47294 21982 47346
rect 22034 47294 22036 47346
rect 21756 47012 21812 47022
rect 21756 45890 21812 46956
rect 21980 46228 22036 47294
rect 22428 47348 22484 47358
rect 22428 47254 22484 47292
rect 21980 46162 22036 46172
rect 21756 45838 21758 45890
rect 21810 45838 21812 45890
rect 21756 45826 21812 45838
rect 22540 45668 22596 49646
rect 22876 49138 22932 49150
rect 22876 49086 22878 49138
rect 22930 49086 22932 49138
rect 22652 48354 22708 48366
rect 22652 48302 22654 48354
rect 22706 48302 22708 48354
rect 22652 46116 22708 48302
rect 22876 47124 22932 49086
rect 23660 48130 23716 48142
rect 23660 48078 23662 48130
rect 23714 48078 23716 48130
rect 22876 47058 22932 47068
rect 23436 47570 23492 47582
rect 23436 47518 23438 47570
rect 23490 47518 23492 47570
rect 22652 46050 22708 46060
rect 23436 45668 23492 47518
rect 23660 47012 23716 48078
rect 23884 48132 23940 48142
rect 23660 46946 23716 46956
rect 23772 47124 23828 47134
rect 23772 46676 23828 47068
rect 23884 46898 23940 48076
rect 23884 46846 23886 46898
rect 23938 46846 23940 46898
rect 23884 46834 23940 46846
rect 23772 46620 23940 46676
rect 23772 46340 23828 46350
rect 23660 46228 23716 46238
rect 23548 45668 23604 45678
rect 23436 45612 23548 45668
rect 22540 45602 22596 45612
rect 23548 45602 23604 45612
rect 23660 45330 23716 46172
rect 23660 45278 23662 45330
rect 23714 45278 23716 45330
rect 23660 45266 23716 45278
rect 21644 44818 21700 44828
rect 23660 44884 23716 44894
rect 23100 44434 23156 44446
rect 23100 44382 23102 44434
rect 23154 44382 23156 44434
rect 20748 44044 21028 44100
rect 22092 44210 22148 44222
rect 22092 44158 22094 44210
rect 22146 44158 22148 44210
rect 20748 43650 20804 44044
rect 20748 43598 20750 43650
rect 20802 43598 20804 43650
rect 20748 43586 20804 43598
rect 20860 43652 20916 43662
rect 20300 41918 20302 41970
rect 20354 41918 20356 41970
rect 20300 41906 20356 41918
rect 20636 41972 20692 41982
rect 20636 41878 20692 41916
rect 19740 41300 19796 41310
rect 19740 41206 19796 41244
rect 20748 40964 20804 40974
rect 20748 40870 20804 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20300 40402 20356 40414
rect 20300 40350 20302 40402
rect 20354 40350 20356 40402
rect 19852 40292 19908 40302
rect 19852 40198 19908 40236
rect 20188 39508 20244 39518
rect 20188 39394 20244 39452
rect 20188 39342 20190 39394
rect 20242 39342 20244 39394
rect 20188 39330 20244 39342
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 38946 20244 38958
rect 20188 38894 20190 38946
rect 20242 38894 20244 38946
rect 20188 38164 20244 38894
rect 20300 38724 20356 40350
rect 20860 39842 20916 43596
rect 21532 43650 21588 43662
rect 21532 43598 21534 43650
rect 21586 43598 21588 43650
rect 21196 42980 21252 42990
rect 21196 42886 21252 42924
rect 21532 41972 21588 43598
rect 21980 42530 22036 42542
rect 21980 42478 21982 42530
rect 22034 42478 22036 42530
rect 21532 41906 21588 41916
rect 21756 42084 21812 42094
rect 20972 41860 21028 41870
rect 20972 40180 21028 41804
rect 21084 41076 21140 41086
rect 21084 40626 21140 41020
rect 21084 40574 21086 40626
rect 21138 40574 21140 40626
rect 21084 40562 21140 40574
rect 21756 40180 21812 42028
rect 21980 41300 22036 42478
rect 22092 42308 22148 44158
rect 23100 42868 23156 44382
rect 23100 42802 23156 42812
rect 22092 42242 22148 42252
rect 21980 41234 22036 41244
rect 23100 42194 23156 42206
rect 23100 42142 23102 42194
rect 23154 42142 23156 42194
rect 22876 40962 22932 40974
rect 22876 40910 22878 40962
rect 22930 40910 22932 40962
rect 22876 40628 22932 40910
rect 21868 40516 21924 40526
rect 22316 40516 22372 40526
rect 21868 40514 22260 40516
rect 21868 40462 21870 40514
rect 21922 40462 22260 40514
rect 21868 40460 22260 40462
rect 21868 40450 21924 40460
rect 20972 40124 21140 40180
rect 20860 39790 20862 39842
rect 20914 39790 20916 39842
rect 20860 39778 20916 39790
rect 20972 39396 21028 39406
rect 20972 39058 21028 39340
rect 20972 39006 20974 39058
rect 21026 39006 21028 39058
rect 20972 38994 21028 39006
rect 21084 39058 21140 40124
rect 21756 40114 21812 40124
rect 22204 39730 22260 40460
rect 22204 39678 22206 39730
rect 22258 39678 22260 39730
rect 22204 39666 22260 39678
rect 21308 39508 21364 39518
rect 21308 39414 21364 39452
rect 21644 39508 21700 39518
rect 22316 39508 22372 40460
rect 21084 39006 21086 39058
rect 21138 39006 21140 39058
rect 21084 38994 21140 39006
rect 20748 38948 20804 38958
rect 20804 38892 20916 38948
rect 20748 38882 20804 38892
rect 20300 38658 20356 38668
rect 20188 38108 20356 38164
rect 19516 37986 19572 37996
rect 19628 37940 19684 37950
rect 18956 36418 19012 36428
rect 19180 37492 19236 37502
rect 19180 35922 19236 37436
rect 19516 36372 19572 36382
rect 19516 36278 19572 36316
rect 19180 35870 19182 35922
rect 19234 35870 19236 35922
rect 19180 35858 19236 35870
rect 19628 35924 19684 37884
rect 19740 37938 19796 37950
rect 19740 37886 19742 37938
rect 19794 37886 19796 37938
rect 19740 37828 19796 37886
rect 20076 37940 20132 37950
rect 20076 37938 20244 37940
rect 20076 37886 20078 37938
rect 20130 37886 20244 37938
rect 20076 37884 20244 37886
rect 20076 37874 20132 37884
rect 19740 37762 19796 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19740 37492 19796 37502
rect 19740 36594 19796 37436
rect 20188 37490 20244 37884
rect 20188 37438 20190 37490
rect 20242 37438 20244 37490
rect 20188 37426 20244 37438
rect 20300 37268 20356 38108
rect 20636 38050 20692 38062
rect 20636 37998 20638 38050
rect 20690 37998 20692 38050
rect 20412 37940 20468 37950
rect 20412 37846 20468 37884
rect 20636 37828 20692 37998
rect 20636 37762 20692 37772
rect 20860 37492 20916 38892
rect 21308 38052 21364 38062
rect 20972 37492 21028 37502
rect 20860 37490 21028 37492
rect 20860 37438 20974 37490
rect 21026 37438 21028 37490
rect 20860 37436 21028 37438
rect 20972 37426 21028 37436
rect 19740 36542 19742 36594
rect 19794 36542 19796 36594
rect 19740 36530 19796 36542
rect 20076 37212 20356 37268
rect 21308 37266 21364 37996
rect 21308 37214 21310 37266
rect 21362 37214 21364 37266
rect 20076 36594 20132 37212
rect 21308 37202 21364 37214
rect 21532 37938 21588 37950
rect 21532 37886 21534 37938
rect 21586 37886 21588 37938
rect 20076 36542 20078 36594
rect 20130 36542 20132 36594
rect 20076 36530 20132 36542
rect 20412 36372 20468 36382
rect 20412 36278 20468 36316
rect 20748 36370 20804 36382
rect 20748 36318 20750 36370
rect 20802 36318 20804 36370
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35924 19796 35934
rect 19628 35922 19796 35924
rect 19628 35870 19742 35922
rect 19794 35870 19796 35922
rect 19628 35868 19796 35870
rect 19740 35858 19796 35868
rect 17388 35758 17390 35810
rect 17442 35758 17444 35810
rect 17388 35746 17444 35758
rect 17612 35812 17668 35822
rect 17612 35698 17668 35756
rect 18172 35812 18228 35822
rect 18172 35718 18228 35756
rect 17612 35646 17614 35698
rect 17666 35646 17668 35698
rect 17612 35634 17668 35646
rect 17164 34916 17220 35532
rect 18396 35586 18452 35598
rect 18396 35534 18398 35586
rect 18450 35534 18452 35586
rect 18396 35364 18452 35534
rect 18956 35588 19012 35598
rect 18956 35494 19012 35532
rect 18396 35298 18452 35308
rect 17164 34822 17220 34860
rect 17724 34916 17780 34926
rect 17724 34822 17780 34860
rect 16492 34638 16494 34690
rect 16546 34638 16548 34690
rect 16492 34626 16548 34638
rect 20188 34690 20244 34702
rect 20188 34638 20190 34690
rect 20242 34638 20244 34690
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 17836 34356 17892 34366
rect 20188 34356 20244 34638
rect 17276 34132 17332 34142
rect 17164 34130 17332 34132
rect 17164 34078 17278 34130
rect 17330 34078 17332 34130
rect 17164 34076 17332 34078
rect 16268 34020 16324 34030
rect 16492 34020 16548 34030
rect 16268 33926 16324 33964
rect 16380 34018 16548 34020
rect 16380 33966 16494 34018
rect 16546 33966 16548 34018
rect 16380 33964 16548 33966
rect 15932 33518 15934 33570
rect 15986 33518 15988 33570
rect 15932 33506 15988 33518
rect 16156 33124 16212 33134
rect 16156 32786 16212 33068
rect 16156 32734 16158 32786
rect 16210 32734 16212 32786
rect 16156 32722 16212 32734
rect 15036 30322 15092 32396
rect 15036 30270 15038 30322
rect 15090 30270 15092 30322
rect 12012 30210 12180 30212
rect 12012 30158 12014 30210
rect 12066 30158 12180 30210
rect 12012 30156 12180 30158
rect 12012 30146 12068 30156
rect 10108 29596 10276 29652
rect 9100 29428 9156 29438
rect 9100 29334 9156 29372
rect 9660 29428 9716 29438
rect 9660 29334 9716 29372
rect 10108 29426 10164 29438
rect 10108 29374 10110 29426
rect 10162 29374 10164 29426
rect 8876 28478 8878 28530
rect 8930 28478 8932 28530
rect 8876 28466 8932 28478
rect 9884 28644 9940 28654
rect 9884 27860 9940 28588
rect 9884 27766 9940 27804
rect 9548 27748 9604 27758
rect 9324 27746 9604 27748
rect 9324 27694 9550 27746
rect 9602 27694 9604 27746
rect 9324 27692 9604 27694
rect 8764 26350 8766 26402
rect 8818 26350 8820 26402
rect 8764 26338 8820 26350
rect 9100 27634 9156 27646
rect 9100 27582 9102 27634
rect 9154 27582 9156 27634
rect 9100 26068 9156 27582
rect 9100 26002 9156 26012
rect 9324 25732 9380 27692
rect 9548 27682 9604 27692
rect 10108 27188 10164 29374
rect 10220 28308 10276 29596
rect 11564 29428 11620 29438
rect 10220 28242 10276 28252
rect 11116 28642 11172 28654
rect 11116 28590 11118 28642
rect 11170 28590 11172 28642
rect 10556 27972 10612 27982
rect 10556 27878 10612 27916
rect 10892 27860 10948 27870
rect 10892 27766 10948 27804
rect 11116 27300 11172 28590
rect 11564 28642 11620 29372
rect 12124 28756 12180 30156
rect 12348 30146 12404 30156
rect 13692 30212 13748 30222
rect 13692 30118 13748 30156
rect 14028 30212 14084 30222
rect 12236 30098 12292 30110
rect 12236 30046 12238 30098
rect 12290 30046 12292 30098
rect 12236 29988 12292 30046
rect 12348 29988 12404 29998
rect 12236 29932 12348 29988
rect 12348 29922 12404 29932
rect 14028 29988 14084 30156
rect 15036 30212 15092 30270
rect 15036 30146 15092 30156
rect 15372 32674 15428 32686
rect 15372 32622 15374 32674
rect 15426 32622 15428 32674
rect 15372 30210 15428 32622
rect 16380 31218 16436 33964
rect 16492 33954 16548 33964
rect 16828 34018 16884 34030
rect 16828 33966 16830 34018
rect 16882 33966 16884 34018
rect 16716 33346 16772 33358
rect 16716 33294 16718 33346
rect 16770 33294 16772 33346
rect 16716 32564 16772 33294
rect 16492 32450 16548 32462
rect 16492 32398 16494 32450
rect 16546 32398 16548 32450
rect 16492 31554 16548 32398
rect 16492 31502 16494 31554
rect 16546 31502 16548 31554
rect 16492 31490 16548 31502
rect 16380 31166 16382 31218
rect 16434 31166 16436 31218
rect 16380 31154 16436 31166
rect 15372 30158 15374 30210
rect 15426 30158 15428 30210
rect 15372 30146 15428 30158
rect 16380 30884 16436 30894
rect 16380 30098 16436 30828
rect 16380 30046 16382 30098
rect 16434 30046 16436 30098
rect 16380 30034 16436 30046
rect 16716 30660 16772 32508
rect 16828 32452 16884 33966
rect 17164 33346 17220 34076
rect 17276 34066 17332 34076
rect 17836 34130 17892 34300
rect 17836 34078 17838 34130
rect 17890 34078 17892 34130
rect 17836 34066 17892 34078
rect 20076 34300 20244 34356
rect 20412 34354 20468 34366
rect 20412 34302 20414 34354
rect 20466 34302 20468 34354
rect 17164 33294 17166 33346
rect 17218 33294 17220 33346
rect 16828 32358 16884 32396
rect 17052 33012 17108 33022
rect 17052 31890 17108 32956
rect 17052 31838 17054 31890
rect 17106 31838 17108 31890
rect 17052 31826 17108 31838
rect 17164 31778 17220 33294
rect 17724 33346 17780 33358
rect 17724 33294 17726 33346
rect 17778 33294 17780 33346
rect 17164 31726 17166 31778
rect 17218 31726 17220 31778
rect 16940 31108 16996 31118
rect 16940 31014 16996 31052
rect 14028 29922 14084 29932
rect 15596 29986 15652 29998
rect 15596 29934 15598 29986
rect 15650 29934 15652 29986
rect 13244 29764 13300 29774
rect 12572 29652 12628 29662
rect 12572 29650 12740 29652
rect 12572 29598 12574 29650
rect 12626 29598 12740 29650
rect 12572 29596 12740 29598
rect 12572 29586 12628 29596
rect 12236 28756 12292 28766
rect 12124 28754 12628 28756
rect 12124 28702 12238 28754
rect 12290 28702 12628 28754
rect 12124 28700 12628 28702
rect 12236 28690 12292 28700
rect 11564 28590 11566 28642
rect 11618 28590 11620 28642
rect 11452 28532 11508 28542
rect 11452 27860 11508 28476
rect 11452 27766 11508 27804
rect 11116 27234 11172 27244
rect 10108 27122 10164 27132
rect 11564 26852 11620 28590
rect 12572 28532 12628 28700
rect 12684 28754 12740 29596
rect 13244 29650 13300 29708
rect 13244 29598 13246 29650
rect 13298 29598 13300 29650
rect 13244 29586 13300 29598
rect 14028 29538 14084 29550
rect 14028 29486 14030 29538
rect 14082 29486 14084 29538
rect 13132 29202 13188 29214
rect 13132 29150 13134 29202
rect 13186 29150 13188 29202
rect 12684 28702 12686 28754
rect 12738 28702 12740 28754
rect 12684 28690 12740 28702
rect 12908 28756 12964 28766
rect 12908 28662 12964 28700
rect 12572 28476 12852 28532
rect 12684 27972 12740 27982
rect 12684 27878 12740 27916
rect 11676 27746 11732 27758
rect 11676 27694 11678 27746
rect 11730 27694 11732 27746
rect 11676 27300 11732 27694
rect 11900 27636 11956 27646
rect 11900 27542 11956 27580
rect 11676 27244 11844 27300
rect 9772 26292 9828 26302
rect 9772 26198 9828 26236
rect 10892 26292 10948 26302
rect 9548 26180 9604 26190
rect 9324 25666 9380 25676
rect 9436 26178 9604 26180
rect 9436 26126 9550 26178
rect 9602 26126 9604 26178
rect 9436 26124 9604 26126
rect 8764 25620 8820 25630
rect 8316 25618 9044 25620
rect 8316 25566 8318 25618
rect 8370 25566 8766 25618
rect 8818 25566 9044 25618
rect 8316 25564 9044 25566
rect 8316 25554 8372 25564
rect 8316 25396 8372 25406
rect 8316 24946 8372 25340
rect 8316 24894 8318 24946
rect 8370 24894 8372 24946
rect 8316 24882 8372 24894
rect 8316 24612 8372 24622
rect 8316 23378 8372 24556
rect 8316 23326 8318 23378
rect 8370 23326 8372 23378
rect 8316 23314 8372 23326
rect 8204 21410 8260 21420
rect 8316 21698 8372 21710
rect 8316 21646 8318 21698
rect 8370 21646 8372 21698
rect 7980 20804 8036 20814
rect 7980 20710 8036 20748
rect 8316 20130 8372 21646
rect 8428 20804 8484 25564
rect 8764 25554 8820 25564
rect 8988 25508 9044 25564
rect 8988 25414 9044 25452
rect 9436 25396 9492 26124
rect 9548 26114 9604 26124
rect 10332 26178 10388 26190
rect 10332 26126 10334 26178
rect 10386 26126 10388 26178
rect 9436 25330 9492 25340
rect 9548 25506 9604 25518
rect 9548 25454 9550 25506
rect 9602 25454 9604 25506
rect 9548 25284 9604 25454
rect 10220 25508 10276 25518
rect 10332 25508 10388 26126
rect 10276 25452 10388 25508
rect 10668 26178 10724 26190
rect 10668 26126 10670 26178
rect 10722 26126 10724 26178
rect 9772 25284 9828 25294
rect 9548 25218 9604 25228
rect 9660 25228 9772 25284
rect 9436 24724 9492 24734
rect 9324 24722 9492 24724
rect 9324 24670 9438 24722
rect 9490 24670 9492 24722
rect 9324 24668 9492 24670
rect 9100 24500 9156 24510
rect 8988 24498 9156 24500
rect 8988 24446 9102 24498
rect 9154 24446 9156 24498
rect 8988 24444 9156 24446
rect 8652 22148 8708 22158
rect 8652 22146 8820 22148
rect 8652 22094 8654 22146
rect 8706 22094 8820 22146
rect 8652 22092 8820 22094
rect 8652 22082 8708 22092
rect 8652 21924 8708 21934
rect 8652 20914 8708 21868
rect 8652 20862 8654 20914
rect 8706 20862 8708 20914
rect 8652 20850 8708 20862
rect 8428 20710 8484 20748
rect 8316 20078 8318 20130
rect 8370 20078 8372 20130
rect 8316 20066 8372 20078
rect 7980 19908 8036 19918
rect 7980 19814 8036 19852
rect 8764 19906 8820 22092
rect 8988 21588 9044 24444
rect 9100 24434 9156 24444
rect 9324 23604 9380 24668
rect 9436 24658 9492 24668
rect 9100 22930 9156 22942
rect 9100 22878 9102 22930
rect 9154 22878 9156 22930
rect 9100 21588 9156 22878
rect 9324 22370 9380 23548
rect 9660 23156 9716 25228
rect 9772 25218 9828 25228
rect 10108 24722 10164 24734
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 9548 23100 9716 23156
rect 9772 23938 9828 23950
rect 9772 23886 9774 23938
rect 9826 23886 9828 23938
rect 9324 22318 9326 22370
rect 9378 22318 9380 22370
rect 9212 22148 9268 22158
rect 9212 22054 9268 22092
rect 9212 21812 9268 21822
rect 9324 21812 9380 22318
rect 9268 21756 9380 21812
rect 9436 22930 9492 22942
rect 9436 22878 9438 22930
rect 9490 22878 9492 22930
rect 9436 21812 9492 22878
rect 9212 21746 9268 21756
rect 9436 21746 9492 21756
rect 9100 21532 9268 21588
rect 8988 21522 9044 21532
rect 9100 21362 9156 21374
rect 9100 21310 9102 21362
rect 9154 21310 9156 21362
rect 8764 19854 8766 19906
rect 8818 19854 8820 19906
rect 8764 19842 8820 19854
rect 8988 19908 9044 19918
rect 8988 19814 9044 19852
rect 8316 19348 8372 19358
rect 8316 19254 8372 19292
rect 7868 18286 7870 18338
rect 7922 18286 7924 18338
rect 7868 18274 7924 18286
rect 6188 17714 6244 17724
rect 8652 17780 8708 17790
rect 8652 17686 8708 17724
rect 9100 17556 9156 21310
rect 9212 20356 9268 21532
rect 9212 20290 9268 20300
rect 9436 21362 9492 21374
rect 9436 21310 9438 21362
rect 9490 21310 9492 21362
rect 9436 18116 9492 21310
rect 9548 19122 9604 23100
rect 9772 22036 9828 23886
rect 10108 23380 10164 24670
rect 10220 23938 10276 25452
rect 10668 24612 10724 26126
rect 10668 24546 10724 24556
rect 10220 23886 10222 23938
rect 10274 23886 10276 23938
rect 10220 23874 10276 23886
rect 10892 23940 10948 26236
rect 11452 26180 11508 26190
rect 11564 26180 11620 26796
rect 11676 27074 11732 27086
rect 11676 27022 11678 27074
rect 11730 27022 11732 27074
rect 11676 26516 11732 27022
rect 11788 26516 11844 27244
rect 12796 27186 12852 28476
rect 12796 27134 12798 27186
rect 12850 27134 12852 27186
rect 12796 27122 12852 27134
rect 11788 26460 12068 26516
rect 11676 26450 11732 26460
rect 11900 26180 11956 26190
rect 11452 26178 11956 26180
rect 11452 26126 11454 26178
rect 11506 26126 11902 26178
rect 11954 26126 11956 26178
rect 11452 26124 11956 26126
rect 11452 25508 11508 26124
rect 11900 26114 11956 26124
rect 11452 24050 11508 25452
rect 12012 25282 12068 26460
rect 12012 25230 12014 25282
rect 12066 25230 12068 25282
rect 12012 25218 12068 25230
rect 12124 26290 12180 26302
rect 12124 26238 12126 26290
rect 12178 26238 12180 26290
rect 11452 23998 11454 24050
rect 11506 23998 11508 24050
rect 11452 23986 11508 23998
rect 10892 23846 10948 23884
rect 11900 23940 11956 23950
rect 11900 23846 11956 23884
rect 10668 23828 10724 23838
rect 10332 23826 10724 23828
rect 10332 23774 10670 23826
rect 10722 23774 10724 23826
rect 10332 23772 10724 23774
rect 10108 23314 10164 23324
rect 10220 23716 10276 23726
rect 10220 23378 10276 23660
rect 10220 23326 10222 23378
rect 10274 23326 10276 23378
rect 10220 23314 10276 23326
rect 9772 21970 9828 21980
rect 9996 22370 10052 22382
rect 9996 22318 9998 22370
rect 10050 22318 10052 22370
rect 9660 21476 9716 21486
rect 9660 20690 9716 21420
rect 9660 20638 9662 20690
rect 9714 20638 9716 20690
rect 9660 20626 9716 20638
rect 9884 21140 9940 21150
rect 9660 20356 9716 20366
rect 9660 20244 9716 20300
rect 9660 20188 9828 20244
rect 9548 19070 9550 19122
rect 9602 19070 9604 19122
rect 9548 19058 9604 19070
rect 9772 18564 9828 20188
rect 9884 20130 9940 21084
rect 9884 20078 9886 20130
rect 9938 20078 9940 20130
rect 9884 20066 9940 20078
rect 9884 18564 9940 18574
rect 9772 18562 9940 18564
rect 9772 18510 9886 18562
rect 9938 18510 9940 18562
rect 9772 18508 9940 18510
rect 9884 18498 9940 18508
rect 9436 18060 9828 18116
rect 9660 17556 9716 17566
rect 9100 17554 9716 17556
rect 9100 17502 9662 17554
rect 9714 17502 9716 17554
rect 9100 17500 9716 17502
rect 9660 17490 9716 17500
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 9772 15988 9828 18060
rect 9996 16210 10052 22318
rect 10220 21812 10276 21822
rect 10332 21812 10388 23772
rect 10668 23762 10724 23772
rect 12124 23604 12180 26238
rect 12684 26290 12740 26302
rect 12684 26238 12686 26290
rect 12738 26238 12740 26290
rect 12684 25620 12740 26238
rect 12684 25554 12740 25564
rect 12684 25282 12740 25294
rect 12684 25230 12686 25282
rect 12738 25230 12740 25282
rect 12348 24836 12404 24846
rect 12236 24834 12404 24836
rect 12236 24782 12350 24834
rect 12402 24782 12404 24834
rect 12236 24780 12404 24782
rect 12236 24050 12292 24780
rect 12348 24770 12404 24780
rect 12684 24836 12740 25230
rect 12684 24770 12740 24780
rect 13132 24724 13188 29150
rect 13916 28756 13972 28766
rect 13804 28642 13860 28654
rect 13804 28590 13806 28642
rect 13858 28590 13860 28642
rect 13692 27972 13748 27982
rect 13692 27186 13748 27916
rect 13692 27134 13694 27186
rect 13746 27134 13748 27186
rect 13692 27122 13748 27134
rect 13804 27076 13860 28590
rect 13804 27010 13860 27020
rect 13916 27074 13972 28700
rect 14028 28084 14084 29486
rect 15596 29316 15652 29934
rect 16380 29428 16436 29438
rect 16380 29426 16660 29428
rect 16380 29374 16382 29426
rect 16434 29374 16660 29426
rect 16380 29372 16660 29374
rect 16380 29362 16436 29372
rect 15596 29250 15652 29260
rect 15708 28756 15764 28766
rect 15708 28662 15764 28700
rect 16380 28756 16436 28766
rect 16380 28662 16436 28700
rect 14028 28018 14084 28028
rect 15036 28420 15092 28430
rect 14924 27858 14980 27870
rect 14924 27806 14926 27858
rect 14978 27806 14980 27858
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 27010 13972 27022
rect 14812 27076 14868 27086
rect 14812 26982 14868 27020
rect 14700 26964 14756 26974
rect 13580 26516 13636 26526
rect 13580 25618 13636 26460
rect 13580 25566 13582 25618
rect 13634 25566 13636 25618
rect 13580 25554 13636 25566
rect 14700 25618 14756 26908
rect 14700 25566 14702 25618
rect 14754 25566 14756 25618
rect 14700 25554 14756 25566
rect 14924 25620 14980 27806
rect 15036 26514 15092 28364
rect 16492 28420 16548 28430
rect 16492 28326 16548 28364
rect 15596 27858 15652 27870
rect 15596 27806 15598 27858
rect 15650 27806 15652 27858
rect 15372 27186 15428 27198
rect 15372 27134 15374 27186
rect 15426 27134 15428 27186
rect 15372 26964 15428 27134
rect 15372 26898 15428 26908
rect 15596 26852 15652 27806
rect 15932 27746 15988 27758
rect 15932 27694 15934 27746
rect 15986 27694 15988 27746
rect 15932 27634 15988 27694
rect 15932 27582 15934 27634
rect 15986 27582 15988 27634
rect 15932 27076 15988 27582
rect 15932 27010 15988 27020
rect 16380 27748 16436 27758
rect 16380 26964 16436 27692
rect 16380 26898 16436 26908
rect 16604 26908 16660 29372
rect 16716 27636 16772 30604
rect 16828 30324 16884 30334
rect 17164 30324 17220 31726
rect 16884 30268 17220 30324
rect 17276 32564 17332 32574
rect 16828 29652 16884 30268
rect 16828 29426 16884 29596
rect 16828 29374 16830 29426
rect 16882 29374 16884 29426
rect 16828 28644 16884 29374
rect 17164 28644 17220 28654
rect 16828 28642 17220 28644
rect 16828 28590 17166 28642
rect 17218 28590 17220 28642
rect 16828 28588 17220 28590
rect 16828 28082 16884 28588
rect 17164 28578 17220 28588
rect 16828 28030 16830 28082
rect 16882 28030 16884 28082
rect 16828 28018 16884 28030
rect 16716 27634 16884 27636
rect 16716 27582 16718 27634
rect 16770 27582 16884 27634
rect 16716 27580 16884 27582
rect 16716 27570 16772 27580
rect 16604 26852 16772 26908
rect 15596 26786 15652 26796
rect 15036 26462 15038 26514
rect 15090 26462 15092 26514
rect 15036 26450 15092 26462
rect 16380 26516 16436 26526
rect 16380 26178 16436 26460
rect 16380 26126 16382 26178
rect 16434 26126 16436 26178
rect 15484 26068 15540 26078
rect 14924 25564 15092 25620
rect 14924 25396 14980 25406
rect 14812 25394 14980 25396
rect 14812 25342 14926 25394
rect 14978 25342 14980 25394
rect 14812 25340 14980 25342
rect 13356 24724 13412 24734
rect 13132 24668 13300 24724
rect 13132 24500 13188 24510
rect 12236 23998 12238 24050
rect 12290 23998 12292 24050
rect 12236 23986 12292 23998
rect 12796 24498 13188 24500
rect 12796 24446 13134 24498
rect 13186 24446 13188 24498
rect 12796 24444 13188 24446
rect 12684 23940 12740 23950
rect 12572 23826 12628 23838
rect 12572 23774 12574 23826
rect 12626 23774 12628 23826
rect 12572 23716 12628 23774
rect 12572 23650 12628 23660
rect 12124 23538 12180 23548
rect 10892 23380 10948 23390
rect 10948 23324 11172 23380
rect 10892 23314 10948 23324
rect 10892 22932 10948 22942
rect 10780 22148 10836 22158
rect 10220 21810 10388 21812
rect 10220 21758 10222 21810
rect 10274 21758 10388 21810
rect 10220 21756 10388 21758
rect 10556 21812 10612 21822
rect 10220 21746 10276 21756
rect 10556 19122 10612 21756
rect 10556 19070 10558 19122
rect 10610 19070 10612 19122
rect 10556 19058 10612 19070
rect 10780 17554 10836 22092
rect 10892 20690 10948 22876
rect 10892 20638 10894 20690
rect 10946 20638 10948 20690
rect 10892 20626 10948 20638
rect 11004 21700 11060 21710
rect 11004 19906 11060 21644
rect 11004 19854 11006 19906
rect 11058 19854 11060 19906
rect 11004 19842 11060 19854
rect 11116 18338 11172 23324
rect 12572 23154 12628 23166
rect 12572 23102 12574 23154
rect 12626 23102 12628 23154
rect 12460 22146 12516 22158
rect 12460 22094 12462 22146
rect 12514 22094 12516 22146
rect 11900 21924 11956 21934
rect 11788 21868 11900 21924
rect 11788 20914 11844 21868
rect 11900 21858 11956 21868
rect 12460 21812 12516 22094
rect 12572 22036 12628 23102
rect 12572 21970 12628 21980
rect 12460 21746 12516 21756
rect 12460 21588 12516 21598
rect 11788 20862 11790 20914
rect 11842 20862 11844 20914
rect 11788 20850 11844 20862
rect 11900 21586 12516 21588
rect 11900 21534 12462 21586
rect 12514 21534 12516 21586
rect 11900 21532 12516 21534
rect 11788 20692 11844 20702
rect 11788 19346 11844 20636
rect 11788 19294 11790 19346
rect 11842 19294 11844 19346
rect 11788 19282 11844 19294
rect 11116 18286 11118 18338
rect 11170 18286 11172 18338
rect 11116 18274 11172 18286
rect 11340 18452 11396 18462
rect 10780 17502 10782 17554
rect 10834 17502 10836 17554
rect 10780 17490 10836 17502
rect 11340 16770 11396 18396
rect 11900 17778 11956 21532
rect 12460 21522 12516 21532
rect 12684 20916 12740 23884
rect 12684 20356 12740 20860
rect 12684 20290 12740 20300
rect 11900 17726 11902 17778
rect 11954 17726 11956 17778
rect 11900 17714 11956 17726
rect 12684 16996 12740 17006
rect 12796 16996 12852 24444
rect 13132 24434 13188 24444
rect 12908 23940 12964 23950
rect 12908 23846 12964 23884
rect 12908 23604 12964 23614
rect 12908 23154 12964 23548
rect 13244 23380 13300 24668
rect 13356 23828 13412 24668
rect 13804 24722 13860 24734
rect 13804 24670 13806 24722
rect 13858 24670 13860 24722
rect 13692 23828 13748 23838
rect 13356 23826 13748 23828
rect 13356 23774 13694 23826
rect 13746 23774 13748 23826
rect 13356 23772 13748 23774
rect 13356 23604 13412 23772
rect 13692 23762 13748 23772
rect 13356 23538 13412 23548
rect 13244 23324 13412 23380
rect 12908 23102 12910 23154
rect 12962 23102 12964 23154
rect 12908 22372 12964 23102
rect 13244 22932 13300 22942
rect 13244 22838 13300 22876
rect 12908 22316 13300 22372
rect 12908 21586 12964 22316
rect 12908 21534 12910 21586
rect 12962 21534 12964 21586
rect 12908 21522 12964 21534
rect 13020 22146 13076 22158
rect 13020 22094 13022 22146
rect 13074 22094 13076 22146
rect 13020 21140 13076 22094
rect 13244 21586 13300 22316
rect 13244 21534 13246 21586
rect 13298 21534 13300 21586
rect 13244 21522 13300 21534
rect 13020 21074 13076 21084
rect 13356 18562 13412 23324
rect 13580 22372 13636 22382
rect 13580 22278 13636 22316
rect 13804 22260 13860 24670
rect 14812 24276 14868 25340
rect 14924 25330 14980 25340
rect 14028 24220 14868 24276
rect 14028 23378 14084 24220
rect 14028 23326 14030 23378
rect 14082 23326 14084 23378
rect 14028 23314 14084 23326
rect 13692 22204 13860 22260
rect 13916 22370 13972 22382
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 13468 20916 13524 20926
rect 13468 20130 13524 20860
rect 13692 20692 13748 22204
rect 13916 21924 13972 22318
rect 13916 21858 13972 21868
rect 13804 21812 13860 21822
rect 13804 20914 13860 21756
rect 13804 20862 13806 20914
rect 13858 20862 13860 20914
rect 13804 20850 13860 20862
rect 13916 21586 13972 21598
rect 13916 21534 13918 21586
rect 13970 21534 13972 21586
rect 13692 20626 13748 20636
rect 13468 20078 13470 20130
rect 13522 20078 13524 20130
rect 13468 20066 13524 20078
rect 13356 18510 13358 18562
rect 13410 18510 13412 18562
rect 13356 18498 13412 18510
rect 12684 16994 12852 16996
rect 12684 16942 12686 16994
rect 12738 16942 12852 16994
rect 12684 16940 12852 16942
rect 12684 16930 12740 16940
rect 11340 16718 11342 16770
rect 11394 16718 11396 16770
rect 11340 16706 11396 16718
rect 9996 16158 9998 16210
rect 10050 16158 10052 16210
rect 9996 16146 10052 16158
rect 13916 16212 13972 21534
rect 15036 20188 15092 25564
rect 15260 25394 15316 25406
rect 15260 25342 15262 25394
rect 15314 25342 15316 25394
rect 15260 20916 15316 25342
rect 15260 20822 15316 20860
rect 15484 20692 15540 26012
rect 15820 26066 15876 26078
rect 15820 26014 15822 26066
rect 15874 26014 15876 26066
rect 15708 25506 15764 25518
rect 15708 25454 15710 25506
rect 15762 25454 15764 25506
rect 15708 24500 15764 25454
rect 15820 25284 15876 26014
rect 16380 25844 16436 26126
rect 16380 25778 16436 25788
rect 16156 25508 16212 25518
rect 16156 25506 16660 25508
rect 16156 25454 16158 25506
rect 16210 25454 16660 25506
rect 16156 25452 16660 25454
rect 16156 25442 16212 25452
rect 15820 25218 15876 25228
rect 15708 24434 15764 24444
rect 16380 24946 16436 24958
rect 16380 24894 16382 24946
rect 16434 24894 16436 24946
rect 16380 24052 16436 24894
rect 16380 23986 16436 23996
rect 16268 23154 16324 23166
rect 16268 23102 16270 23154
rect 16322 23102 16324 23154
rect 15820 22372 15876 22382
rect 15596 21252 15652 21262
rect 15596 20914 15652 21196
rect 15596 20862 15598 20914
rect 15650 20862 15652 20914
rect 15596 20850 15652 20862
rect 15708 20804 15764 20814
rect 15484 20636 15652 20692
rect 14476 20132 15092 20188
rect 14476 18338 14532 20132
rect 14924 20018 14980 20030
rect 14924 19966 14926 20018
rect 14978 19966 14980 20018
rect 14924 19684 14980 19966
rect 15484 19908 15540 19918
rect 15484 19814 15540 19852
rect 14924 19618 14980 19628
rect 15596 19122 15652 20636
rect 15596 19070 15598 19122
rect 15650 19070 15652 19122
rect 15596 19058 15652 19070
rect 14476 18286 14478 18338
rect 14530 18286 14532 18338
rect 14476 18274 14532 18286
rect 15596 16772 15652 16782
rect 15708 16772 15764 20748
rect 15820 20802 15876 22316
rect 16156 21698 16212 21710
rect 16156 21646 16158 21698
rect 16210 21646 16212 21698
rect 16156 21252 16212 21646
rect 16268 21700 16324 23102
rect 16268 21634 16324 21644
rect 16380 22148 16436 22158
rect 16156 21186 16212 21196
rect 16380 21028 16436 22092
rect 15820 20750 15822 20802
rect 15874 20750 15876 20802
rect 15820 20738 15876 20750
rect 16156 20972 16436 21028
rect 16492 22146 16548 22158
rect 16492 22094 16494 22146
rect 16546 22094 16548 22146
rect 15596 16770 15764 16772
rect 15596 16718 15598 16770
rect 15650 16718 15764 16770
rect 15596 16716 15764 16718
rect 15596 16706 15652 16716
rect 14812 16212 14868 16222
rect 13916 16210 14868 16212
rect 13916 16158 14814 16210
rect 14866 16158 14868 16210
rect 13916 16156 14868 16158
rect 14812 16146 14868 16156
rect 9884 15988 9940 15998
rect 9772 15932 9884 15988
rect 9884 15922 9940 15932
rect 10892 15988 10948 15998
rect 10892 15894 10948 15932
rect 16156 15986 16212 20972
rect 16380 20804 16436 20842
rect 16380 20738 16436 20748
rect 16380 20580 16436 20590
rect 16380 18340 16436 20524
rect 16492 20130 16548 22094
rect 16492 20078 16494 20130
rect 16546 20078 16548 20130
rect 16492 20066 16548 20078
rect 16492 18340 16548 18350
rect 16380 18284 16492 18340
rect 16492 18274 16548 18284
rect 16604 17778 16660 25452
rect 16716 21140 16772 26852
rect 16828 26178 16884 27580
rect 17276 26908 17332 32508
rect 17612 32452 17668 32462
rect 17612 31108 17668 32396
rect 17724 32228 17780 33294
rect 20076 33348 20132 34300
rect 20412 33460 20468 34302
rect 20748 34132 20804 36318
rect 21532 35252 21588 37886
rect 21644 37828 21700 39452
rect 21868 39452 22372 39508
rect 22428 39618 22484 39630
rect 22428 39566 22430 39618
rect 22482 39566 22484 39618
rect 22428 39508 22484 39566
rect 21868 39058 21924 39452
rect 22428 39442 22484 39452
rect 22876 39508 22932 40572
rect 23100 39730 23156 42142
rect 23660 41860 23716 44828
rect 23772 43538 23828 46284
rect 23884 43708 23940 46620
rect 23996 43876 24052 49868
rect 24332 49026 24388 49038
rect 24332 48974 24334 49026
rect 24386 48974 24388 49026
rect 24220 48580 24276 48590
rect 24220 45666 24276 48524
rect 24332 47572 24388 48974
rect 24332 47506 24388 47516
rect 24444 46676 24500 51436
rect 27132 51268 27188 51278
rect 26908 51266 27188 51268
rect 26908 51214 27134 51266
rect 27186 51214 27188 51266
rect 26908 51212 27188 51214
rect 24556 50708 24612 50718
rect 24556 50706 24836 50708
rect 24556 50654 24558 50706
rect 24610 50654 24836 50706
rect 24556 50652 24836 50654
rect 24556 50642 24612 50652
rect 24780 49026 24836 50652
rect 25340 50482 25396 50494
rect 25340 50430 25342 50482
rect 25394 50430 25396 50482
rect 24780 48974 24782 49026
rect 24834 48974 24836 49026
rect 24780 48962 24836 48974
rect 25228 49698 25284 49710
rect 25228 49646 25230 49698
rect 25282 49646 25284 49698
rect 25228 48580 25284 49646
rect 25228 48514 25284 48524
rect 25340 48356 25396 50430
rect 26572 50482 26628 50494
rect 26572 50430 26574 50482
rect 26626 50430 26628 50482
rect 24892 48300 25396 48356
rect 25452 49810 25508 49822
rect 25452 49758 25454 49810
rect 25506 49758 25508 49810
rect 25452 49700 25508 49758
rect 24668 47348 24724 47358
rect 24668 47254 24724 47292
rect 24444 46620 24612 46676
rect 24444 46452 24500 46462
rect 24444 46358 24500 46396
rect 24220 45614 24222 45666
rect 24274 45614 24276 45666
rect 24220 45602 24276 45614
rect 24332 45668 24388 45678
rect 24108 44884 24164 44894
rect 24108 44434 24164 44828
rect 24108 44382 24110 44434
rect 24162 44382 24164 44434
rect 24108 44370 24164 44382
rect 24220 43876 24276 43886
rect 23996 43820 24220 43876
rect 24220 43810 24276 43820
rect 23884 43652 24276 43708
rect 23772 43486 23774 43538
rect 23826 43486 23828 43538
rect 23772 43474 23828 43486
rect 24220 42754 24276 43652
rect 24220 42702 24222 42754
rect 24274 42702 24276 42754
rect 24220 42690 24276 42702
rect 23772 42644 23828 42654
rect 23772 41970 23828 42588
rect 24332 42084 24388 45612
rect 24444 45332 24500 45342
rect 24556 45332 24612 46620
rect 24892 46114 24948 48300
rect 25340 48132 25396 48142
rect 25452 48132 25508 49644
rect 25676 49812 25732 49822
rect 25676 49476 25732 49756
rect 26124 49700 26180 49710
rect 26124 49606 26180 49644
rect 25340 48130 25508 48132
rect 25340 48078 25342 48130
rect 25394 48078 25508 48130
rect 25340 48076 25508 48078
rect 25564 49420 25732 49476
rect 25340 48020 25396 48076
rect 24892 46062 24894 46114
rect 24946 46062 24948 46114
rect 24892 46050 24948 46062
rect 25116 47572 25172 47582
rect 25116 47458 25172 47516
rect 25116 47406 25118 47458
rect 25170 47406 25172 47458
rect 25116 46676 25172 47406
rect 25340 47460 25396 47964
rect 25340 47394 25396 47404
rect 25564 47458 25620 49420
rect 26572 48916 26628 50430
rect 26572 48850 26628 48860
rect 25900 48242 25956 48254
rect 25900 48190 25902 48242
rect 25954 48190 25956 48242
rect 25676 48132 25732 48142
rect 25676 48038 25732 48076
rect 25900 48020 25956 48190
rect 25900 47954 25956 47964
rect 26460 48242 26516 48254
rect 26460 48190 26462 48242
rect 26514 48190 26516 48242
rect 25564 47406 25566 47458
rect 25618 47406 25620 47458
rect 25564 47394 25620 47406
rect 24444 45330 24612 45332
rect 24444 45278 24446 45330
rect 24498 45278 24612 45330
rect 24444 45276 24612 45278
rect 25116 45892 25172 46620
rect 24444 45266 24500 45276
rect 24892 44996 24948 45006
rect 24556 44322 24612 44334
rect 24556 44270 24558 44322
rect 24610 44270 24612 44322
rect 24556 44100 24612 44270
rect 24892 44322 24948 44940
rect 24892 44270 24894 44322
rect 24946 44270 24948 44322
rect 24892 44258 24948 44270
rect 25116 44100 25172 45836
rect 25564 47012 25620 47022
rect 25564 45890 25620 46956
rect 25564 45838 25566 45890
rect 25618 45838 25620 45890
rect 25564 45826 25620 45838
rect 25676 46786 25732 46798
rect 25676 46734 25678 46786
rect 25730 46734 25732 46786
rect 25676 45220 25732 46734
rect 26460 46676 26516 48190
rect 26908 48242 26964 51212
rect 27132 51202 27188 51212
rect 27244 49812 27300 52222
rect 28140 52052 28196 52062
rect 28028 52050 28196 52052
rect 28028 51998 28142 52050
rect 28194 51998 28196 52050
rect 28028 51996 28196 51998
rect 27916 51492 27972 51502
rect 27804 51436 27916 51492
rect 27580 50708 27636 50718
rect 27580 50706 27748 50708
rect 27580 50654 27582 50706
rect 27634 50654 27748 50706
rect 27580 50652 27748 50654
rect 27580 50642 27636 50652
rect 27692 50428 27748 50652
rect 27244 49746 27300 49756
rect 27580 50372 27748 50428
rect 27356 48804 27412 48814
rect 27356 48710 27412 48748
rect 26908 48190 26910 48242
rect 26962 48190 26964 48242
rect 26908 48178 26964 48190
rect 27132 47348 27188 47358
rect 27188 47292 27300 47348
rect 27132 47282 27188 47292
rect 26460 46610 26516 46620
rect 25676 45154 25732 45164
rect 26572 46562 26628 46574
rect 26572 46510 26574 46562
rect 26626 46510 26628 46562
rect 24556 44044 25172 44100
rect 24556 43708 24612 44044
rect 24444 43652 24612 43708
rect 24780 43876 24836 43886
rect 24444 43538 24500 43652
rect 24444 43486 24446 43538
rect 24498 43486 24500 43538
rect 24444 43474 24500 43486
rect 24780 42532 24836 43820
rect 25116 43708 25172 44044
rect 24892 43652 25172 43708
rect 25788 44100 25844 44110
rect 24892 42754 24948 43652
rect 24892 42702 24894 42754
rect 24946 42702 24948 42754
rect 24892 42690 24948 42702
rect 25676 43650 25732 43662
rect 25676 43598 25678 43650
rect 25730 43598 25732 43650
rect 25004 42532 25060 42542
rect 24780 42530 25060 42532
rect 24780 42478 25006 42530
rect 25058 42478 25060 42530
rect 24780 42476 25060 42478
rect 25004 42466 25060 42476
rect 24220 42028 24388 42084
rect 25004 42308 25060 42318
rect 23772 41918 23774 41970
rect 23826 41918 23828 41970
rect 23772 41906 23828 41918
rect 23996 41972 24052 41982
rect 23996 41878 24052 41916
rect 23660 41794 23716 41804
rect 23548 41186 23604 41198
rect 23548 41134 23550 41186
rect 23602 41134 23604 41186
rect 23548 40964 23604 41134
rect 23548 40898 23604 40908
rect 24108 40404 24164 40414
rect 24108 40310 24164 40348
rect 23100 39678 23102 39730
rect 23154 39678 23156 39730
rect 23100 39666 23156 39678
rect 22876 39414 22932 39452
rect 23996 39618 24052 39630
rect 23996 39566 23998 39618
rect 24050 39566 24052 39618
rect 21868 39006 21870 39058
rect 21922 39006 21924 39058
rect 21868 38994 21924 39006
rect 22204 39060 22260 39070
rect 21644 37762 21700 37772
rect 21644 37268 21700 37278
rect 21644 37174 21700 37212
rect 21532 35186 21588 35196
rect 21756 36370 21812 36382
rect 21756 36318 21758 36370
rect 21810 36318 21812 36370
rect 20860 34690 20916 34702
rect 20860 34638 20862 34690
rect 20914 34638 20916 34690
rect 20860 34244 20916 34638
rect 20972 34692 21028 34702
rect 20972 34354 21028 34636
rect 20972 34302 20974 34354
rect 21026 34302 21028 34354
rect 20972 34290 21028 34302
rect 20860 34178 20916 34188
rect 20748 34066 20804 34076
rect 21084 34130 21140 34142
rect 21084 34078 21086 34130
rect 21138 34078 21140 34130
rect 20412 33394 20468 33404
rect 20076 33282 20132 33292
rect 20300 33122 20356 33134
rect 20300 33070 20302 33122
rect 20354 33070 20356 33122
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 18396 32564 18452 32574
rect 18396 32470 18452 32508
rect 17724 32162 17780 32172
rect 19516 32452 19572 32462
rect 17724 31780 17780 31790
rect 17724 31686 17780 31724
rect 18844 31556 18900 31566
rect 17836 31218 17892 31230
rect 17836 31166 17838 31218
rect 17890 31166 17892 31218
rect 17724 31108 17780 31118
rect 17612 31106 17780 31108
rect 17612 31054 17726 31106
rect 17778 31054 17780 31106
rect 17612 31052 17780 31054
rect 17724 31042 17780 31052
rect 17836 30884 17892 31166
rect 17836 30818 17892 30828
rect 18508 30882 18564 30894
rect 18508 30830 18510 30882
rect 18562 30830 18564 30882
rect 18508 30660 18564 30830
rect 18508 30594 18564 30604
rect 18620 30212 18676 30222
rect 18620 30118 18676 30156
rect 17500 29652 17556 29662
rect 17500 29558 17556 29596
rect 17948 29652 18004 29662
rect 17948 29558 18004 29596
rect 18844 29538 18900 31500
rect 19516 30994 19572 32396
rect 20076 32004 20132 32014
rect 20076 31666 20132 31948
rect 20076 31614 20078 31666
rect 20130 31614 20132 31666
rect 20076 31602 20132 31614
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19516 30942 19518 30994
rect 19570 30942 19572 30994
rect 19292 30884 19348 30894
rect 19516 30884 19572 30942
rect 20188 30994 20244 31006
rect 20188 30942 20190 30994
rect 20242 30942 20244 30994
rect 19292 30882 19684 30884
rect 19292 30830 19294 30882
rect 19346 30830 19684 30882
rect 19292 30828 19684 30830
rect 19068 30210 19124 30222
rect 19068 30158 19070 30210
rect 19122 30158 19124 30210
rect 19068 29652 19124 30158
rect 19292 29652 19348 30828
rect 19628 30322 19684 30828
rect 20188 30548 20244 30942
rect 20300 30996 20356 33070
rect 20860 33122 20916 33134
rect 20860 33070 20862 33122
rect 20914 33070 20916 33122
rect 20860 32676 20916 33070
rect 20860 32610 20916 32620
rect 21084 32452 21140 34078
rect 21644 34130 21700 34142
rect 21644 34078 21646 34130
rect 21698 34078 21700 34130
rect 21644 33796 21700 34078
rect 21756 33908 21812 36318
rect 22092 36372 22148 36382
rect 21756 33842 21812 33852
rect 21980 34132 22036 34142
rect 21644 33730 21700 33740
rect 21420 33460 21476 33470
rect 21420 33366 21476 33404
rect 21644 33234 21700 33246
rect 21644 33182 21646 33234
rect 21698 33182 21700 33234
rect 21084 32386 21140 32396
rect 21196 32788 21252 32798
rect 21196 31890 21252 32732
rect 21644 32452 21700 33182
rect 21644 32386 21700 32396
rect 21196 31838 21198 31890
rect 21250 31838 21252 31890
rect 21196 31826 21252 31838
rect 20972 31780 21028 31790
rect 20860 31668 20916 31678
rect 20860 31574 20916 31612
rect 20300 30930 20356 30940
rect 20188 30482 20244 30492
rect 19628 30270 19630 30322
rect 19682 30270 19684 30322
rect 19628 30258 19684 30270
rect 20300 30324 20356 30334
rect 20300 30210 20356 30268
rect 20300 30158 20302 30210
rect 20354 30158 20356 30210
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19124 29596 19348 29652
rect 19068 29586 19124 29596
rect 18844 29486 18846 29538
rect 18898 29486 18900 29538
rect 18844 29474 18900 29486
rect 17724 28980 17780 28990
rect 17724 28642 17780 28924
rect 17724 28590 17726 28642
rect 17778 28590 17780 28642
rect 17724 28578 17780 28590
rect 17948 28084 18004 28094
rect 17948 27990 18004 28028
rect 19292 28082 19348 29596
rect 20300 29652 20356 30158
rect 20748 30324 20804 30334
rect 20748 30210 20804 30268
rect 20748 30158 20750 30210
rect 20802 30158 20804 30210
rect 20748 30146 20804 30158
rect 20300 29558 20356 29596
rect 20860 29652 20916 29662
rect 20972 29652 21028 31724
rect 21980 31666 22036 34076
rect 22092 33460 22148 36316
rect 22204 35698 22260 39004
rect 22764 38724 22820 38734
rect 22652 38164 22708 38174
rect 22652 38070 22708 38108
rect 22652 36596 22708 36606
rect 22652 36502 22708 36540
rect 22204 35646 22206 35698
rect 22258 35646 22260 35698
rect 22204 35634 22260 35646
rect 22764 34914 22820 38668
rect 23996 38052 24052 39566
rect 24220 38834 24276 42028
rect 24332 41860 24388 41870
rect 24332 41766 24388 41804
rect 24780 41860 24836 41870
rect 24444 41300 24500 41310
rect 24444 41206 24500 41244
rect 24780 41298 24836 41804
rect 25004 41410 25060 42252
rect 25004 41358 25006 41410
rect 25058 41358 25060 41410
rect 25004 41346 25060 41358
rect 25452 41860 25508 41870
rect 24780 41246 24782 41298
rect 24834 41246 24836 41298
rect 24780 41234 24836 41246
rect 24668 40404 24724 40414
rect 24332 39620 24388 39630
rect 24332 39526 24388 39564
rect 24220 38782 24222 38834
rect 24274 38782 24276 38834
rect 24220 38770 24276 38782
rect 24668 38834 24724 40348
rect 25340 40292 25396 40302
rect 24780 40180 24836 40190
rect 24836 40124 24948 40180
rect 24780 40114 24836 40124
rect 24668 38782 24670 38834
rect 24722 38782 24724 38834
rect 23996 37958 24052 37996
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24556 37940 24612 37998
rect 24668 38052 24724 38782
rect 24668 37986 24724 37996
rect 24780 39956 24836 39966
rect 24556 37874 24612 37884
rect 23324 37826 23380 37838
rect 23324 37774 23326 37826
rect 23378 37774 23380 37826
rect 23212 36258 23268 36270
rect 23212 36206 23214 36258
rect 23266 36206 23268 36258
rect 23212 35924 23268 36206
rect 23324 36260 23380 37774
rect 24220 37490 24276 37502
rect 24220 37438 24222 37490
rect 24274 37438 24276 37490
rect 24220 37380 24276 37438
rect 24780 37490 24836 39900
rect 24780 37438 24782 37490
rect 24834 37438 24836 37490
rect 24780 37426 24836 37438
rect 24220 37314 24276 37324
rect 24220 36482 24276 36494
rect 24220 36430 24222 36482
rect 24274 36430 24276 36482
rect 23660 36260 23716 36270
rect 24220 36260 24276 36430
rect 24556 36484 24612 36494
rect 24556 36390 24612 36428
rect 23324 36258 24276 36260
rect 23324 36206 23662 36258
rect 23714 36206 24276 36258
rect 23324 36204 24276 36206
rect 23660 36194 23716 36204
rect 23268 35868 23492 35924
rect 23212 35858 23268 35868
rect 23436 35810 23492 35868
rect 23436 35758 23438 35810
rect 23490 35758 23492 35810
rect 23436 35746 23492 35758
rect 22876 35700 22932 35710
rect 22876 35606 22932 35644
rect 24220 35700 24276 36204
rect 24220 35028 24276 35644
rect 24444 35700 24500 35710
rect 24444 35586 24500 35644
rect 24444 35534 24446 35586
rect 24498 35534 24500 35586
rect 24444 35522 24500 35534
rect 24220 34962 24276 34972
rect 22764 34862 22766 34914
rect 22818 34862 22820 34914
rect 22764 33572 22820 34862
rect 24220 34354 24276 34366
rect 24220 34302 24222 34354
rect 24274 34302 24276 34354
rect 22428 33516 22708 33572
rect 22204 33460 22260 33470
rect 22428 33460 22484 33516
rect 22092 33458 22484 33460
rect 22092 33406 22206 33458
rect 22258 33406 22484 33458
rect 22092 33404 22484 33406
rect 22204 31892 22260 33404
rect 22540 33348 22596 33358
rect 22652 33348 22708 33516
rect 22764 33506 22820 33516
rect 23548 33572 23604 33582
rect 22764 33348 22820 33358
rect 22652 33346 22820 33348
rect 22652 33294 22766 33346
rect 22818 33294 22820 33346
rect 22652 33292 22820 33294
rect 22540 33254 22596 33292
rect 22764 33282 22820 33292
rect 23548 33234 23604 33516
rect 23548 33182 23550 33234
rect 23602 33182 23604 33234
rect 23548 32564 23604 33182
rect 24220 32676 24276 34302
rect 24780 34356 24836 34366
rect 24892 34356 24948 40124
rect 25228 37380 25284 37390
rect 25228 37286 25284 37324
rect 25340 36932 25396 40236
rect 25452 38722 25508 41804
rect 25676 41860 25732 43598
rect 25788 42642 25844 44044
rect 25788 42590 25790 42642
rect 25842 42590 25844 42642
rect 25788 42578 25844 42590
rect 25900 42308 25956 42318
rect 25676 41794 25732 41804
rect 25788 41858 25844 41870
rect 25788 41806 25790 41858
rect 25842 41806 25844 41858
rect 25788 41748 25844 41806
rect 25788 41300 25844 41692
rect 25676 41244 25844 41300
rect 25564 40516 25620 40526
rect 25564 40422 25620 40460
rect 25452 38670 25454 38722
rect 25506 38670 25508 38722
rect 25452 38658 25508 38670
rect 25676 40404 25732 41244
rect 25788 41076 25844 41086
rect 25900 41076 25956 42252
rect 26572 42084 26628 46510
rect 26684 45108 26740 45118
rect 26684 45014 26740 45052
rect 26572 42018 26628 42028
rect 26684 43426 26740 43438
rect 26684 43374 26686 43426
rect 26738 43374 26740 43426
rect 26124 41860 26180 41870
rect 26124 41858 26404 41860
rect 26124 41806 26126 41858
rect 26178 41806 26404 41858
rect 26124 41804 26404 41806
rect 26124 41794 26180 41804
rect 25788 41074 25956 41076
rect 25788 41022 25790 41074
rect 25842 41022 25956 41074
rect 25788 41020 25956 41022
rect 25788 41010 25844 41020
rect 26348 40740 26404 41804
rect 26460 41858 26516 41870
rect 26460 41806 26462 41858
rect 26514 41806 26516 41858
rect 26460 41748 26516 41806
rect 26460 41682 26516 41692
rect 26684 41300 26740 43374
rect 27132 41972 27188 41982
rect 27132 41878 27188 41916
rect 26684 41234 26740 41244
rect 26796 41858 26852 41870
rect 26796 41806 26798 41858
rect 26850 41806 26852 41858
rect 26348 40684 26740 40740
rect 25788 40628 25844 40638
rect 25788 40404 25844 40572
rect 25676 40402 25844 40404
rect 25676 40350 25790 40402
rect 25842 40350 25844 40402
rect 25676 40348 25844 40350
rect 25564 37380 25620 37390
rect 25676 37380 25732 40348
rect 25788 40338 25844 40348
rect 26460 40514 26516 40526
rect 26460 40462 26462 40514
rect 26514 40462 26516 40514
rect 25564 37378 25732 37380
rect 25564 37326 25566 37378
rect 25618 37326 25732 37378
rect 25564 37324 25732 37326
rect 25564 37314 25620 37324
rect 26124 37268 26180 37278
rect 25340 36866 25396 36876
rect 26012 37266 26180 37268
rect 26012 37214 26126 37266
rect 26178 37214 26180 37266
rect 26012 37212 26180 37214
rect 24780 34354 24948 34356
rect 24780 34302 24782 34354
rect 24834 34302 24948 34354
rect 24780 34300 24948 34302
rect 25340 35700 25396 35710
rect 24780 34290 24836 34300
rect 25340 34130 25396 35644
rect 26012 35700 26068 37212
rect 26124 37202 26180 37212
rect 26460 36484 26516 40462
rect 26684 39506 26740 40684
rect 26796 39620 26852 41806
rect 27244 41636 27300 47292
rect 27356 45220 27412 45230
rect 27356 41748 27412 45164
rect 27468 44098 27524 44110
rect 27468 44046 27470 44098
rect 27522 44046 27524 44098
rect 27468 41970 27524 44046
rect 27580 42756 27636 50372
rect 27804 43652 27860 51436
rect 27916 51426 27972 51436
rect 27916 49700 27972 49710
rect 27916 49606 27972 49644
rect 27916 49252 27972 49262
rect 28028 49252 28084 51996
rect 28140 51986 28196 51996
rect 28476 51490 28532 51502
rect 28476 51438 28478 51490
rect 28530 51438 28532 51490
rect 27916 49250 28084 49252
rect 27916 49198 27918 49250
rect 27970 49198 28084 49250
rect 27916 49196 28084 49198
rect 28140 49700 28196 49710
rect 27916 49186 27972 49196
rect 28140 49138 28196 49644
rect 28252 49700 28308 49710
rect 28252 49698 28420 49700
rect 28252 49646 28254 49698
rect 28306 49646 28420 49698
rect 28252 49644 28420 49646
rect 28252 49634 28308 49644
rect 28140 49086 28142 49138
rect 28194 49086 28196 49138
rect 28140 49074 28196 49086
rect 28028 48916 28084 48926
rect 27916 47236 27972 47246
rect 27916 45778 27972 47180
rect 27916 45726 27918 45778
rect 27970 45726 27972 45778
rect 27916 45714 27972 45726
rect 28028 44546 28084 48860
rect 28252 48804 28308 48814
rect 28252 48710 28308 48748
rect 28140 47234 28196 47246
rect 28140 47182 28142 47234
rect 28194 47182 28196 47234
rect 28140 46900 28196 47182
rect 28140 46834 28196 46844
rect 28140 46676 28196 46686
rect 28140 45444 28196 46620
rect 28364 46340 28420 49644
rect 28476 48804 28532 51438
rect 28476 48738 28532 48748
rect 28588 46674 28644 53788
rect 30380 53844 30436 53854
rect 33628 53844 33684 53854
rect 38556 53844 38612 53854
rect 41356 53844 41412 53854
rect 30380 53750 30436 53788
rect 33516 53842 33684 53844
rect 33516 53790 33630 53842
rect 33682 53790 33684 53842
rect 33516 53788 33684 53790
rect 31388 53618 31444 53630
rect 31388 53566 31390 53618
rect 31442 53566 31444 53618
rect 31052 52834 31108 52846
rect 31052 52782 31054 52834
rect 31106 52782 31108 52834
rect 30716 52050 30772 52062
rect 30716 51998 30718 52050
rect 30770 51998 30772 52050
rect 29036 51492 29092 51502
rect 29036 51398 29092 51436
rect 30156 51268 30212 51278
rect 30044 51266 30212 51268
rect 30044 51214 30158 51266
rect 30210 51214 30212 51266
rect 30044 51212 30212 51214
rect 29372 49922 29428 49934
rect 29372 49870 29374 49922
rect 29426 49870 29428 49922
rect 28700 48916 28756 48926
rect 28700 47682 28756 48860
rect 29260 48914 29316 48926
rect 29260 48862 29262 48914
rect 29314 48862 29316 48914
rect 28700 47630 28702 47682
rect 28754 47630 28756 47682
rect 28700 47618 28756 47630
rect 28812 48804 28868 48814
rect 28588 46622 28590 46674
rect 28642 46622 28644 46674
rect 28588 46610 28644 46622
rect 28364 46274 28420 46284
rect 28700 46116 28756 46126
rect 28812 46116 28868 48748
rect 29260 48466 29316 48862
rect 29260 48414 29262 48466
rect 29314 48414 29316 48466
rect 29260 48402 29316 48414
rect 29036 47458 29092 47470
rect 29036 47406 29038 47458
rect 29090 47406 29092 47458
rect 29036 46676 29092 47406
rect 29036 46610 29092 46620
rect 28700 46114 28868 46116
rect 28700 46062 28702 46114
rect 28754 46062 28868 46114
rect 28700 46060 28868 46062
rect 29036 46116 29092 46126
rect 28700 46050 28756 46060
rect 29036 46022 29092 46060
rect 28140 45388 28644 45444
rect 28028 44494 28030 44546
rect 28082 44494 28084 44546
rect 28028 44482 28084 44494
rect 28588 45218 28644 45388
rect 28588 45166 28590 45218
rect 28642 45166 28644 45218
rect 28252 44212 28308 44222
rect 28028 44210 28308 44212
rect 28028 44158 28254 44210
rect 28306 44158 28308 44210
rect 28028 44156 28308 44158
rect 27916 43652 27972 43662
rect 27804 43650 27972 43652
rect 27804 43598 27918 43650
rect 27970 43598 27972 43650
rect 27804 43596 27972 43598
rect 27916 43586 27972 43596
rect 27692 43428 27748 43438
rect 28028 43428 28084 44156
rect 28252 44146 28308 44156
rect 28364 44100 28420 44110
rect 28364 44006 28420 44044
rect 27692 43426 28196 43428
rect 27692 43374 27694 43426
rect 27746 43374 28196 43426
rect 27692 43372 28196 43374
rect 27692 43362 27748 43372
rect 28028 42756 28084 42766
rect 27580 42754 28084 42756
rect 27580 42702 28030 42754
rect 28082 42702 28084 42754
rect 27580 42700 28084 42702
rect 28028 42690 28084 42700
rect 27468 41918 27470 41970
rect 27522 41918 27524 41970
rect 27468 41906 27524 41918
rect 27916 42532 27972 42542
rect 27916 41970 27972 42476
rect 27916 41918 27918 41970
rect 27970 41918 27972 41970
rect 27916 41906 27972 41918
rect 28140 41972 28196 43372
rect 28028 41748 28084 41758
rect 27356 41692 27636 41748
rect 27244 41580 27524 41636
rect 27132 40964 27188 40974
rect 26796 39564 26964 39620
rect 26684 39454 26686 39506
rect 26738 39454 26740 39506
rect 26684 39442 26740 39454
rect 26908 37938 26964 39564
rect 26908 37886 26910 37938
rect 26962 37886 26964 37938
rect 26908 37874 26964 37886
rect 26460 36418 26516 36428
rect 26012 35606 26068 35644
rect 27020 36258 27076 36270
rect 27020 36206 27022 36258
rect 27074 36206 27076 36258
rect 26348 35028 26404 35038
rect 26348 34934 26404 34972
rect 27020 35026 27076 36206
rect 27020 34974 27022 35026
rect 27074 34974 27076 35026
rect 27020 34962 27076 34974
rect 25340 34078 25342 34130
rect 25394 34078 25396 34130
rect 25340 34066 25396 34078
rect 27132 34242 27188 40908
rect 27468 39842 27524 41580
rect 27468 39790 27470 39842
rect 27522 39790 27524 39842
rect 27468 39778 27524 39790
rect 27580 36708 27636 41692
rect 27916 41636 27972 41646
rect 27692 40290 27748 40302
rect 27692 40238 27694 40290
rect 27746 40238 27748 40290
rect 27692 38668 27748 40238
rect 27916 40180 27972 41580
rect 28028 41186 28084 41692
rect 28028 41134 28030 41186
rect 28082 41134 28084 41186
rect 28028 41122 28084 41134
rect 28140 40626 28196 41916
rect 28252 42868 28308 42878
rect 28252 41970 28308 42812
rect 28588 42754 28644 45166
rect 29148 45108 29204 45118
rect 28700 43652 28756 43662
rect 28700 43558 28756 43596
rect 28588 42702 28590 42754
rect 28642 42702 28644 42754
rect 28476 42532 28532 42542
rect 28588 42532 28644 42702
rect 28532 42476 28644 42532
rect 28476 42466 28532 42476
rect 28252 41918 28254 41970
rect 28306 41918 28308 41970
rect 28252 41906 28308 41918
rect 28588 41186 28644 41198
rect 28588 41134 28590 41186
rect 28642 41134 28644 41186
rect 28140 40574 28142 40626
rect 28194 40574 28196 40626
rect 28140 40562 28196 40574
rect 28476 40740 28532 40750
rect 27916 40124 28084 40180
rect 27916 39732 27972 39742
rect 27916 39638 27972 39676
rect 28028 39058 28084 40124
rect 28476 39394 28532 40684
rect 28588 40404 28644 41134
rect 28588 40338 28644 40348
rect 28700 40516 28756 40526
rect 28700 40068 28756 40460
rect 28588 40012 28756 40068
rect 28924 40404 28980 40414
rect 28588 39730 28644 40012
rect 28588 39678 28590 39730
rect 28642 39678 28644 39730
rect 28588 39666 28644 39678
rect 28476 39342 28478 39394
rect 28530 39342 28532 39394
rect 28476 39330 28532 39342
rect 28028 39006 28030 39058
rect 28082 39006 28084 39058
rect 28028 38994 28084 39006
rect 28812 38948 28868 38958
rect 28812 38854 28868 38892
rect 27804 38836 27860 38846
rect 27804 38834 27972 38836
rect 27804 38782 27806 38834
rect 27858 38782 27972 38834
rect 27804 38780 27972 38782
rect 27804 38770 27860 38780
rect 27916 38724 27972 38780
rect 28028 38724 28084 38734
rect 27916 38668 28028 38724
rect 27692 38612 27860 38668
rect 27692 38388 27748 38398
rect 27692 38274 27748 38332
rect 27692 38222 27694 38274
rect 27746 38222 27748 38274
rect 27692 38210 27748 38222
rect 27804 37268 27860 38612
rect 27804 37202 27860 37212
rect 28028 38162 28084 38668
rect 28028 38110 28030 38162
rect 28082 38110 28084 38162
rect 28028 37154 28084 38110
rect 28028 37102 28030 37154
rect 28082 37102 28084 37154
rect 28028 37090 28084 37102
rect 28364 38276 28420 38286
rect 27692 36708 27748 36718
rect 27580 36706 27748 36708
rect 27580 36654 27694 36706
rect 27746 36654 27748 36706
rect 27580 36652 27748 36654
rect 27692 36642 27748 36652
rect 28028 36258 28084 36270
rect 28028 36206 28030 36258
rect 28082 36206 28084 36258
rect 27804 35586 27860 35598
rect 27804 35534 27806 35586
rect 27858 35534 27860 35586
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 25788 33348 25844 33358
rect 24556 33012 24612 33022
rect 24332 32676 24388 32686
rect 24220 32674 24388 32676
rect 24220 32622 24334 32674
rect 24386 32622 24388 32674
rect 24220 32620 24388 32622
rect 24332 32610 24388 32620
rect 22204 31826 22260 31836
rect 22316 32452 22372 32462
rect 21980 31614 21982 31666
rect 22034 31614 22036 31666
rect 21980 31602 22036 31614
rect 21308 30996 21364 31006
rect 21364 30940 21476 30996
rect 21308 30930 21364 30940
rect 20860 29650 21028 29652
rect 20860 29598 20862 29650
rect 20914 29598 21028 29650
rect 20860 29596 21028 29598
rect 21308 30324 21364 30334
rect 20860 29586 20916 29596
rect 21308 29426 21364 30268
rect 21420 30322 21476 30940
rect 21420 30270 21422 30322
rect 21474 30270 21476 30322
rect 21420 30258 21476 30270
rect 21644 30212 21700 30222
rect 21644 30118 21700 30156
rect 22316 30212 22372 32396
rect 22988 32450 23044 32462
rect 22988 32398 22990 32450
rect 23042 32398 23044 32450
rect 22988 32004 23044 32398
rect 23324 32452 23380 32462
rect 23324 32358 23380 32396
rect 22988 31938 23044 31948
rect 22540 31218 22596 31230
rect 22540 31166 22542 31218
rect 22594 31166 22596 31218
rect 22540 30322 22596 31166
rect 23548 30884 23604 32508
rect 23772 32562 23828 32574
rect 23772 32510 23774 32562
rect 23826 32510 23828 32562
rect 23772 32452 23828 32510
rect 23772 32386 23828 32396
rect 23884 32450 23940 32462
rect 23884 32398 23886 32450
rect 23938 32398 23940 32450
rect 23548 30790 23604 30828
rect 23212 30770 23268 30782
rect 23212 30718 23214 30770
rect 23266 30718 23268 30770
rect 23212 30436 23268 30718
rect 23212 30370 23268 30380
rect 22540 30270 22542 30322
rect 22594 30270 22596 30322
rect 22540 30258 22596 30270
rect 22316 30118 22372 30156
rect 23548 29986 23604 29998
rect 23548 29934 23550 29986
rect 23602 29934 23604 29986
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 21308 29362 21364 29374
rect 21644 29428 21700 29438
rect 21644 29334 21700 29372
rect 19852 29316 19908 29326
rect 19852 29222 19908 29260
rect 22540 29204 22596 29214
rect 21532 28642 21588 28654
rect 21532 28590 21534 28642
rect 21586 28590 21588 28642
rect 20300 28418 20356 28430
rect 20860 28420 20916 28430
rect 21308 28420 21364 28430
rect 20300 28366 20302 28418
rect 20354 28366 20356 28418
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19292 28030 19294 28082
rect 19346 28030 19348 28082
rect 19292 28018 19348 28030
rect 18172 27858 18228 27870
rect 18172 27806 18174 27858
rect 18226 27806 18228 27858
rect 17612 27748 17668 27758
rect 17612 27654 17668 27692
rect 18172 27748 18228 27806
rect 18172 27682 18228 27692
rect 19740 27748 19796 27758
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 24724 16884 26126
rect 17164 26852 17332 26908
rect 17388 27074 17444 27086
rect 17388 27022 17390 27074
rect 17442 27022 17444 27074
rect 17164 25844 17220 26852
rect 17276 26068 17332 26106
rect 17276 26002 17332 26012
rect 17276 25844 17332 25854
rect 17164 25788 17276 25844
rect 16828 24668 17108 24724
rect 16828 24500 16884 24510
rect 16828 23154 16884 24444
rect 16828 23102 16830 23154
rect 16882 23102 16884 23154
rect 16828 23090 16884 23102
rect 16940 24498 16996 24510
rect 16940 24446 16942 24498
rect 16994 24446 16996 24498
rect 16940 21588 16996 24446
rect 17052 23716 17108 24668
rect 17276 23938 17332 25788
rect 17388 25284 17444 27022
rect 17388 25218 17444 25228
rect 17724 27074 17780 27086
rect 17724 27022 17726 27074
rect 17778 27022 17780 27074
rect 17612 24724 17668 24734
rect 17612 24630 17668 24668
rect 17276 23886 17278 23938
rect 17330 23886 17332 23938
rect 17276 23874 17332 23886
rect 17052 23660 17444 23716
rect 17276 22930 17332 22942
rect 17276 22878 17278 22930
rect 17330 22878 17332 22930
rect 17164 22372 17220 22382
rect 17164 22278 17220 22316
rect 17052 22148 17108 22158
rect 17052 22054 17108 22092
rect 17276 21812 17332 22878
rect 17276 21746 17332 21756
rect 16940 21532 17332 21588
rect 16940 21362 16996 21374
rect 16940 21310 16942 21362
rect 16994 21310 16996 21362
rect 16716 21084 16884 21140
rect 16716 20916 16772 20926
rect 16716 20188 16772 20860
rect 16828 20580 16884 21084
rect 16828 20514 16884 20524
rect 16716 20132 16884 20188
rect 16828 20130 16884 20132
rect 16828 20078 16830 20130
rect 16882 20078 16884 20130
rect 16828 20020 16884 20078
rect 16828 19954 16884 19964
rect 16828 19348 16884 19358
rect 16828 19254 16884 19292
rect 16940 19124 16996 21310
rect 16604 17726 16606 17778
rect 16658 17726 16660 17778
rect 16604 17714 16660 17726
rect 16716 19068 16996 19124
rect 16716 16994 16772 19068
rect 17276 17556 17332 21532
rect 17388 21586 17444 23660
rect 17388 21534 17390 21586
rect 17442 21534 17444 21586
rect 17388 19908 17444 21534
rect 17500 22372 17556 22382
rect 17500 20132 17556 22316
rect 17500 20038 17556 20076
rect 17612 22036 17668 22046
rect 17388 19012 17444 19852
rect 17500 19012 17556 19022
rect 17388 18956 17500 19012
rect 17500 18946 17556 18956
rect 17500 17556 17556 17566
rect 17276 17554 17556 17556
rect 17276 17502 17502 17554
rect 17554 17502 17556 17554
rect 17276 17500 17556 17502
rect 17500 17490 17556 17500
rect 16716 16942 16718 16994
rect 16770 16942 16772 16994
rect 16716 16930 16772 16942
rect 16156 15934 16158 15986
rect 16210 15934 16212 15986
rect 16156 15922 16212 15934
rect 17612 15148 17668 21980
rect 17724 19348 17780 27022
rect 19740 27076 19796 27692
rect 19740 27010 19796 27020
rect 19964 27634 20020 27646
rect 19964 27582 19966 27634
rect 20018 27582 20020 27634
rect 19964 26852 20020 27582
rect 20300 27300 20356 28366
rect 20300 27234 20356 27244
rect 20636 28418 20916 28420
rect 20636 28366 20862 28418
rect 20914 28366 20916 28418
rect 20636 28364 20916 28366
rect 20076 26964 20132 26974
rect 20636 26908 20692 28364
rect 20860 28354 20916 28364
rect 20972 28418 21364 28420
rect 20972 28366 21310 28418
rect 21362 28366 21364 28418
rect 20972 28364 21364 28366
rect 20972 28196 21028 28364
rect 21308 28354 21364 28364
rect 20748 28140 21028 28196
rect 20748 28082 20804 28140
rect 20748 28030 20750 28082
rect 20802 28030 20804 28082
rect 20748 28018 20804 28030
rect 20076 26870 20132 26908
rect 19964 26786 20020 26796
rect 20524 26852 20692 26908
rect 20748 27748 20804 27758
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18284 26516 18340 26526
rect 18060 26402 18116 26414
rect 18060 26350 18062 26402
rect 18114 26350 18116 26402
rect 18060 25732 18116 26350
rect 18060 25666 18116 25676
rect 17948 25060 18004 25070
rect 17948 24724 18004 25004
rect 17948 24630 18004 24668
rect 18060 23266 18116 23278
rect 18060 23214 18062 23266
rect 18114 23214 18116 23266
rect 17836 22370 17892 22382
rect 17836 22318 17838 22370
rect 17890 22318 17892 22370
rect 17836 20356 17892 22318
rect 17836 20290 17892 20300
rect 18060 20244 18116 23214
rect 18060 20178 18116 20188
rect 18172 20580 18228 20590
rect 18172 20130 18228 20524
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20066 18228 20078
rect 17836 20020 17892 20030
rect 17836 19926 17892 19964
rect 17724 19282 17780 19292
rect 18284 18562 18340 26460
rect 19516 26292 19572 26302
rect 19404 25732 19460 25742
rect 19404 25638 19460 25676
rect 19180 25396 19236 25406
rect 18956 25394 19236 25396
rect 18956 25342 19182 25394
rect 19234 25342 19236 25394
rect 18956 25340 19236 25342
rect 18396 25282 18452 25294
rect 18396 25230 18398 25282
rect 18450 25230 18452 25282
rect 18396 24610 18452 25230
rect 18396 24558 18398 24610
rect 18450 24558 18452 24610
rect 18396 24546 18452 24558
rect 18844 24500 18900 24510
rect 18732 20580 18788 20590
rect 18732 20486 18788 20524
rect 18620 20356 18676 20366
rect 18844 20356 18900 24444
rect 18508 20244 18564 20254
rect 18508 20130 18564 20188
rect 18508 20078 18510 20130
rect 18562 20078 18564 20130
rect 18508 20066 18564 20078
rect 18508 19572 18564 19582
rect 18508 18788 18564 19516
rect 18284 18510 18286 18562
rect 18338 18510 18340 18562
rect 18284 18498 18340 18510
rect 18396 18732 18564 18788
rect 18396 16994 18452 18732
rect 18396 16942 18398 16994
rect 18450 16942 18452 16994
rect 18396 16930 18452 16942
rect 18620 16212 18676 20300
rect 18732 20300 18900 20356
rect 18732 19122 18788 20300
rect 18844 20020 18900 20030
rect 18844 19926 18900 19964
rect 18732 19070 18734 19122
rect 18786 19070 18788 19122
rect 18732 19058 18788 19070
rect 18732 17556 18788 17566
rect 18956 17556 19012 25340
rect 19180 25330 19236 25340
rect 19292 25396 19348 25406
rect 19180 25172 19236 25182
rect 19180 24946 19236 25116
rect 19180 24894 19182 24946
rect 19234 24894 19236 24946
rect 19180 24836 19236 24894
rect 19180 24770 19236 24780
rect 19068 24052 19124 24062
rect 19068 23958 19124 23996
rect 19292 23938 19348 25340
rect 19292 23886 19294 23938
rect 19346 23886 19348 23938
rect 19068 21812 19124 21822
rect 19124 21756 19236 21812
rect 19068 21746 19124 21756
rect 19068 20132 19124 20142
rect 19068 20018 19124 20076
rect 19068 19966 19070 20018
rect 19122 19966 19124 20018
rect 19068 19954 19124 19966
rect 18732 17554 19012 17556
rect 18732 17502 18734 17554
rect 18786 17502 19012 17554
rect 18732 17500 19012 17502
rect 19068 18564 19124 18574
rect 18732 17490 18788 17500
rect 18732 16212 18788 16222
rect 18620 16210 18788 16212
rect 18620 16158 18734 16210
rect 18786 16158 18788 16210
rect 18620 16156 18788 16158
rect 18732 16146 18788 16156
rect 17612 15092 17892 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 17836 14644 17892 15092
rect 18172 14644 18228 14654
rect 17836 14642 18228 14644
rect 17836 14590 18174 14642
rect 18226 14590 18228 14642
rect 17836 14588 18228 14590
rect 18172 14578 18228 14588
rect 19068 14420 19124 18508
rect 19180 16436 19236 21756
rect 19292 21362 19348 23886
rect 19516 23380 19572 26236
rect 20412 26290 20468 26302
rect 20412 26238 20414 26290
rect 20466 26238 20468 26290
rect 19628 25506 19684 25518
rect 19628 25454 19630 25506
rect 19682 25454 19684 25506
rect 19628 25172 19684 25454
rect 20188 25508 20244 25518
rect 19628 25106 19684 25116
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 25452
rect 20076 24892 20244 24948
rect 20300 25284 20356 25294
rect 19628 24836 19684 24846
rect 19628 24742 19684 24780
rect 19852 24500 19908 24510
rect 19852 24406 19908 24444
rect 19964 24052 20020 24062
rect 20076 24052 20132 24892
rect 19964 24050 20132 24052
rect 19964 23998 19966 24050
rect 20018 23998 20132 24050
rect 19964 23996 20132 23998
rect 20300 24050 20356 25228
rect 20300 23998 20302 24050
rect 20354 23998 20356 24050
rect 19964 23986 20020 23996
rect 20300 23940 20356 23998
rect 20300 23874 20356 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19516 23324 19684 23380
rect 19516 23156 19572 23166
rect 19292 21310 19294 21362
rect 19346 21310 19348 21362
rect 19292 20916 19348 21310
rect 19292 20020 19348 20860
rect 19292 19954 19348 19964
rect 19404 23100 19516 23156
rect 19404 16770 19460 23100
rect 19516 23090 19572 23100
rect 19516 20578 19572 20590
rect 19516 20526 19518 20578
rect 19570 20526 19572 20578
rect 19516 19572 19572 20526
rect 19628 20244 19684 23324
rect 20300 23156 20356 23166
rect 20300 23062 20356 23100
rect 20188 22146 20244 22158
rect 20188 22094 20190 22146
rect 20242 22094 20244 22146
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22094
rect 20076 21756 20244 21812
rect 19740 20916 19796 20926
rect 19740 20822 19796 20860
rect 20076 20914 20132 21756
rect 20412 21588 20468 26238
rect 20076 20862 20078 20914
rect 20130 20862 20132 20914
rect 20076 20850 20132 20862
rect 20188 21532 20468 21588
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19628 20188 19796 20244
rect 19516 19506 19572 19516
rect 19628 20018 19684 20030
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 19516 19236 19572 19246
rect 19516 18338 19572 19180
rect 19516 18286 19518 18338
rect 19570 18286 19572 18338
rect 19516 18274 19572 18286
rect 19404 16718 19406 16770
rect 19458 16718 19460 16770
rect 19404 16706 19460 16718
rect 19628 16660 19684 19966
rect 19740 19346 19796 20188
rect 19740 19294 19742 19346
rect 19794 19294 19796 19346
rect 19740 19282 19796 19294
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18452 20244 21532
rect 20412 21364 20468 21374
rect 20300 21362 20468 21364
rect 20300 21310 20414 21362
rect 20466 21310 20468 21362
rect 20300 21308 20468 21310
rect 20300 19236 20356 21308
rect 20412 21298 20468 21308
rect 20412 20916 20468 20926
rect 20412 20822 20468 20860
rect 20300 19180 20468 19236
rect 20300 19012 20356 19022
rect 20300 18918 20356 18956
rect 19740 18396 20244 18452
rect 19740 17778 19796 18396
rect 19740 17726 19742 17778
rect 19794 17726 19796 17778
rect 19740 17714 19796 17726
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20412 16772 20468 19180
rect 20524 16996 20580 26852
rect 20636 25508 20692 25546
rect 20748 25508 20804 27692
rect 21308 27300 21364 27310
rect 21308 27206 21364 27244
rect 21532 27076 21588 28590
rect 22316 28642 22372 28654
rect 22316 28590 22318 28642
rect 22370 28590 22372 28642
rect 22316 27860 22372 28590
rect 22316 27794 22372 27804
rect 21532 26908 21588 27020
rect 22428 27076 22484 27086
rect 22428 26982 22484 27020
rect 20860 26850 20916 26862
rect 20860 26798 20862 26850
rect 20914 26798 20916 26850
rect 20860 26516 20916 26798
rect 20860 26450 20916 26460
rect 21308 26852 21588 26908
rect 22204 26852 22260 26862
rect 20692 25452 20804 25508
rect 20860 26292 20916 26302
rect 21084 26292 21140 26302
rect 20860 26290 21140 26292
rect 20860 26238 20862 26290
rect 20914 26238 21086 26290
rect 21138 26238 21140 26290
rect 20860 26236 21140 26238
rect 20636 25442 20692 25452
rect 20636 25282 20692 25294
rect 20636 25230 20638 25282
rect 20690 25230 20692 25282
rect 20636 24946 20692 25230
rect 20748 25284 20804 25294
rect 20860 25284 20916 26236
rect 21084 26226 21140 26236
rect 20804 25228 20916 25284
rect 20748 25218 20804 25228
rect 20636 24894 20638 24946
rect 20690 24894 20692 24946
rect 20636 24882 20692 24894
rect 20748 24948 20804 24958
rect 20748 24050 20804 24892
rect 21308 24948 21364 26852
rect 21868 26850 22260 26852
rect 21868 26798 22206 26850
rect 22258 26798 22260 26850
rect 21868 26796 22260 26798
rect 21532 26740 21588 26750
rect 21532 26068 21588 26684
rect 21756 26404 21812 26414
rect 21644 26292 21700 26302
rect 21644 26198 21700 26236
rect 21532 26012 21700 26068
rect 21420 25396 21476 25406
rect 21420 25302 21476 25340
rect 21308 24882 21364 24892
rect 20748 23998 20750 24050
rect 20802 23998 20804 24050
rect 20748 23986 20804 23998
rect 21196 23940 21252 23950
rect 21196 23846 21252 23884
rect 20748 23154 20804 23166
rect 20748 23102 20750 23154
rect 20802 23102 20804 23154
rect 20748 22372 20804 23102
rect 21084 22932 21140 22942
rect 21084 22930 21588 22932
rect 21084 22878 21086 22930
rect 21138 22878 21588 22930
rect 21084 22876 21588 22878
rect 21084 22866 21140 22876
rect 20748 22306 20804 22316
rect 20860 22148 20916 22158
rect 20860 22146 21364 22148
rect 20860 22094 20862 22146
rect 20914 22094 21364 22146
rect 20860 22092 21364 22094
rect 20860 22082 20916 22092
rect 20972 21812 21028 21822
rect 20636 21810 21028 21812
rect 20636 21758 20974 21810
rect 21026 21758 21028 21810
rect 20636 21756 21028 21758
rect 20636 20914 20692 21756
rect 20972 21746 21028 21756
rect 20636 20862 20638 20914
rect 20690 20862 20692 20914
rect 20636 20850 20692 20862
rect 20636 20132 20692 20142
rect 20636 19348 20692 20076
rect 20636 19254 20692 19292
rect 20972 16996 21028 17006
rect 20524 16994 21028 16996
rect 20524 16942 20974 16994
rect 21026 16942 21028 16994
rect 20524 16940 21028 16942
rect 20972 16930 21028 16940
rect 20412 16706 20468 16716
rect 19740 16660 19796 16670
rect 19628 16604 19740 16660
rect 19740 16594 19796 16604
rect 20300 16660 20356 16670
rect 19180 16380 19796 16436
rect 19740 15986 19796 16380
rect 19740 15934 19742 15986
rect 19794 15934 19796 15986
rect 19740 15922 19796 15934
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15202 20356 16604
rect 21308 15426 21364 22092
rect 21420 19348 21476 19358
rect 21420 19254 21476 19292
rect 21532 18452 21588 22876
rect 21644 20690 21700 26012
rect 21756 25618 21812 26348
rect 21756 25566 21758 25618
rect 21810 25566 21812 25618
rect 21756 25554 21812 25566
rect 21756 23938 21812 23950
rect 21756 23886 21758 23938
rect 21810 23886 21812 23938
rect 21756 23156 21812 23886
rect 21868 23378 21924 26796
rect 22204 26786 22260 26796
rect 22540 25394 22596 29148
rect 23548 29092 23604 29934
rect 23884 29652 23940 32398
rect 23996 31780 24052 31790
rect 23996 31218 24052 31724
rect 24220 31778 24276 31790
rect 24220 31726 24222 31778
rect 24274 31726 24276 31778
rect 24220 31668 24276 31726
rect 24220 31602 24276 31612
rect 23996 31166 23998 31218
rect 24050 31166 24052 31218
rect 23996 30324 24052 31166
rect 23996 30258 24052 30268
rect 24332 30436 24388 30446
rect 24332 30098 24388 30380
rect 24332 30046 24334 30098
rect 24386 30046 24388 30098
rect 24332 30034 24388 30046
rect 23996 29652 24052 29662
rect 23884 29650 24052 29652
rect 23884 29598 23998 29650
rect 24050 29598 24052 29650
rect 23884 29596 24052 29598
rect 23996 29586 24052 29596
rect 24556 29316 24612 32956
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 24668 31780 24724 31790
rect 24668 31686 24724 31724
rect 25788 31666 25844 33292
rect 25788 31614 25790 31666
rect 25842 31614 25844 31666
rect 25788 31602 25844 31614
rect 25900 32564 25956 32574
rect 25004 31556 25060 31566
rect 25004 31462 25060 31500
rect 25452 31220 25508 31230
rect 25452 31126 25508 31164
rect 25900 30660 25956 32508
rect 27132 32564 27188 34190
rect 27132 32498 27188 32508
rect 27244 34804 27300 34814
rect 27580 34804 27636 34814
rect 27244 34802 27636 34804
rect 27244 34750 27246 34802
rect 27298 34750 27582 34802
rect 27634 34750 27636 34802
rect 27244 34748 27636 34750
rect 27244 32674 27300 34748
rect 27580 34738 27636 34748
rect 27692 34690 27748 34702
rect 27692 34638 27694 34690
rect 27746 34638 27748 34690
rect 27692 33348 27748 34638
rect 27692 33282 27748 33292
rect 27244 32622 27246 32674
rect 27298 32622 27300 32674
rect 26684 32452 26740 32462
rect 26684 31948 26740 32396
rect 27244 31948 27300 32622
rect 26684 31892 27524 31948
rect 26572 31668 26628 31678
rect 26012 30884 26068 30894
rect 26068 30828 26180 30884
rect 26012 30790 26068 30828
rect 25956 30604 26068 30660
rect 25900 30594 25956 30604
rect 24556 29250 24612 29260
rect 25116 29988 25172 29998
rect 24780 29204 24836 29214
rect 24780 29202 25060 29204
rect 24780 29150 24782 29202
rect 24834 29150 25060 29202
rect 24780 29148 25060 29150
rect 24780 29138 24836 29148
rect 24444 29092 24500 29102
rect 23548 29026 23604 29036
rect 24332 29036 24444 29092
rect 22540 25342 22542 25394
rect 22594 25342 22596 25394
rect 22540 25330 22596 25342
rect 22652 28642 22708 28654
rect 22652 28590 22654 28642
rect 22706 28590 22708 28642
rect 21868 23326 21870 23378
rect 21922 23326 21924 23378
rect 21868 23314 21924 23326
rect 21756 23100 22260 23156
rect 22092 22596 22148 22606
rect 21644 20638 21646 20690
rect 21698 20638 21700 20690
rect 21644 20626 21700 20638
rect 21756 20916 21812 20926
rect 21756 20188 21812 20860
rect 21756 20132 21924 20188
rect 21868 19346 21924 20132
rect 21868 19294 21870 19346
rect 21922 19294 21924 19346
rect 21868 19282 21924 19294
rect 21980 20130 22036 20142
rect 21980 20078 21982 20130
rect 22034 20078 22036 20130
rect 21980 19010 22036 20078
rect 22092 19236 22148 22540
rect 22092 19170 22148 19180
rect 21980 18958 21982 19010
rect 22034 18958 22036 19010
rect 21980 18946 22036 18958
rect 21532 18386 21588 18396
rect 21868 18340 21924 18350
rect 21868 18246 21924 18284
rect 22204 16212 22260 23100
rect 22652 20914 22708 28590
rect 24220 28196 24276 28206
rect 23772 27972 23828 27982
rect 22988 27858 23044 27870
rect 22988 27806 22990 27858
rect 23042 27806 23044 27858
rect 22876 24724 22932 24734
rect 22764 24722 22932 24724
rect 22764 24670 22878 24722
rect 22930 24670 22932 24722
rect 22764 24668 22932 24670
rect 22764 22596 22820 24668
rect 22876 24658 22932 24668
rect 22988 22820 23044 27806
rect 23212 27860 23268 27870
rect 22764 22530 22820 22540
rect 22876 22764 23044 22820
rect 23100 27636 23156 27646
rect 22764 22372 22820 22382
rect 22764 22278 22820 22316
rect 22652 20862 22654 20914
rect 22706 20862 22708 20914
rect 22652 20850 22708 20862
rect 22876 20692 22932 22764
rect 23100 22708 23156 27580
rect 23212 27074 23268 27804
rect 23660 27860 23716 27870
rect 23660 27766 23716 27804
rect 23212 27022 23214 27074
rect 23266 27022 23268 27074
rect 23212 27010 23268 27022
rect 23660 27076 23716 27086
rect 23660 26982 23716 27020
rect 23772 26908 23828 27916
rect 24220 27970 24276 28140
rect 24220 27918 24222 27970
rect 24274 27918 24276 27970
rect 24108 27860 24164 27870
rect 23548 26852 23828 26908
rect 23884 27746 23940 27758
rect 23884 27694 23886 27746
rect 23938 27694 23940 27746
rect 23884 26964 23940 27694
rect 23884 26898 23940 26908
rect 23548 25618 23604 26852
rect 23996 26404 24052 26414
rect 23996 26310 24052 26348
rect 23548 25566 23550 25618
rect 23602 25566 23604 25618
rect 23548 25554 23604 25566
rect 24108 25618 24164 27804
rect 24220 27748 24276 27918
rect 24220 27682 24276 27692
rect 24108 25566 24110 25618
rect 24162 25566 24164 25618
rect 24108 25554 24164 25566
rect 24332 24948 24388 29036
rect 24444 29026 24500 29036
rect 24668 27748 24724 27758
rect 24668 27188 24724 27692
rect 24668 27122 24724 27132
rect 25004 26964 25060 29148
rect 25116 28418 25172 29932
rect 25340 29428 25396 29438
rect 25340 29334 25396 29372
rect 25788 29426 25844 29438
rect 25788 29374 25790 29426
rect 25842 29374 25844 29426
rect 25788 29092 25844 29374
rect 25788 29026 25844 29036
rect 25788 28868 25844 28878
rect 25788 28774 25844 28812
rect 25116 28366 25118 28418
rect 25170 28366 25172 28418
rect 25116 28354 25172 28366
rect 26012 28642 26068 30604
rect 26012 28590 26014 28642
rect 26066 28590 26068 28642
rect 26012 28084 26068 28590
rect 26012 28018 26068 28028
rect 25228 27858 25284 27870
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 25228 27748 25284 27806
rect 25228 27682 25284 27692
rect 25788 27636 25844 27646
rect 25788 27634 25956 27636
rect 25788 27582 25790 27634
rect 25842 27582 25956 27634
rect 25788 27580 25956 27582
rect 25788 27570 25844 27580
rect 25004 26908 25396 26964
rect 25900 26962 25956 27580
rect 25900 26910 25902 26962
rect 25954 26910 25956 26962
rect 25340 26852 25508 26908
rect 25900 26898 25956 26910
rect 25116 26290 25172 26302
rect 25116 26238 25118 26290
rect 25170 26238 25172 26290
rect 24780 26068 24836 26078
rect 24332 24882 24388 24892
rect 24444 26066 24836 26068
rect 24444 26014 24782 26066
rect 24834 26014 24836 26066
rect 24444 26012 24836 26014
rect 23324 24724 23380 24734
rect 23324 23940 23380 24668
rect 23324 23874 23380 23884
rect 24108 24498 24164 24510
rect 24108 24446 24110 24498
rect 24162 24446 24164 24498
rect 24108 23826 24164 24446
rect 24108 23774 24110 23826
rect 24162 23774 24164 23826
rect 24108 23762 24164 23774
rect 24332 23716 24388 23726
rect 24220 23156 24276 23166
rect 22316 20636 22932 20692
rect 22988 22652 23156 22708
rect 24108 23154 24276 23156
rect 24108 23102 24222 23154
rect 24274 23102 24276 23154
rect 24108 23100 24276 23102
rect 22316 16770 22372 20636
rect 22764 19794 22820 19806
rect 22764 19742 22766 19794
rect 22818 19742 22820 19794
rect 22540 19348 22596 19358
rect 22540 19234 22596 19292
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22540 19170 22596 19182
rect 22316 16718 22318 16770
rect 22370 16718 22372 16770
rect 22316 16706 22372 16718
rect 22652 16212 22708 16222
rect 22204 16210 22708 16212
rect 22204 16158 22654 16210
rect 22706 16158 22708 16210
rect 22204 16156 22708 16158
rect 22652 16146 22708 16156
rect 21308 15374 21310 15426
rect 21362 15374 21364 15426
rect 21308 15362 21364 15374
rect 22540 15428 22596 15438
rect 22764 15428 22820 19742
rect 22988 18562 23044 22652
rect 23548 22258 23604 22270
rect 23548 22206 23550 22258
rect 23602 22206 23604 22258
rect 23548 21812 23604 22206
rect 23996 22148 24052 22158
rect 23324 21756 23940 21812
rect 23212 20580 23268 20590
rect 23324 20580 23380 21756
rect 23212 20578 23380 20580
rect 23212 20526 23214 20578
rect 23266 20526 23380 20578
rect 23212 20524 23380 20526
rect 23436 21586 23492 21598
rect 23436 21534 23438 21586
rect 23490 21534 23492 21586
rect 23212 20244 23268 20524
rect 23212 19348 23268 20188
rect 23212 19282 23268 19292
rect 22988 18510 22990 18562
rect 23042 18510 23044 18562
rect 22988 18498 23044 18510
rect 23100 19234 23156 19246
rect 23100 19182 23102 19234
rect 23154 19182 23156 19234
rect 22540 15426 22820 15428
rect 22540 15374 22542 15426
rect 22594 15374 22820 15426
rect 22540 15372 22820 15374
rect 22540 15362 22596 15372
rect 20300 15150 20302 15202
rect 20354 15150 20356 15202
rect 20300 15138 20356 15150
rect 23100 15148 23156 19182
rect 23436 18564 23492 21534
rect 23884 21588 23940 21756
rect 23884 21494 23940 21532
rect 23884 20916 23940 20926
rect 23996 20916 24052 22092
rect 23884 20914 24052 20916
rect 23884 20862 23886 20914
rect 23938 20862 24052 20914
rect 23884 20860 24052 20862
rect 23884 20850 23940 20860
rect 23996 20578 24052 20590
rect 23996 20526 23998 20578
rect 24050 20526 24052 20578
rect 23548 20020 23604 20030
rect 23548 19926 23604 19964
rect 23772 19794 23828 19806
rect 23772 19742 23774 19794
rect 23826 19742 23828 19794
rect 23772 19124 23828 19742
rect 23772 19058 23828 19068
rect 23884 19348 23940 19358
rect 23884 18674 23940 19292
rect 23884 18622 23886 18674
rect 23938 18622 23940 18674
rect 23884 18610 23940 18622
rect 23996 18564 24052 20526
rect 23436 18508 23604 18564
rect 23548 15202 23604 18508
rect 23996 18498 24052 18508
rect 23660 18452 23716 18462
rect 23660 15986 23716 18396
rect 24108 17780 24164 23100
rect 24220 23090 24276 23100
rect 24220 20244 24276 20254
rect 24220 20150 24276 20188
rect 24108 17714 24164 17724
rect 23772 17556 23828 17566
rect 24332 17556 24388 23660
rect 24444 21700 24500 26012
rect 24780 26002 24836 26012
rect 24780 25506 24836 25518
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24556 25284 24612 25294
rect 24780 25284 24836 25454
rect 25116 25284 25172 26238
rect 24556 25282 25116 25284
rect 24556 25230 24558 25282
rect 24610 25230 25116 25282
rect 24556 25228 25116 25230
rect 24556 24724 24612 25228
rect 24556 24658 24612 24668
rect 24668 24836 24724 24846
rect 24668 24722 24724 24780
rect 24668 24670 24670 24722
rect 24722 24670 24724 24722
rect 24668 21700 24724 24670
rect 25004 23940 25060 25228
rect 25116 25190 25172 25228
rect 25228 26292 25284 26302
rect 25228 25060 25284 26236
rect 24780 23938 25060 23940
rect 24780 23886 25006 23938
rect 25058 23886 25060 23938
rect 24780 23884 25060 23886
rect 24780 23156 24836 23884
rect 25004 23874 25060 23884
rect 25116 25004 25284 25060
rect 25340 25506 25396 25518
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 24892 23716 24948 23726
rect 24892 23622 24948 23660
rect 25116 23380 25172 25004
rect 24780 23062 24836 23100
rect 24892 23324 25172 23380
rect 25228 24724 25284 24734
rect 24444 21644 24612 21700
rect 24444 21474 24500 21486
rect 24444 21422 24446 21474
rect 24498 21422 24500 21474
rect 24444 21362 24500 21422
rect 24444 21310 24446 21362
rect 24498 21310 24500 21362
rect 24444 21298 24500 21310
rect 23772 17554 24388 17556
rect 23772 17502 23774 17554
rect 23826 17502 24388 17554
rect 23772 17500 24388 17502
rect 23772 17490 23828 17500
rect 23660 15934 23662 15986
rect 23714 15934 23716 15986
rect 23660 15922 23716 15934
rect 24332 16772 24388 16782
rect 23548 15150 23550 15202
rect 23602 15150 23604 15202
rect 23100 15092 23268 15148
rect 23548 15138 23604 15150
rect 23212 14644 23268 15092
rect 23324 14644 23380 14654
rect 23212 14642 23380 14644
rect 23212 14590 23326 14642
rect 23378 14590 23380 14642
rect 23212 14588 23380 14590
rect 23324 14578 23380 14588
rect 19180 14420 19236 14430
rect 19068 14418 19236 14420
rect 19068 14366 19182 14418
rect 19234 14366 19236 14418
rect 19068 14364 19236 14366
rect 19180 14354 19236 14364
rect 24332 14418 24388 16716
rect 24556 15988 24612 21644
rect 24668 21362 24724 21644
rect 24668 21310 24670 21362
rect 24722 21310 24724 21362
rect 24668 20242 24724 21310
rect 24780 21476 24836 21486
rect 24780 20690 24836 21420
rect 24780 20638 24782 20690
rect 24834 20638 24836 20690
rect 24780 20626 24836 20638
rect 24668 20190 24670 20242
rect 24722 20190 24724 20242
rect 24668 20020 24724 20190
rect 24668 19954 24724 19964
rect 24780 17780 24836 17790
rect 24892 17780 24948 23324
rect 25116 23156 25172 23166
rect 25116 22148 25172 23100
rect 25228 22372 25284 24668
rect 25340 22484 25396 25454
rect 25340 22418 25396 22428
rect 25228 22306 25284 22316
rect 25172 22092 25396 22148
rect 25116 22054 25172 22092
rect 25340 21924 25396 22092
rect 25340 21810 25396 21868
rect 25340 21758 25342 21810
rect 25394 21758 25396 21810
rect 25340 21746 25396 21758
rect 25452 20132 25508 26852
rect 25676 26292 25732 26302
rect 25676 26198 25732 26236
rect 26124 24724 26180 30828
rect 26348 30882 26404 30894
rect 26348 30830 26350 30882
rect 26402 30830 26404 30882
rect 26348 30436 26404 30830
rect 26348 30370 26404 30380
rect 26236 30212 26292 30222
rect 26236 29428 26292 30156
rect 26236 28082 26292 29372
rect 26236 28030 26238 28082
rect 26290 28030 26292 28082
rect 26236 27860 26292 28030
rect 26572 28196 26628 31612
rect 26684 31106 26740 31892
rect 26684 31054 26686 31106
rect 26738 31054 26740 31106
rect 26684 31042 26740 31054
rect 27132 30994 27188 31006
rect 27132 30942 27134 30994
rect 27186 30942 27188 30994
rect 27132 30884 27188 30942
rect 27132 30818 27188 30828
rect 26684 30212 26740 30222
rect 27244 30212 27300 30222
rect 26684 30210 26852 30212
rect 26684 30158 26686 30210
rect 26738 30158 26852 30210
rect 26684 30156 26852 30158
rect 26684 30146 26740 30156
rect 26572 28084 26628 28140
rect 26684 28084 26740 28094
rect 26572 28082 26740 28084
rect 26572 28030 26686 28082
rect 26738 28030 26740 28082
rect 26572 28028 26740 28030
rect 26684 28018 26740 28028
rect 26236 27634 26292 27804
rect 26236 27582 26238 27634
rect 26290 27582 26292 27634
rect 26236 27570 26292 27582
rect 26796 26964 26852 30156
rect 27244 30118 27300 30156
rect 27468 30210 27524 31892
rect 27804 31668 27860 35534
rect 28028 35028 28084 36206
rect 28364 35922 28420 38220
rect 28924 37268 28980 40348
rect 29148 39732 29204 45052
rect 29372 44884 29428 49870
rect 29708 49924 29764 49934
rect 29596 48914 29652 48926
rect 29596 48862 29598 48914
rect 29650 48862 29652 48914
rect 29596 48804 29652 48862
rect 29596 48738 29652 48748
rect 29708 47458 29764 49868
rect 29932 49252 29988 49262
rect 29932 48466 29988 49196
rect 29932 48414 29934 48466
rect 29986 48414 29988 48466
rect 29932 48402 29988 48414
rect 29708 47406 29710 47458
rect 29762 47406 29764 47458
rect 29708 47394 29764 47406
rect 29372 44818 29428 44828
rect 29484 46900 29540 46910
rect 29484 44434 29540 46844
rect 29820 45780 29876 45790
rect 29820 45686 29876 45724
rect 29484 44382 29486 44434
rect 29538 44382 29540 44434
rect 29484 44370 29540 44382
rect 29820 44436 29876 44446
rect 29820 44342 29876 44380
rect 29260 42756 29316 42766
rect 29260 42662 29316 42700
rect 29708 42756 29764 42766
rect 30044 42756 30100 51212
rect 30156 51202 30212 51212
rect 30268 48914 30324 48926
rect 30268 48862 30270 48914
rect 30322 48862 30324 48914
rect 30156 48802 30212 48814
rect 30156 48750 30158 48802
rect 30210 48750 30212 48802
rect 30156 47236 30212 48750
rect 30268 48804 30324 48862
rect 30716 48916 30772 51998
rect 31052 49924 31108 52782
rect 31052 49858 31108 49868
rect 30716 48850 30772 48860
rect 31052 49698 31108 49710
rect 31052 49646 31054 49698
rect 31106 49646 31108 49698
rect 30268 48244 30324 48748
rect 30268 48178 30324 48188
rect 30828 48244 30884 48254
rect 30828 48150 30884 48188
rect 30156 47170 30212 47180
rect 30940 48130 30996 48142
rect 30940 48078 30942 48130
rect 30994 48078 30996 48130
rect 30940 46898 30996 48078
rect 30940 46846 30942 46898
rect 30994 46846 30996 46898
rect 30940 46834 30996 46846
rect 30940 45108 30996 45118
rect 30940 45014 30996 45052
rect 30492 44322 30548 44334
rect 30492 44270 30494 44322
rect 30546 44270 30548 44322
rect 29708 42754 30100 42756
rect 29708 42702 29710 42754
rect 29762 42702 30100 42754
rect 29708 42700 30100 42702
rect 30268 44210 30324 44222
rect 30268 44158 30270 44210
rect 30322 44158 30324 44210
rect 29708 42690 29764 42700
rect 30268 42308 30324 44158
rect 30268 42242 30324 42252
rect 29148 39620 29204 39676
rect 29372 42084 29428 42094
rect 29148 39618 29316 39620
rect 29148 39566 29150 39618
rect 29202 39566 29316 39618
rect 29148 39564 29316 39566
rect 29148 39554 29204 39564
rect 29148 37940 29204 37950
rect 28924 37266 29092 37268
rect 28924 37214 28926 37266
rect 28978 37214 29092 37266
rect 28924 37212 29092 37214
rect 28924 37202 28980 37212
rect 29036 36482 29092 37212
rect 29036 36430 29038 36482
rect 29090 36430 29092 36482
rect 29036 36418 29092 36430
rect 28364 35870 28366 35922
rect 28418 35870 28420 35922
rect 28364 35858 28420 35870
rect 29148 35922 29204 37884
rect 29148 35870 29150 35922
rect 29202 35870 29204 35922
rect 29148 35858 29204 35870
rect 28028 34692 28084 34972
rect 28476 34804 28532 34814
rect 28364 34692 28420 34702
rect 28028 34690 28420 34692
rect 28028 34638 28366 34690
rect 28418 34638 28420 34690
rect 28028 34636 28420 34638
rect 28364 34130 28420 34636
rect 28364 34078 28366 34130
rect 28418 34078 28420 34130
rect 28364 31948 28420 34078
rect 28476 33346 28532 34748
rect 29260 34690 29316 39564
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 28476 33294 28478 33346
rect 28530 33294 28532 33346
rect 28476 33282 28532 33294
rect 28700 34130 28756 34142
rect 28700 34078 28702 34130
rect 28754 34078 28756 34130
rect 28700 33012 28756 34078
rect 28700 32946 28756 32956
rect 28476 32564 28532 32574
rect 28476 32470 28532 32508
rect 28700 32338 28756 32350
rect 28700 32286 28702 32338
rect 28754 32286 28756 32338
rect 28140 31892 28196 31902
rect 28364 31892 28644 31948
rect 28140 31778 28196 31836
rect 28140 31726 28142 31778
rect 28194 31726 28196 31778
rect 28140 31714 28196 31726
rect 28588 31778 28644 31892
rect 28588 31726 28590 31778
rect 28642 31726 28644 31778
rect 27804 31602 27860 31612
rect 28588 31220 28644 31726
rect 28588 31154 28644 31164
rect 27468 30158 27470 30210
rect 27522 30158 27524 30210
rect 27468 30146 27524 30158
rect 28252 30212 28308 30222
rect 28252 30118 28308 30156
rect 27580 29988 27636 29998
rect 27580 29894 27636 29932
rect 28140 29650 28196 29662
rect 28140 29598 28142 29650
rect 28194 29598 28196 29650
rect 27244 28084 27300 28094
rect 27300 28028 27412 28084
rect 27244 27990 27300 28028
rect 27020 27634 27076 27646
rect 27020 27582 27022 27634
rect 27074 27582 27076 27634
rect 27020 27186 27076 27582
rect 27020 27134 27022 27186
rect 27074 27134 27076 27186
rect 27020 27122 27076 27134
rect 26796 26908 27188 26964
rect 26684 26852 26740 26862
rect 26684 26758 26740 26796
rect 26124 24658 26180 24668
rect 25676 23940 25732 23950
rect 25676 23938 25844 23940
rect 25676 23886 25678 23938
rect 25730 23886 25844 23938
rect 25676 23884 25844 23886
rect 25676 23874 25732 23884
rect 25676 23154 25732 23166
rect 25676 23102 25678 23154
rect 25730 23102 25732 23154
rect 25676 20580 25732 23102
rect 25788 22036 25844 23884
rect 27020 22594 27076 22606
rect 27020 22542 27022 22594
rect 27074 22542 27076 22594
rect 25788 21970 25844 21980
rect 26460 22484 26516 22494
rect 25788 21700 25844 21710
rect 25788 21586 25844 21644
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25788 21522 25844 21534
rect 25900 21476 25956 21486
rect 25900 21382 25956 21420
rect 25676 20524 26180 20580
rect 26012 20132 26068 20142
rect 25452 20130 26068 20132
rect 25452 20078 26014 20130
rect 26066 20078 26068 20130
rect 25452 20076 26068 20078
rect 26012 20066 26068 20076
rect 25340 20020 25396 20030
rect 25340 19908 25396 19964
rect 25452 19908 25508 19918
rect 25340 19906 25508 19908
rect 25340 19854 25454 19906
rect 25506 19854 25508 19906
rect 25340 19852 25508 19854
rect 25452 19842 25508 19852
rect 25452 19124 25508 19134
rect 25452 19030 25508 19068
rect 26124 18228 26180 20524
rect 26236 19012 26292 19022
rect 26236 19010 26404 19012
rect 26236 18958 26238 19010
rect 26290 18958 26404 19010
rect 26236 18956 26404 18958
rect 26236 18946 26292 18956
rect 26124 18162 26180 18172
rect 24780 17778 24948 17780
rect 24780 17726 24782 17778
rect 24834 17726 24948 17778
rect 24780 17724 24948 17726
rect 24780 17714 24836 17724
rect 24556 15922 24612 15932
rect 24332 14366 24334 14418
rect 24386 14366 24388 14418
rect 24332 14354 24388 14366
rect 26348 14418 26404 18956
rect 26460 16210 26516 22428
rect 27020 22482 27076 22542
rect 27020 22430 27022 22482
rect 27074 22430 27076 22482
rect 27020 22418 27076 22430
rect 26908 22372 26964 22382
rect 26908 21810 26964 22316
rect 26908 21758 26910 21810
rect 26962 21758 26964 21810
rect 26908 21746 26964 21758
rect 27020 20802 27076 20814
rect 27020 20750 27022 20802
rect 27074 20750 27076 20802
rect 26572 19348 26628 19358
rect 26572 19254 26628 19292
rect 26460 16158 26462 16210
rect 26514 16158 26516 16210
rect 26460 16146 26516 16158
rect 27020 14644 27076 20750
rect 27132 19906 27188 26908
rect 27132 19854 27134 19906
rect 27186 19854 27188 19906
rect 27132 19842 27188 19854
rect 27244 24948 27300 24958
rect 27132 17780 27188 17790
rect 27244 17780 27300 24892
rect 27356 22596 27412 28028
rect 27468 27636 27524 27646
rect 27468 27542 27524 27580
rect 28140 27188 28196 29598
rect 28364 28756 28420 28766
rect 28364 28754 28644 28756
rect 28364 28702 28366 28754
rect 28418 28702 28644 28754
rect 28364 28700 28644 28702
rect 28364 28690 28420 28700
rect 28252 28644 28308 28654
rect 28252 28082 28308 28588
rect 28252 28030 28254 28082
rect 28306 28030 28308 28082
rect 28252 28018 28308 28030
rect 28588 28532 28644 28700
rect 28252 27188 28308 27198
rect 28140 27186 28308 27188
rect 28140 27134 28254 27186
rect 28306 27134 28308 27186
rect 28140 27132 28308 27134
rect 28252 27122 28308 27132
rect 28588 27186 28644 28476
rect 28588 27134 28590 27186
rect 28642 27134 28644 27186
rect 28028 27076 28084 27086
rect 27468 26964 27524 26974
rect 27916 26964 27972 26974
rect 27468 26962 27972 26964
rect 27468 26910 27470 26962
rect 27522 26910 27918 26962
rect 27970 26910 27972 26962
rect 27468 26908 27972 26910
rect 27468 25284 27524 26908
rect 27916 26898 27972 26908
rect 27468 25218 27524 25228
rect 27916 25282 27972 25294
rect 27916 25230 27918 25282
rect 27970 25230 27972 25282
rect 27916 24052 27972 25230
rect 27916 23986 27972 23996
rect 27356 22502 27412 22540
rect 27916 23156 27972 23166
rect 27468 22484 27524 22494
rect 27916 22484 27972 23100
rect 27468 22482 27972 22484
rect 27468 22430 27470 22482
rect 27522 22430 27918 22482
rect 27970 22430 27972 22482
rect 27468 22428 27972 22430
rect 27132 17778 27300 17780
rect 27132 17726 27134 17778
rect 27186 17726 27300 17778
rect 27132 17724 27300 17726
rect 27356 22036 27412 22046
rect 27132 17714 27188 17724
rect 27356 16772 27412 21980
rect 27468 21924 27524 22428
rect 27916 22418 27972 22428
rect 27468 20916 27524 21868
rect 27580 21588 27636 21598
rect 27804 21588 27860 21598
rect 27636 21586 27860 21588
rect 27636 21534 27806 21586
rect 27858 21534 27860 21586
rect 27636 21532 27860 21534
rect 27580 21494 27636 21532
rect 27804 21522 27860 21532
rect 28028 21140 28084 27020
rect 28364 26852 28420 26862
rect 28252 26516 28308 26526
rect 28252 26422 28308 26460
rect 28140 25396 28196 25406
rect 28140 23714 28196 25340
rect 28140 23662 28142 23714
rect 28194 23662 28196 23714
rect 28140 23650 28196 23662
rect 28252 23378 28308 23390
rect 28252 23326 28254 23378
rect 28306 23326 28308 23378
rect 28252 22482 28308 23326
rect 28252 22430 28254 22482
rect 28306 22430 28308 22482
rect 28252 22418 28308 22430
rect 28028 21084 28308 21140
rect 28140 20916 28196 20926
rect 27468 20914 28196 20916
rect 27468 20862 28142 20914
rect 28194 20862 28196 20914
rect 27468 20860 28196 20862
rect 27468 20802 27524 20860
rect 28140 20850 28196 20860
rect 27468 20750 27470 20802
rect 27522 20750 27524 20802
rect 27468 20738 27524 20750
rect 28252 20692 28308 21084
rect 27804 20636 28308 20692
rect 27804 18338 27860 20636
rect 27804 18286 27806 18338
rect 27858 18286 27860 18338
rect 27804 18274 27860 18286
rect 28252 17780 28308 17790
rect 27468 16772 27524 16782
rect 27356 16770 27524 16772
rect 27356 16718 27470 16770
rect 27522 16718 27524 16770
rect 27356 16716 27524 16718
rect 27468 16706 27524 16716
rect 27244 15988 27300 15998
rect 27244 15894 27300 15932
rect 28252 15202 28308 17724
rect 28364 17554 28420 26796
rect 28588 26740 28644 27134
rect 28588 26674 28644 26684
rect 28476 25282 28532 25294
rect 28476 25230 28478 25282
rect 28530 25230 28532 25282
rect 28476 23604 28532 25230
rect 28700 24276 28756 32286
rect 29260 31948 29316 34638
rect 29036 31892 29316 31948
rect 29372 31892 29428 42028
rect 29484 41076 29540 41086
rect 29484 40402 29540 41020
rect 29484 40350 29486 40402
rect 29538 40350 29540 40402
rect 29484 40338 29540 40350
rect 29932 41074 29988 41086
rect 29932 41022 29934 41074
rect 29986 41022 29988 41074
rect 29932 39844 29988 41022
rect 30492 40516 30548 44270
rect 31052 43538 31108 49646
rect 31388 49252 31444 53566
rect 32060 53060 32116 53070
rect 31388 49186 31444 49196
rect 31500 53058 32116 53060
rect 31500 53006 32062 53058
rect 32114 53006 32116 53058
rect 31500 53004 32116 53006
rect 31052 43486 31054 43538
rect 31106 43486 31108 43538
rect 31052 43474 31108 43486
rect 31164 48356 31220 48366
rect 30604 42082 30660 42094
rect 30604 42030 30606 42082
rect 30658 42030 30660 42082
rect 30604 40740 30660 42030
rect 31164 41748 31220 48300
rect 31500 46900 31556 53004
rect 32060 52994 32116 53004
rect 32060 52276 32116 52286
rect 33404 52276 33460 52286
rect 32060 52274 32228 52276
rect 32060 52222 32062 52274
rect 32114 52222 32228 52274
rect 32060 52220 32228 52222
rect 32060 52210 32116 52220
rect 32060 49924 32116 49934
rect 31836 49922 32116 49924
rect 31836 49870 32062 49922
rect 32114 49870 32116 49922
rect 31836 49868 32116 49870
rect 31724 49026 31780 49038
rect 31724 48974 31726 49026
rect 31778 48974 31780 49026
rect 31612 48130 31668 48142
rect 31612 48078 31614 48130
rect 31666 48078 31668 48130
rect 31612 47124 31668 48078
rect 31724 47460 31780 48974
rect 31724 47394 31780 47404
rect 31612 47068 31780 47124
rect 31612 46900 31668 46910
rect 31500 46898 31668 46900
rect 31500 46846 31614 46898
rect 31666 46846 31668 46898
rect 31500 46844 31668 46846
rect 31612 46834 31668 46844
rect 31724 45780 31780 47068
rect 31724 45714 31780 45724
rect 31500 44324 31556 44334
rect 31388 43540 31444 43550
rect 31500 43540 31556 44268
rect 31388 43538 31556 43540
rect 31388 43486 31390 43538
rect 31442 43486 31556 43538
rect 31388 43484 31556 43486
rect 31388 42756 31444 43484
rect 31388 42690 31444 42700
rect 31836 42532 31892 49868
rect 32060 49858 32116 49868
rect 32060 49028 32116 49038
rect 32060 48934 32116 48972
rect 31948 48244 32004 48254
rect 31948 48150 32004 48188
rect 32172 47908 32228 52220
rect 32956 52052 33012 52062
rect 32620 50706 32676 50718
rect 32620 50654 32622 50706
rect 32674 50654 32676 50706
rect 32620 48356 32676 50654
rect 32620 48290 32676 48300
rect 32732 48916 32788 48926
rect 31948 47852 32228 47908
rect 32284 48244 32340 48254
rect 31948 45892 32004 47852
rect 32060 47234 32116 47246
rect 32060 47182 32062 47234
rect 32114 47182 32116 47234
rect 32060 46116 32116 47182
rect 32284 46674 32340 48188
rect 32284 46622 32286 46674
rect 32338 46622 32340 46674
rect 32060 46060 32228 46116
rect 32060 45892 32116 45902
rect 31948 45890 32116 45892
rect 31948 45838 32062 45890
rect 32114 45838 32116 45890
rect 31948 45836 32116 45838
rect 32060 45826 32116 45836
rect 32060 45668 32116 45678
rect 32060 44322 32116 45612
rect 32172 45218 32228 46060
rect 32172 45166 32174 45218
rect 32226 45166 32228 45218
rect 32172 45154 32228 45166
rect 32284 45108 32340 46622
rect 32620 48132 32676 48142
rect 32508 46562 32564 46574
rect 32508 46510 32510 46562
rect 32562 46510 32564 46562
rect 32508 45332 32564 46510
rect 32620 45444 32676 48076
rect 32732 47682 32788 48860
rect 32732 47630 32734 47682
rect 32786 47630 32788 47682
rect 32732 47618 32788 47630
rect 32844 47460 32900 47470
rect 32844 47012 32900 47404
rect 32732 46956 32900 47012
rect 32732 45890 32788 46956
rect 32732 45838 32734 45890
rect 32786 45838 32788 45890
rect 32732 45826 32788 45838
rect 32844 45890 32900 45902
rect 32844 45838 32846 45890
rect 32898 45838 32900 45890
rect 32620 45388 32788 45444
rect 32508 45266 32564 45276
rect 32396 45108 32452 45118
rect 32732 45108 32788 45388
rect 32284 45106 32452 45108
rect 32284 45054 32398 45106
rect 32450 45054 32452 45106
rect 32284 45052 32452 45054
rect 32284 44436 32340 45052
rect 32396 45042 32452 45052
rect 32508 45052 32788 45108
rect 32284 44370 32340 44380
rect 32060 44270 32062 44322
rect 32114 44270 32116 44322
rect 32060 44258 32116 44270
rect 32396 43538 32452 43550
rect 32396 43486 32398 43538
rect 32450 43486 32452 43538
rect 31388 42476 31892 42532
rect 32172 43426 32228 43438
rect 32172 43374 32174 43426
rect 32226 43374 32228 43426
rect 32172 42530 32228 43374
rect 32172 42478 32174 42530
rect 32226 42478 32228 42530
rect 31388 41970 31444 42476
rect 32172 42466 32228 42478
rect 32396 43428 32452 43486
rect 31388 41918 31390 41970
rect 31442 41918 31444 41970
rect 31388 41906 31444 41918
rect 31724 41970 31780 41982
rect 31724 41918 31726 41970
rect 31778 41918 31780 41970
rect 31164 41682 31220 41692
rect 30604 40674 30660 40684
rect 30940 41298 30996 41310
rect 30940 41246 30942 41298
rect 30994 41246 30996 41298
rect 30604 40516 30660 40526
rect 30492 40460 30604 40516
rect 30604 40450 30660 40460
rect 30940 39956 30996 41246
rect 31724 40516 31780 41918
rect 31836 41858 31892 41870
rect 31836 41806 31838 41858
rect 31890 41806 31892 41858
rect 31836 40626 31892 41806
rect 32396 41748 32452 43372
rect 32508 42084 32564 45052
rect 32620 44884 32676 44894
rect 32620 42756 32676 44828
rect 32844 44324 32900 45838
rect 32956 45330 33012 51996
rect 33404 50428 33460 52220
rect 33292 50372 33460 50428
rect 33180 49924 33236 49934
rect 33068 48242 33124 48254
rect 33068 48190 33070 48242
rect 33122 48190 33124 48242
rect 33068 48132 33124 48190
rect 33068 48066 33124 48076
rect 32956 45278 32958 45330
rect 33010 45278 33012 45330
rect 32956 45266 33012 45278
rect 32844 44258 32900 44268
rect 33068 43652 33124 43662
rect 33068 43558 33124 43596
rect 33180 43428 33236 49868
rect 33292 45892 33348 50372
rect 33404 49028 33460 49038
rect 33516 49028 33572 53788
rect 33628 53778 33684 53788
rect 37436 53842 38612 53844
rect 37436 53790 38558 53842
rect 38610 53790 38612 53842
rect 37436 53788 38612 53790
rect 34636 53618 34692 53630
rect 34636 53566 34638 53618
rect 34690 53566 34692 53618
rect 34412 52276 34468 52286
rect 34412 52182 34468 52220
rect 33964 50482 34020 50494
rect 33964 50430 33966 50482
rect 34018 50430 34020 50482
rect 33964 50428 34020 50430
rect 33460 48972 33572 49028
rect 33852 50372 34020 50428
rect 33404 48962 33460 48972
rect 33516 48804 33572 48814
rect 33516 47458 33572 48748
rect 33516 47406 33518 47458
rect 33570 47406 33572 47458
rect 33516 47394 33572 47406
rect 33404 45892 33460 45902
rect 33292 45890 33460 45892
rect 33292 45838 33406 45890
rect 33458 45838 33460 45890
rect 33292 45836 33460 45838
rect 33404 45826 33460 45836
rect 33740 45332 33796 45342
rect 33740 45238 33796 45276
rect 33740 44436 33796 44446
rect 33628 44100 33684 44110
rect 32732 43372 33236 43428
rect 33292 43538 33348 43550
rect 33292 43486 33294 43538
rect 33346 43486 33348 43538
rect 33292 43428 33348 43486
rect 32732 42978 32788 43372
rect 33292 43362 33348 43372
rect 32732 42926 32734 42978
rect 32786 42926 32788 42978
rect 32732 42914 32788 42926
rect 32844 42756 32900 42766
rect 32620 42754 32900 42756
rect 32620 42702 32846 42754
rect 32898 42702 32900 42754
rect 32620 42700 32900 42702
rect 32844 42690 32900 42700
rect 33628 42642 33684 44044
rect 33740 43428 33796 44380
rect 33852 43652 33908 50372
rect 34076 49700 34132 49710
rect 33964 49698 34132 49700
rect 33964 49646 34078 49698
rect 34130 49646 34132 49698
rect 33964 49644 34132 49646
rect 33964 45668 34020 49644
rect 34076 49634 34132 49644
rect 34636 48916 34692 53566
rect 37324 53620 37380 53630
rect 35868 53058 35924 53070
rect 35868 53006 35870 53058
rect 35922 53006 35924 53058
rect 34636 48850 34692 48860
rect 34860 52834 34916 52846
rect 34860 52782 34862 52834
rect 34914 52782 34916 52834
rect 34412 48804 34468 48814
rect 33964 45602 34020 45612
rect 34188 48802 34468 48804
rect 34188 48750 34414 48802
rect 34466 48750 34468 48802
rect 34188 48748 34468 48750
rect 33852 43596 34020 43652
rect 33852 43428 33908 43438
rect 33740 43426 33908 43428
rect 33740 43374 33854 43426
rect 33906 43374 33908 43426
rect 33740 43372 33908 43374
rect 33852 43362 33908 43372
rect 33628 42590 33630 42642
rect 33682 42590 33684 42642
rect 33628 42578 33684 42590
rect 32508 42028 32788 42084
rect 32508 41970 32564 42028
rect 32508 41918 32510 41970
rect 32562 41918 32564 41970
rect 32508 41906 32564 41918
rect 32732 41972 32788 42028
rect 33292 41972 33348 41982
rect 32732 41970 33348 41972
rect 32732 41918 33294 41970
rect 33346 41918 33348 41970
rect 32732 41916 33348 41918
rect 31836 40574 31838 40626
rect 31890 40574 31892 40626
rect 31836 40562 31892 40574
rect 32172 41186 32228 41198
rect 32172 41134 32174 41186
rect 32226 41134 32228 41186
rect 31724 40450 31780 40460
rect 30940 39890 30996 39900
rect 31164 40404 31220 40414
rect 29932 39778 29988 39788
rect 31164 39732 31220 40348
rect 31948 40404 32004 40414
rect 32172 40404 32228 41134
rect 32004 40348 32228 40404
rect 31948 40338 32004 40348
rect 32172 40292 32228 40348
rect 32172 40226 32228 40236
rect 32284 40516 32340 40526
rect 32396 40516 32452 41692
rect 32620 41860 32676 41870
rect 32620 40626 32676 41804
rect 32732 41188 32788 41198
rect 32732 41094 32788 41132
rect 32620 40574 32622 40626
rect 32674 40574 32676 40626
rect 32620 40562 32676 40574
rect 32340 40460 32452 40516
rect 32060 39956 32116 39966
rect 31164 39730 31444 39732
rect 31164 39678 31166 39730
rect 31218 39678 31444 39730
rect 31164 39676 31444 39678
rect 31164 39666 31220 39676
rect 31164 38836 31220 38846
rect 31164 38742 31220 38780
rect 31388 38836 31444 39676
rect 31948 38948 32004 38958
rect 31948 38854 32004 38892
rect 31500 38836 31556 38846
rect 31388 38834 31556 38836
rect 31388 38782 31502 38834
rect 31554 38782 31556 38834
rect 31388 38780 31556 38782
rect 30940 38164 30996 38174
rect 30828 37940 30884 37950
rect 30828 37846 30884 37884
rect 29484 37268 29540 37278
rect 29484 37174 29540 37212
rect 29596 36932 29652 36942
rect 29596 36482 29652 36876
rect 29596 36430 29598 36482
rect 29650 36430 29652 36482
rect 29596 36418 29652 36430
rect 29932 36260 29988 36270
rect 29932 35028 29988 36204
rect 29932 35026 30212 35028
rect 29932 34974 29934 35026
rect 29986 34974 30212 35026
rect 29932 34972 30212 34974
rect 29932 34962 29988 34972
rect 30156 34914 30212 34972
rect 30156 34862 30158 34914
rect 30210 34862 30212 34914
rect 30156 34850 30212 34862
rect 30604 33348 30660 33358
rect 30604 33254 30660 33292
rect 30940 33346 30996 38108
rect 31388 38050 31444 38780
rect 31500 38770 31556 38780
rect 31388 37998 31390 38050
rect 31442 37998 31444 38050
rect 31388 37986 31444 37998
rect 31948 38052 32004 38062
rect 32060 38052 32116 39900
rect 32284 38946 32340 40460
rect 32284 38894 32286 38946
rect 32338 38894 32340 38946
rect 32284 38882 32340 38894
rect 32620 39844 32676 39854
rect 31948 38050 32116 38052
rect 31948 37998 31950 38050
rect 32002 37998 32116 38050
rect 31948 37996 32116 37998
rect 31948 37986 32004 37996
rect 31164 37940 31220 37950
rect 31164 37846 31220 37884
rect 32620 37490 32676 39788
rect 33292 38948 33348 41916
rect 33964 40628 34020 43596
rect 34188 43650 34244 48748
rect 34412 48738 34468 48748
rect 34860 48804 34916 52782
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35756 52276 35812 52286
rect 35644 52220 35756 52276
rect 35420 52052 35476 52062
rect 35420 51958 35476 51996
rect 34860 48738 34916 48748
rect 34972 51492 35028 51502
rect 34188 43598 34190 43650
rect 34242 43598 34244 43650
rect 34188 43586 34244 43598
rect 34300 46562 34356 46574
rect 34300 46510 34302 46562
rect 34354 46510 34356 46562
rect 34076 41748 34132 41758
rect 34076 41654 34132 41692
rect 33964 40562 34020 40572
rect 33516 40402 33572 40414
rect 33516 40350 33518 40402
rect 33570 40350 33572 40402
rect 33516 40292 33572 40350
rect 34188 40404 34244 40414
rect 34300 40404 34356 46510
rect 34972 44548 35028 51436
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 50820 35252 50830
rect 35196 49588 35252 50764
rect 35308 49924 35364 49934
rect 35308 49830 35364 49868
rect 35084 49532 35252 49588
rect 35084 49252 35140 49532
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 49252 35252 49262
rect 35084 49250 35252 49252
rect 35084 49198 35198 49250
rect 35250 49198 35252 49250
rect 35084 49196 35252 49198
rect 35196 49186 35252 49196
rect 35420 48244 35476 48254
rect 35420 48130 35476 48188
rect 35420 48078 35422 48130
rect 35474 48078 35476 48130
rect 35420 48066 35476 48078
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35420 46788 35476 46798
rect 35420 46786 35588 46788
rect 35420 46734 35422 46786
rect 35474 46734 35588 46786
rect 35420 46732 35588 46734
rect 35420 46722 35476 46732
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 44548 35252 44558
rect 34972 44546 35252 44548
rect 34972 44494 35198 44546
rect 35250 44494 35252 44546
rect 34972 44492 35252 44494
rect 35196 44482 35252 44492
rect 34636 44100 34692 44110
rect 34636 44098 34804 44100
rect 34636 44046 34638 44098
rect 34690 44046 34804 44098
rect 34636 44044 34804 44046
rect 34636 44034 34692 44044
rect 34188 40402 34356 40404
rect 34188 40350 34190 40402
rect 34242 40350 34356 40402
rect 34188 40348 34356 40350
rect 34188 40338 34244 40348
rect 34524 40292 34580 40302
rect 33572 40236 33908 40292
rect 33516 40226 33572 40236
rect 33292 38724 33348 38892
rect 33852 38834 33908 40236
rect 33852 38782 33854 38834
rect 33906 38782 33908 38834
rect 33852 38770 33908 38782
rect 34524 38834 34580 40236
rect 34748 39730 34804 44044
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34748 39678 34750 39730
rect 34802 39678 34804 39730
rect 34748 39666 34804 39678
rect 34972 41748 35028 41758
rect 34972 39618 35028 41692
rect 35532 41636 35588 46732
rect 35644 45108 35700 52220
rect 35756 52210 35812 52220
rect 35868 50820 35924 53006
rect 36652 53060 36708 53070
rect 35868 50754 35924 50764
rect 36428 52836 36484 52846
rect 36316 49924 36372 49934
rect 36092 49028 36148 49038
rect 36092 49026 36260 49028
rect 36092 48974 36094 49026
rect 36146 48974 36260 49026
rect 36092 48972 36260 48974
rect 36092 48962 36148 48972
rect 36092 48802 36148 48814
rect 36092 48750 36094 48802
rect 36146 48750 36148 48802
rect 36092 48692 36148 48750
rect 35756 48636 36148 48692
rect 35756 45778 35812 48636
rect 36092 48468 36148 48478
rect 35868 48466 36148 48468
rect 35868 48414 36094 48466
rect 36146 48414 36148 48466
rect 35868 48412 36148 48414
rect 35868 47234 35924 48412
rect 36092 48402 36148 48412
rect 36092 48244 36148 48254
rect 36204 48244 36260 48972
rect 36148 48188 36260 48244
rect 36092 48150 36148 48188
rect 35868 47182 35870 47234
rect 35922 47182 35924 47234
rect 35868 47170 35924 47182
rect 35980 47460 36036 47470
rect 35980 46674 36036 47404
rect 35980 46622 35982 46674
rect 36034 46622 36036 46674
rect 35980 46610 36036 46622
rect 36316 46004 36372 49868
rect 36428 46674 36484 52780
rect 36540 49588 36596 49598
rect 36540 47682 36596 49532
rect 36540 47630 36542 47682
rect 36594 47630 36596 47682
rect 36540 47618 36596 47630
rect 36428 46622 36430 46674
rect 36482 46622 36484 46674
rect 36428 46610 36484 46622
rect 36540 46116 36596 46126
rect 36652 46116 36708 53004
rect 36764 51268 36820 51278
rect 36764 51266 36932 51268
rect 36764 51214 36766 51266
rect 36818 51214 36932 51266
rect 36764 51212 36932 51214
rect 36764 51202 36820 51212
rect 36764 48244 36820 48254
rect 36764 47460 36820 48188
rect 36764 47394 36820 47404
rect 36540 46114 36708 46116
rect 36540 46062 36542 46114
rect 36594 46062 36708 46114
rect 36540 46060 36708 46062
rect 36540 46050 36596 46060
rect 35756 45726 35758 45778
rect 35810 45726 35812 45778
rect 35756 45714 35812 45726
rect 36092 45948 36372 46004
rect 35980 45108 36036 45118
rect 35644 45106 36036 45108
rect 35644 45054 35982 45106
rect 36034 45054 36036 45106
rect 35644 45052 36036 45054
rect 35980 45042 36036 45052
rect 36092 44884 36148 45948
rect 36876 45892 36932 51212
rect 36988 49924 37044 49934
rect 36988 49830 37044 49868
rect 37324 46116 37380 53564
rect 37436 48242 37492 53788
rect 38556 53778 38612 53788
rect 40348 53842 41412 53844
rect 40348 53790 41358 53842
rect 41410 53790 41412 53842
rect 40348 53788 41412 53790
rect 39564 53620 39620 53630
rect 39564 53526 39620 53564
rect 38668 53060 38724 53070
rect 38668 52966 38724 53004
rect 37660 52836 37716 52846
rect 37660 52742 37716 52780
rect 37996 52276 38052 52286
rect 37996 52182 38052 52220
rect 39452 52276 39508 52286
rect 39116 52050 39172 52062
rect 39116 51998 39118 52050
rect 39170 51998 39172 52050
rect 37772 51492 37828 51502
rect 37772 51398 37828 51436
rect 39004 50708 39060 50718
rect 38220 50596 38276 50606
rect 38108 49700 38164 49710
rect 37436 48190 37438 48242
rect 37490 48190 37492 48242
rect 37436 48178 37492 48190
rect 37548 49698 38164 49700
rect 37548 49646 38110 49698
rect 38162 49646 38164 49698
rect 37548 49644 38164 49646
rect 37436 46116 37492 46126
rect 37324 46114 37492 46116
rect 37324 46062 37438 46114
rect 37490 46062 37492 46114
rect 37324 46060 37492 46062
rect 37436 46050 37492 46060
rect 35868 44828 36148 44884
rect 36204 45836 36932 45892
rect 35868 41970 35924 44828
rect 35980 44210 36036 44222
rect 35980 44158 35982 44210
rect 36034 44158 36036 44210
rect 35980 44100 36036 44158
rect 35980 44034 36036 44044
rect 35980 42756 36036 42766
rect 36204 42756 36260 45836
rect 36428 45108 36484 45118
rect 36764 45108 36820 45118
rect 36428 45106 36820 45108
rect 36428 45054 36430 45106
rect 36482 45054 36766 45106
rect 36818 45054 36820 45106
rect 36428 45052 36820 45054
rect 36428 44324 36484 45052
rect 36764 45042 36820 45052
rect 37436 45108 37492 45118
rect 37436 45014 37492 45052
rect 37548 44548 37604 49644
rect 38108 49634 38164 49644
rect 37996 49026 38052 49038
rect 37996 48974 37998 49026
rect 38050 48974 38052 49026
rect 37996 48244 38052 48974
rect 37996 48178 38052 48188
rect 38220 47460 38276 50540
rect 38892 50484 38948 50494
rect 37324 44492 37604 44548
rect 37660 47404 38276 47460
rect 38332 50482 38948 50484
rect 38332 50430 38894 50482
rect 38946 50430 38948 50482
rect 38332 50428 38948 50430
rect 35980 42754 36260 42756
rect 35980 42702 35982 42754
rect 36034 42702 36260 42754
rect 35980 42700 36260 42702
rect 36316 44210 36372 44222
rect 36316 44158 36318 44210
rect 36370 44158 36372 44210
rect 35980 42690 36036 42700
rect 36316 42644 36372 44158
rect 36428 42756 36484 44268
rect 36988 44324 37044 44334
rect 36988 44230 37044 44268
rect 36540 43540 36596 43550
rect 36540 43446 36596 43484
rect 36876 42756 36932 42766
rect 36428 42754 36876 42756
rect 36428 42702 36430 42754
rect 36482 42702 36876 42754
rect 36428 42700 36876 42702
rect 37324 42756 37380 44492
rect 37436 44324 37492 44334
rect 37660 44324 37716 47404
rect 38220 47236 38276 47246
rect 38220 45778 38276 47180
rect 38220 45726 38222 45778
rect 38274 45726 38276 45778
rect 38220 45714 38276 45726
rect 38332 44884 38388 50428
rect 38892 50418 38948 50428
rect 38668 49028 38724 49038
rect 39004 49028 39060 50652
rect 39116 49588 39172 51998
rect 39116 49522 39172 49532
rect 38668 49026 39060 49028
rect 38668 48974 38670 49026
rect 38722 48974 39060 49026
rect 38668 48972 39060 48974
rect 39116 49028 39172 49038
rect 38668 48962 38724 48972
rect 38892 48132 38948 48142
rect 38892 46898 38948 48076
rect 38892 46846 38894 46898
rect 38946 46846 38948 46898
rect 38892 46834 38948 46846
rect 37436 44322 37716 44324
rect 37436 44270 37438 44322
rect 37490 44270 37716 44322
rect 37436 44268 37716 44270
rect 37772 44828 38388 44884
rect 37436 44258 37492 44268
rect 37660 43988 37716 43998
rect 37436 42756 37492 42766
rect 37324 42754 37492 42756
rect 37324 42702 37438 42754
rect 37490 42702 37492 42754
rect 37324 42700 37492 42702
rect 36428 42690 36484 42700
rect 36876 42662 36932 42700
rect 37436 42690 37492 42700
rect 35868 41918 35870 41970
rect 35922 41918 35924 41970
rect 35868 41906 35924 41918
rect 36092 42588 36372 42644
rect 36092 41748 36148 42588
rect 35196 41580 35460 41590
rect 35532 41580 35812 41636
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35756 41412 35812 41580
rect 35868 41412 35924 41422
rect 35756 41410 35924 41412
rect 35756 41358 35870 41410
rect 35922 41358 35924 41410
rect 35756 41356 35924 41358
rect 35868 41346 35924 41356
rect 36092 41298 36148 41692
rect 36092 41246 36094 41298
rect 36146 41246 36148 41298
rect 36092 41234 36148 41246
rect 36316 42084 36372 42094
rect 35196 40964 35252 40974
rect 35196 40870 35252 40908
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34972 39566 34974 39618
rect 35026 39566 35028 39618
rect 34972 39554 35028 39566
rect 34524 38782 34526 38834
rect 34578 38782 34580 38834
rect 34524 38770 34580 38782
rect 33292 38658 33348 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 38276 35140 38286
rect 35084 38182 35140 38220
rect 32620 37438 32622 37490
rect 32674 37438 32676 37490
rect 32620 37426 32676 37438
rect 33404 37940 33460 37950
rect 31836 37378 31892 37390
rect 31836 37326 31838 37378
rect 31890 37326 31892 37378
rect 30940 33294 30942 33346
rect 30994 33294 30996 33346
rect 30940 33282 30996 33294
rect 31164 36596 31220 36606
rect 29820 33236 29876 33246
rect 29484 33234 29876 33236
rect 29484 33182 29822 33234
rect 29874 33182 29876 33234
rect 29484 33180 29876 33182
rect 29484 32786 29540 33180
rect 29820 33170 29876 33180
rect 30156 33236 30212 33246
rect 30156 33142 30212 33180
rect 29484 32734 29486 32786
rect 29538 32734 29540 32786
rect 29484 32722 29540 32734
rect 29036 30884 29092 31892
rect 29372 31826 29428 31836
rect 31164 31892 31220 36540
rect 31836 35924 31892 37326
rect 33404 37380 33460 37884
rect 34300 37826 34356 37838
rect 34300 37774 34302 37826
rect 34354 37774 34356 37826
rect 34300 37490 34356 37774
rect 34300 37438 34302 37490
rect 34354 37438 34356 37490
rect 34300 37426 34356 37438
rect 34188 37380 34244 37390
rect 33404 37286 33460 37324
rect 34076 37324 34188 37380
rect 33068 37156 33124 37166
rect 32956 37154 33124 37156
rect 32956 37102 33070 37154
rect 33122 37102 33124 37154
rect 32956 37100 33124 37102
rect 32732 36484 32788 36494
rect 32732 36390 32788 36428
rect 32172 36260 32228 36270
rect 32956 36260 33012 37100
rect 33068 37090 33124 37100
rect 33516 36596 33572 36606
rect 33068 36484 33124 36494
rect 33068 36390 33124 36428
rect 33516 36482 33572 36540
rect 33516 36430 33518 36482
rect 33570 36430 33572 36482
rect 33516 36418 33572 36430
rect 32172 36258 33012 36260
rect 32172 36206 32174 36258
rect 32226 36206 33012 36258
rect 32172 36204 33012 36206
rect 32172 36194 32228 36204
rect 31836 35858 31892 35868
rect 33068 35812 33124 35822
rect 33068 35718 33124 35756
rect 33404 35812 33460 35822
rect 33404 35718 33460 35756
rect 34076 35812 34132 37324
rect 34188 37286 34244 37324
rect 35644 37266 35700 37278
rect 35644 37214 35646 37266
rect 35698 37214 35700 37266
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34076 35718 34132 35756
rect 34860 36484 34916 36494
rect 31388 35698 31444 35710
rect 31388 35646 31390 35698
rect 31442 35646 31444 35698
rect 31276 34356 31332 34366
rect 31276 34262 31332 34300
rect 31164 31826 31220 31836
rect 29036 30818 29092 30828
rect 29260 31780 29316 31790
rect 29260 30212 29316 31724
rect 29708 31780 29764 31790
rect 29708 31778 30324 31780
rect 29708 31726 29710 31778
rect 29762 31726 30324 31778
rect 29708 31724 30324 31726
rect 29708 31714 29764 31724
rect 28812 29202 28868 29214
rect 28812 29150 28814 29202
rect 28866 29150 28868 29202
rect 28812 26292 28868 29150
rect 28924 29204 28980 29214
rect 28924 29110 28980 29148
rect 29260 28754 29316 30156
rect 29260 28702 29262 28754
rect 29314 28702 29316 28754
rect 29260 28690 29316 28702
rect 29596 30210 29652 30222
rect 29596 30158 29598 30210
rect 29650 30158 29652 30210
rect 29596 27972 29652 30158
rect 29708 29540 29764 29550
rect 29708 29446 29764 29484
rect 29708 28644 29764 28654
rect 29708 28550 29764 28588
rect 29932 28642 29988 28654
rect 29932 28590 29934 28642
rect 29986 28590 29988 28642
rect 29932 28532 29988 28590
rect 29932 28466 29988 28476
rect 29596 27906 29652 27916
rect 30156 28420 30212 28430
rect 29260 27074 29316 27086
rect 29260 27022 29262 27074
rect 29314 27022 29316 27074
rect 28812 26236 28980 26292
rect 28700 24210 28756 24220
rect 28812 26066 28868 26078
rect 28812 26014 28814 26066
rect 28866 26014 28868 26066
rect 28812 23828 28868 26014
rect 28924 24612 28980 26236
rect 29148 26290 29204 26302
rect 29148 26238 29150 26290
rect 29202 26238 29204 26290
rect 29148 25284 29204 26238
rect 29260 25508 29316 27022
rect 29708 27074 29764 27086
rect 29708 27022 29710 27074
rect 29762 27022 29764 27074
rect 29372 26740 29428 26750
rect 29428 26684 29540 26740
rect 29372 26674 29428 26684
rect 29260 25442 29316 25452
rect 29372 26516 29428 26526
rect 29148 25218 29204 25228
rect 29372 25282 29428 26460
rect 29372 25230 29374 25282
rect 29426 25230 29428 25282
rect 29372 25218 29428 25230
rect 29484 25732 29540 26684
rect 29484 25618 29540 25676
rect 29484 25566 29486 25618
rect 29538 25566 29540 25618
rect 28924 24546 28980 24556
rect 29148 24052 29204 24062
rect 29148 23958 29204 23996
rect 29484 24050 29540 25566
rect 29484 23998 29486 24050
rect 29538 23998 29540 24050
rect 29484 23986 29540 23998
rect 29596 26290 29652 26302
rect 29596 26238 29598 26290
rect 29650 26238 29652 26290
rect 28812 23772 29428 23828
rect 28700 23716 28756 23726
rect 28700 23714 29316 23716
rect 28700 23662 28702 23714
rect 28754 23662 29316 23714
rect 28700 23660 29316 23662
rect 28700 23650 28756 23660
rect 28476 23548 28644 23604
rect 28588 22484 28644 23548
rect 29148 23156 29204 23166
rect 29148 23062 29204 23100
rect 28812 22930 28868 22942
rect 28812 22878 28814 22930
rect 28866 22878 28868 22930
rect 28588 22428 28756 22484
rect 28588 22260 28644 22270
rect 28588 22166 28644 22204
rect 28476 21586 28532 21598
rect 28476 21534 28478 21586
rect 28530 21534 28532 21586
rect 28476 18564 28532 21534
rect 28476 18498 28532 18508
rect 28364 17502 28366 17554
rect 28418 17502 28420 17554
rect 28364 17490 28420 17502
rect 28700 16994 28756 22428
rect 28812 20356 28868 22878
rect 29148 22820 29204 22830
rect 28812 20290 28868 20300
rect 28924 22764 29148 22820
rect 28924 18562 28980 22764
rect 29148 22754 29204 22764
rect 29148 22596 29204 22606
rect 29148 22370 29204 22540
rect 29148 22318 29150 22370
rect 29202 22318 29204 22370
rect 29148 22306 29204 22318
rect 28924 18510 28926 18562
rect 28978 18510 28980 18562
rect 28924 18498 28980 18510
rect 28700 16942 28702 16994
rect 28754 16942 28756 16994
rect 28700 16930 28756 16942
rect 29260 16996 29316 23660
rect 29372 18564 29428 23772
rect 29596 23604 29652 26238
rect 29708 25620 29764 27022
rect 29708 25554 29764 25564
rect 30044 25284 30100 25294
rect 30044 24834 30100 25228
rect 30044 24782 30046 24834
rect 30098 24782 30100 24834
rect 30044 24770 30100 24782
rect 30044 24612 30100 24622
rect 29596 23538 29652 23548
rect 29708 24276 29764 24286
rect 29596 23154 29652 23166
rect 29596 23102 29598 23154
rect 29650 23102 29652 23154
rect 29484 21588 29540 21598
rect 29484 19572 29540 21532
rect 29596 20244 29652 23102
rect 29596 20178 29652 20188
rect 29708 20130 29764 24220
rect 29932 23714 29988 23726
rect 29932 23662 29934 23714
rect 29986 23662 29988 23714
rect 29932 23156 29988 23662
rect 29932 23090 29988 23100
rect 29708 20078 29710 20130
rect 29762 20078 29764 20130
rect 29708 20066 29764 20078
rect 29484 19516 29652 19572
rect 29484 18564 29540 18574
rect 29372 18562 29540 18564
rect 29372 18510 29486 18562
rect 29538 18510 29540 18562
rect 29372 18508 29540 18510
rect 29484 18498 29540 18508
rect 29372 16996 29428 17006
rect 29260 16994 29428 16996
rect 29260 16942 29374 16994
rect 29426 16942 29428 16994
rect 29260 16940 29428 16942
rect 29372 16930 29428 16940
rect 29596 15426 29652 19516
rect 30044 19122 30100 24556
rect 30156 22820 30212 28364
rect 30156 22754 30212 22764
rect 30156 22260 30212 22270
rect 30156 22146 30212 22204
rect 30156 22094 30158 22146
rect 30210 22094 30212 22146
rect 30156 22082 30212 22094
rect 30268 19908 30324 31724
rect 30492 29540 30548 29550
rect 30492 28754 30548 29484
rect 31164 29428 31220 29438
rect 30492 28702 30494 28754
rect 30546 28702 30548 28754
rect 30492 28690 30548 28702
rect 30716 28756 30772 28766
rect 30716 28662 30772 28700
rect 30940 28420 30996 28430
rect 30940 28326 30996 28364
rect 30604 27860 30660 27870
rect 30604 27858 31108 27860
rect 30604 27806 30606 27858
rect 30658 27806 31108 27858
rect 30604 27804 31108 27806
rect 30604 27794 30660 27804
rect 30380 25732 30436 25742
rect 30436 25676 30548 25732
rect 30380 25666 30436 25676
rect 30492 25618 30548 25676
rect 30492 25566 30494 25618
rect 30546 25566 30548 25618
rect 30492 25554 30548 25566
rect 30828 25620 30884 25630
rect 30380 25396 30436 25406
rect 30380 25282 30436 25340
rect 30380 25230 30382 25282
rect 30434 25230 30436 25282
rect 30380 25218 30436 25230
rect 30604 23828 30660 23838
rect 30492 23826 30660 23828
rect 30492 23774 30606 23826
rect 30658 23774 30660 23826
rect 30492 23772 30660 23774
rect 30492 23044 30548 23772
rect 30604 23762 30660 23772
rect 30716 23714 30772 23726
rect 30716 23662 30718 23714
rect 30770 23662 30772 23714
rect 30492 22260 30548 22988
rect 30492 22194 30548 22204
rect 30604 23604 30660 23614
rect 30604 21588 30660 23548
rect 30716 21810 30772 23662
rect 30716 21758 30718 21810
rect 30770 21758 30772 21810
rect 30716 21746 30772 21758
rect 30604 21532 30772 21588
rect 30604 19908 30660 19918
rect 30268 19906 30660 19908
rect 30268 19854 30606 19906
rect 30658 19854 30660 19906
rect 30268 19852 30660 19854
rect 30604 19842 30660 19852
rect 30044 19070 30046 19122
rect 30098 19070 30100 19122
rect 30044 19058 30100 19070
rect 29596 15374 29598 15426
rect 29650 15374 29652 15426
rect 29596 15362 29652 15374
rect 30156 18564 30212 18574
rect 28252 15150 28254 15202
rect 28306 15150 28308 15202
rect 28252 15138 28308 15150
rect 27356 14644 27412 14654
rect 27020 14642 27412 14644
rect 27020 14590 27358 14642
rect 27410 14590 27412 14642
rect 27020 14588 27412 14590
rect 27356 14578 27412 14588
rect 30156 14642 30212 18508
rect 30716 16770 30772 21532
rect 30828 18338 30884 25564
rect 30940 25284 30996 25294
rect 30940 25190 30996 25228
rect 30940 24724 30996 24734
rect 30940 24630 30996 24668
rect 31052 19346 31108 27804
rect 31164 27858 31220 29372
rect 31164 27806 31166 27858
rect 31218 27806 31220 27858
rect 31164 27794 31220 27806
rect 31388 27188 31444 35646
rect 31948 35698 32004 35710
rect 31948 35646 31950 35698
rect 32002 35646 32004 35698
rect 31836 35252 31892 35262
rect 31836 34354 31892 35196
rect 31836 34302 31838 34354
rect 31890 34302 31892 34354
rect 31836 34290 31892 34302
rect 31948 33684 32004 35646
rect 32396 35700 32452 35710
rect 32060 34244 32116 34254
rect 32060 34150 32116 34188
rect 32396 34242 32452 35644
rect 34860 35698 34916 36428
rect 35644 36484 35700 37214
rect 36316 37266 36372 42028
rect 36652 42082 36708 42094
rect 36652 42030 36654 42082
rect 36706 42030 36708 42082
rect 36652 41300 36708 42030
rect 36652 41234 36708 41244
rect 36988 41748 37044 41758
rect 36988 41298 37044 41692
rect 36988 41246 36990 41298
rect 37042 41246 37044 41298
rect 36988 41234 37044 41246
rect 36428 41074 36484 41086
rect 36428 41022 36430 41074
rect 36482 41022 36484 41074
rect 36428 40626 36484 41022
rect 37100 40964 37156 40974
rect 37100 40870 37156 40908
rect 36428 40574 36430 40626
rect 36482 40574 36484 40626
rect 36428 40562 36484 40574
rect 37212 40628 37268 40638
rect 37212 40534 37268 40572
rect 37436 39394 37492 39406
rect 37436 39342 37438 39394
rect 37490 39342 37492 39394
rect 36316 37214 36318 37266
rect 36370 37214 36372 37266
rect 36316 37202 36372 37214
rect 36876 39058 36932 39070
rect 36876 39006 36878 39058
rect 36930 39006 36932 39058
rect 36876 37044 36932 39006
rect 37436 38948 37492 39342
rect 37548 39060 37604 39070
rect 37660 39060 37716 43932
rect 37772 39842 37828 44828
rect 39116 43708 39172 48972
rect 39452 46898 39508 52220
rect 40012 50706 40068 50718
rect 40012 50654 40014 50706
rect 40066 50654 40068 50706
rect 40012 48692 40068 50654
rect 39452 46846 39454 46898
rect 39506 46846 39508 46898
rect 39452 46834 39508 46846
rect 39676 48636 40068 48692
rect 39676 43708 39732 48636
rect 39900 48466 39956 48478
rect 39900 48414 39902 48466
rect 39954 48414 39956 48466
rect 39900 46788 39956 48414
rect 40348 47348 40404 53788
rect 41356 53778 41412 53788
rect 41244 53060 41300 53070
rect 40572 53058 41300 53060
rect 40572 53006 41246 53058
rect 41298 53006 41300 53058
rect 40572 53004 41300 53006
rect 40460 50484 40516 50494
rect 40460 48466 40516 50428
rect 40460 48414 40462 48466
rect 40514 48414 40516 48466
rect 40460 48402 40516 48414
rect 40460 47572 40516 47582
rect 40460 47478 40516 47516
rect 40348 47292 40516 47348
rect 40012 46788 40068 46798
rect 39900 46786 40068 46788
rect 39900 46734 40014 46786
rect 40066 46734 40068 46786
rect 39900 46732 40068 46734
rect 40012 46722 40068 46732
rect 40348 46788 40404 46798
rect 40348 46694 40404 46732
rect 40460 45890 40516 47292
rect 40460 45838 40462 45890
rect 40514 45838 40516 45890
rect 40460 45826 40516 45838
rect 39900 45330 39956 45342
rect 39900 45278 39902 45330
rect 39954 45278 39956 45330
rect 39900 45220 39956 45278
rect 40460 45332 40516 45342
rect 40572 45332 40628 53004
rect 41244 52994 41300 53004
rect 40796 52274 40852 52286
rect 40796 52222 40798 52274
rect 40850 52222 40852 52274
rect 40460 45330 40628 45332
rect 40460 45278 40462 45330
rect 40514 45278 40628 45330
rect 40460 45276 40628 45278
rect 40684 52052 40740 52062
rect 40460 45266 40516 45276
rect 40684 45220 40740 51996
rect 40796 50596 40852 52222
rect 40796 50530 40852 50540
rect 41356 50148 41412 50158
rect 41244 50092 41356 50148
rect 41132 48804 41188 48814
rect 41132 48710 41188 48748
rect 41244 48580 41300 50092
rect 41356 50082 41412 50092
rect 41132 48524 41300 48580
rect 41356 48916 41412 48926
rect 40908 48132 40964 48142
rect 40908 48038 40964 48076
rect 40796 47572 40852 47582
rect 40796 46674 40852 47516
rect 40796 46622 40798 46674
rect 40850 46622 40852 46674
rect 40796 45892 40852 46622
rect 41020 46004 41076 46014
rect 40908 45892 40964 45902
rect 40796 45890 40964 45892
rect 40796 45838 40910 45890
rect 40962 45838 40964 45890
rect 40796 45836 40964 45838
rect 40908 45826 40964 45836
rect 41020 45330 41076 45948
rect 41020 45278 41022 45330
rect 41074 45278 41076 45330
rect 41020 45266 41076 45278
rect 39900 45154 39956 45164
rect 40572 45164 40740 45220
rect 40572 45108 40628 45164
rect 40460 45052 40628 45108
rect 38892 43652 39172 43708
rect 39452 43652 39732 43708
rect 39900 44098 39956 44110
rect 39900 44046 39902 44098
rect 39954 44046 39956 44098
rect 38892 41970 38948 43652
rect 38892 41918 38894 41970
rect 38946 41918 38948 41970
rect 38892 41906 38948 41918
rect 39004 43426 39060 43438
rect 39004 43374 39006 43426
rect 39058 43374 39060 43426
rect 39004 42756 39060 43374
rect 39004 41972 39060 42700
rect 38220 41300 38276 41310
rect 38220 41206 38276 41244
rect 39004 41186 39060 41916
rect 39004 41134 39006 41186
rect 39058 41134 39060 41186
rect 39004 41122 39060 41134
rect 39452 41186 39508 43652
rect 39564 41972 39620 41982
rect 39564 41878 39620 41916
rect 39900 41858 39956 44046
rect 40460 42980 40516 45052
rect 41132 44884 41188 48524
rect 41244 48356 41300 48366
rect 41356 48356 41412 48860
rect 41244 48354 41412 48356
rect 41244 48302 41246 48354
rect 41298 48302 41412 48354
rect 41244 48300 41412 48302
rect 41244 46788 41300 48300
rect 41244 46722 41300 46732
rect 41468 46674 41524 54348
rect 42700 54404 42756 54414
rect 42700 54310 42756 54348
rect 43036 53844 43092 53854
rect 42364 53618 42420 53630
rect 42364 53566 42366 53618
rect 42418 53566 42420 53618
rect 42364 52276 42420 53566
rect 42588 52836 42644 52846
rect 42588 52834 42756 52836
rect 42588 52782 42590 52834
rect 42642 52782 42756 52834
rect 42588 52780 42756 52782
rect 42588 52770 42644 52780
rect 42364 52210 42420 52220
rect 41692 52164 41748 52174
rect 41468 46622 41470 46674
rect 41522 46622 41524 46674
rect 41468 46610 41524 46622
rect 41580 49252 41636 49262
rect 41580 46452 41636 49196
rect 41692 49250 41748 52108
rect 41804 52052 41860 52062
rect 41804 51958 41860 51996
rect 41692 49198 41694 49250
rect 41746 49198 41748 49250
rect 41692 49186 41748 49198
rect 41916 51266 41972 51278
rect 41916 51214 41918 51266
rect 41970 51214 41972 51266
rect 41916 49028 41972 51214
rect 42588 50706 42644 50718
rect 42588 50654 42590 50706
rect 42642 50654 42644 50706
rect 42476 50372 42532 50382
rect 42252 49812 42308 49822
rect 41916 48962 41972 48972
rect 42028 49810 42308 49812
rect 42028 49758 42254 49810
rect 42306 49758 42308 49810
rect 42028 49756 42308 49758
rect 41916 48244 41972 48254
rect 42028 48244 42084 49756
rect 42252 49746 42308 49756
rect 42252 48916 42308 48926
rect 42252 48822 42308 48860
rect 41916 48242 42084 48244
rect 41916 48190 41918 48242
rect 41970 48190 42084 48242
rect 41916 48188 42084 48190
rect 42140 48802 42196 48814
rect 42140 48750 42142 48802
rect 42194 48750 42196 48802
rect 41916 47572 41972 48188
rect 41916 47506 41972 47516
rect 42028 47236 42084 47246
rect 42140 47236 42196 48750
rect 42252 48244 42308 48254
rect 42476 48244 42532 50316
rect 42252 48242 42532 48244
rect 42252 48190 42254 48242
rect 42306 48190 42532 48242
rect 42252 48188 42532 48190
rect 42252 48178 42308 48188
rect 42476 48020 42532 48030
rect 42364 47964 42476 48020
rect 42084 47180 42196 47236
rect 42252 47458 42308 47470
rect 42252 47406 42254 47458
rect 42306 47406 42308 47458
rect 42252 47236 42308 47406
rect 42028 47170 42084 47180
rect 42252 47170 42308 47180
rect 40572 44828 41188 44884
rect 41244 46396 41636 46452
rect 40572 44546 40628 44828
rect 40572 44494 40574 44546
rect 40626 44494 40628 44546
rect 40572 44482 40628 44494
rect 40908 44100 40964 44110
rect 40908 44098 41076 44100
rect 40908 44046 40910 44098
rect 40962 44046 41076 44098
rect 40908 44044 41076 44046
rect 40908 44034 40964 44044
rect 40908 43876 40964 43886
rect 40908 43538 40964 43820
rect 40908 43486 40910 43538
rect 40962 43486 40964 43538
rect 40572 42980 40628 42990
rect 40460 42978 40628 42980
rect 40460 42926 40574 42978
rect 40626 42926 40628 42978
rect 40460 42924 40628 42926
rect 40572 42914 40628 42924
rect 40908 42754 40964 43486
rect 41020 43540 41076 44044
rect 41076 43484 41188 43540
rect 41020 43474 41076 43484
rect 40908 42702 40910 42754
rect 40962 42702 40964 42754
rect 40908 42690 40964 42702
rect 39900 41806 39902 41858
rect 39954 41806 39956 41858
rect 39900 41794 39956 41806
rect 40012 42530 40068 42542
rect 40012 42478 40014 42530
rect 40066 42478 40068 42530
rect 40012 41300 40068 42478
rect 40796 41972 40852 41982
rect 40796 41878 40852 41916
rect 40012 41234 40068 41244
rect 40124 41858 40180 41870
rect 40124 41806 40126 41858
rect 40178 41806 40180 41858
rect 39452 41134 39454 41186
rect 39506 41134 39508 41186
rect 39452 41122 39508 41134
rect 38556 41076 38612 41086
rect 38556 40982 38612 41020
rect 40124 41076 40180 41806
rect 40124 41010 40180 41020
rect 39452 40514 39508 40526
rect 39452 40462 39454 40514
rect 39506 40462 39508 40514
rect 38556 40404 38612 40414
rect 38444 40292 38500 40302
rect 38444 40198 38500 40236
rect 37772 39790 37774 39842
rect 37826 39790 37828 39842
rect 37772 39778 37828 39790
rect 38556 39506 38612 40348
rect 38556 39454 38558 39506
rect 38610 39454 38612 39506
rect 38556 39442 38612 39454
rect 37548 39058 37716 39060
rect 37548 39006 37550 39058
rect 37602 39006 37716 39058
rect 37548 39004 37716 39006
rect 37548 38994 37604 39004
rect 37436 38882 37492 38892
rect 37996 38610 38052 38622
rect 37996 38558 37998 38610
rect 38050 38558 38052 38610
rect 37436 38164 37492 38174
rect 37436 37380 37492 38108
rect 36876 36988 37156 37044
rect 36540 36708 36596 36718
rect 36540 36614 36596 36652
rect 35644 36418 35700 36428
rect 35980 36372 36036 36382
rect 35980 36258 36036 36316
rect 36988 36372 37044 36382
rect 36988 36278 37044 36316
rect 35980 36206 35982 36258
rect 36034 36206 36036 36258
rect 35980 36194 36036 36206
rect 34860 35646 34862 35698
rect 34914 35646 34916 35698
rect 34860 35634 34916 35646
rect 35532 36036 35588 36046
rect 35532 35698 35588 35980
rect 35532 35646 35534 35698
rect 35586 35646 35588 35698
rect 35532 35634 35588 35646
rect 32620 35588 32676 35598
rect 33740 35588 33796 35598
rect 32396 34190 32398 34242
rect 32450 34190 32452 34242
rect 32396 34178 32452 34190
rect 32508 35586 32676 35588
rect 32508 35534 32622 35586
rect 32674 35534 32676 35586
rect 32508 35532 32676 35534
rect 31836 33628 32004 33684
rect 31836 33348 31892 33628
rect 31836 33282 31892 33292
rect 32508 33460 32564 35532
rect 32620 35522 32676 35532
rect 33628 35586 33796 35588
rect 33628 35534 33742 35586
rect 33794 35534 33796 35586
rect 33628 35532 33796 35534
rect 33628 34132 33684 35532
rect 33740 35522 33796 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 37100 35026 37156 36988
rect 37100 34974 37102 35026
rect 37154 34974 37156 35026
rect 37100 34962 37156 34974
rect 37324 36596 37380 36606
rect 37436 36596 37492 37324
rect 37324 36594 37492 36596
rect 37324 36542 37326 36594
rect 37378 36542 37492 36594
rect 37324 36540 37492 36542
rect 37660 38162 37716 38174
rect 37660 38110 37662 38162
rect 37714 38110 37716 38162
rect 37324 35026 37380 36540
rect 37660 35924 37716 38110
rect 37996 38164 38052 38558
rect 38108 38164 38164 38174
rect 38052 38162 38164 38164
rect 38052 38110 38110 38162
rect 38162 38110 38164 38162
rect 38052 38108 38164 38110
rect 37996 38070 38052 38108
rect 38108 38098 38164 38108
rect 39228 38050 39284 38062
rect 39228 37998 39230 38050
rect 39282 37998 39284 38050
rect 38444 37938 38500 37950
rect 38444 37886 38446 37938
rect 38498 37886 38500 37938
rect 38444 37492 38500 37886
rect 38556 37492 38612 37502
rect 38444 37490 38612 37492
rect 38444 37438 38558 37490
rect 38610 37438 38612 37490
rect 38444 37436 38612 37438
rect 38556 37426 38612 37436
rect 38556 37268 38612 37278
rect 38444 37212 38556 37268
rect 39228 37268 39284 37998
rect 39452 37492 39508 40462
rect 40908 39620 40964 39630
rect 40908 39526 40964 39564
rect 40908 39172 40964 39182
rect 40236 38948 40292 38958
rect 40236 38834 40292 38892
rect 40908 38836 40964 39116
rect 41132 38948 41188 43484
rect 41244 42754 41300 46396
rect 41804 46004 41860 46014
rect 41804 45890 41860 45948
rect 41804 45838 41806 45890
rect 41858 45838 41860 45890
rect 41804 45826 41860 45838
rect 42364 45330 42420 47964
rect 42476 47954 42532 47964
rect 42364 45278 42366 45330
rect 42418 45278 42420 45330
rect 42364 45266 42420 45278
rect 41468 45220 41524 45230
rect 41468 45126 41524 45164
rect 41692 45106 41748 45118
rect 41692 45054 41694 45106
rect 41746 45054 41748 45106
rect 41468 44996 41524 45006
rect 41468 43538 41524 44940
rect 41692 44212 41748 45054
rect 41692 44146 41748 44156
rect 41804 44434 41860 44446
rect 41804 44382 41806 44434
rect 41858 44382 41860 44434
rect 41468 43486 41470 43538
rect 41522 43486 41524 43538
rect 41468 43474 41524 43486
rect 41244 42702 41246 42754
rect 41298 42702 41300 42754
rect 41244 42690 41300 42702
rect 41468 42868 41524 42878
rect 41468 41970 41524 42812
rect 41804 42084 41860 44382
rect 42588 42868 42644 50654
rect 42700 44996 42756 52780
rect 42924 49812 42980 49822
rect 43036 49812 43092 53788
rect 43708 52164 43764 54574
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 45836 53844 45892 53854
rect 45836 53750 45892 53788
rect 43708 52098 43764 52108
rect 44492 53620 44548 53630
rect 42924 49810 43092 49812
rect 42924 49758 42926 49810
rect 42978 49758 43092 49810
rect 42924 49756 43092 49758
rect 43148 51490 43204 51502
rect 43148 51438 43150 51490
rect 43202 51438 43204 51490
rect 42924 49746 42980 49756
rect 42924 48916 42980 48926
rect 42924 48822 42980 48860
rect 42812 48804 42868 48814
rect 42812 48710 42868 48748
rect 43148 48020 43204 51438
rect 43932 50482 43988 50494
rect 43932 50430 43934 50482
rect 43986 50430 43988 50482
rect 43372 49028 43428 49038
rect 43372 49026 43540 49028
rect 43372 48974 43374 49026
rect 43426 48974 43540 49026
rect 43372 48972 43540 48974
rect 43372 48962 43428 48972
rect 43148 47954 43204 47964
rect 43484 48916 43540 48972
rect 42924 47236 42980 47246
rect 42924 45668 42980 47180
rect 43484 46004 43540 48860
rect 43596 48914 43652 48926
rect 43596 48862 43598 48914
rect 43650 48862 43652 48914
rect 43596 47068 43652 48862
rect 43596 47012 43764 47068
rect 43708 46898 43764 47012
rect 43708 46846 43710 46898
rect 43762 46846 43764 46898
rect 43708 46834 43764 46846
rect 43596 46004 43652 46014
rect 43484 46002 43652 46004
rect 43484 45950 43598 46002
rect 43650 45950 43652 46002
rect 43484 45948 43652 45950
rect 42924 45602 42980 45612
rect 43148 45220 43204 45230
rect 43148 45126 43204 45164
rect 42700 44930 42756 44940
rect 43596 44996 43652 45948
rect 43596 44930 43652 44940
rect 42812 44210 42868 44222
rect 42812 44158 42814 44210
rect 42866 44158 42868 44210
rect 42812 43988 42868 44158
rect 43596 44212 43652 44222
rect 43596 44118 43652 44156
rect 42812 43922 42868 43932
rect 43708 44098 43764 44110
rect 43708 44046 43710 44098
rect 43762 44046 43764 44098
rect 43708 43762 43764 44046
rect 43708 43710 43710 43762
rect 43762 43710 43764 43762
rect 43708 43698 43764 43710
rect 43932 43708 43988 50430
rect 44268 48244 44324 48254
rect 44268 47570 44324 48188
rect 44268 47518 44270 47570
rect 44322 47518 44324 47570
rect 44268 47506 44324 47518
rect 44380 47236 44436 47246
rect 44380 46676 44436 47180
rect 44492 46898 44548 53564
rect 47068 53620 47124 53630
rect 47068 53526 47124 53564
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 44492 46846 44494 46898
rect 44546 46846 44548 46898
rect 44492 46834 44548 46846
rect 44604 53060 44660 53070
rect 44604 46898 44660 53004
rect 45948 53060 46004 53070
rect 45948 52966 46004 53004
rect 51100 53058 51156 53070
rect 51100 53006 51102 53058
rect 51154 53006 51156 53058
rect 44940 52834 44996 52846
rect 50092 52836 50148 52846
rect 44940 52782 44942 52834
rect 44994 52782 44996 52834
rect 44716 51266 44772 51278
rect 44716 51214 44718 51266
rect 44770 51214 44772 51266
rect 44716 49252 44772 51214
rect 44940 50372 44996 52782
rect 49196 52834 50148 52836
rect 49196 52782 50094 52834
rect 50146 52782 50148 52834
rect 49196 52780 50148 52782
rect 46060 52276 46116 52286
rect 48636 52276 48692 52286
rect 46060 52274 46340 52276
rect 46060 52222 46062 52274
rect 46114 52222 46340 52274
rect 46060 52220 46340 52222
rect 46060 52210 46116 52220
rect 44940 50306 44996 50316
rect 45724 51490 45780 51502
rect 45724 51438 45726 51490
rect 45778 51438 45780 51490
rect 45724 50148 45780 51438
rect 45948 51492 46004 51502
rect 45836 50708 45892 50718
rect 45836 50614 45892 50652
rect 45724 50082 45780 50092
rect 45388 50034 45444 50046
rect 45388 49982 45390 50034
rect 45442 49982 45444 50034
rect 45388 49924 45444 49982
rect 45948 50034 46004 51436
rect 45948 49982 45950 50034
rect 46002 49982 46004 50034
rect 45948 49970 46004 49982
rect 46060 50708 46116 50718
rect 45388 49858 45444 49868
rect 45612 49812 45668 49822
rect 45500 49756 45612 49812
rect 44716 49186 44772 49196
rect 44828 49700 44884 49710
rect 44828 48466 44884 49644
rect 45388 49588 45444 49598
rect 44828 48414 44830 48466
rect 44882 48414 44884 48466
rect 44828 48402 44884 48414
rect 44940 49026 44996 49038
rect 44940 48974 44942 49026
rect 44994 48974 44996 49026
rect 44604 46846 44606 46898
rect 44658 46846 44660 46898
rect 44604 46834 44660 46846
rect 44828 48244 44884 48254
rect 44716 46788 44772 46798
rect 44380 46620 44548 46676
rect 43932 43652 44436 43708
rect 44380 42978 44436 43652
rect 44492 43650 44548 46620
rect 44716 43708 44772 46732
rect 44828 46004 44884 48188
rect 44940 47458 44996 48974
rect 45388 48466 45444 49532
rect 45388 48414 45390 48466
rect 45442 48414 45444 48466
rect 45388 48402 45444 48414
rect 44940 47406 44942 47458
rect 44994 47406 44996 47458
rect 44940 47124 44996 47406
rect 45388 47460 45444 47470
rect 45500 47460 45556 49756
rect 45612 49746 45668 49756
rect 45612 49140 45668 49150
rect 45612 49026 45668 49084
rect 45612 48974 45614 49026
rect 45666 48974 45668 49026
rect 45612 48962 45668 48974
rect 45612 48244 45668 48254
rect 45612 48150 45668 48188
rect 45388 47458 45556 47460
rect 45388 47406 45390 47458
rect 45442 47406 45556 47458
rect 45388 47404 45556 47406
rect 45388 47394 45444 47404
rect 44940 47058 44996 47068
rect 45388 46786 45444 46798
rect 45388 46734 45390 46786
rect 45442 46734 45444 46786
rect 44940 46004 44996 46014
rect 44884 46002 44996 46004
rect 44884 45950 44942 46002
rect 44994 45950 44996 46002
rect 44884 45948 44996 45950
rect 44828 45910 44884 45948
rect 44492 43598 44494 43650
rect 44546 43598 44548 43650
rect 44492 43586 44548 43598
rect 44604 43652 44772 43708
rect 44380 42926 44382 42978
rect 44434 42926 44436 42978
rect 44380 42914 44436 42926
rect 42588 42802 42644 42812
rect 41804 42018 41860 42028
rect 43596 42530 43652 42542
rect 43596 42478 43598 42530
rect 43650 42478 43652 42530
rect 41468 41918 41470 41970
rect 41522 41918 41524 41970
rect 41468 41906 41524 41918
rect 43596 41412 43652 42478
rect 43932 42194 43988 42206
rect 43932 42142 43934 42194
rect 43986 42142 43988 42194
rect 43596 41356 43876 41412
rect 43372 41300 43428 41310
rect 43372 41206 43428 41244
rect 42476 41188 42532 41198
rect 42476 41094 42532 41132
rect 42700 41074 42756 41086
rect 42700 41022 42702 41074
rect 42754 41022 42756 41074
rect 41692 40962 41748 40974
rect 41692 40910 41694 40962
rect 41746 40910 41748 40962
rect 41244 39618 41300 39630
rect 41244 39566 41246 39618
rect 41298 39566 41300 39618
rect 41244 39172 41300 39566
rect 41692 39620 41748 40910
rect 42700 40404 42756 41022
rect 43036 41076 43092 41086
rect 43708 41076 43764 41086
rect 43036 41074 43204 41076
rect 43036 41022 43038 41074
rect 43090 41022 43204 41074
rect 43036 41020 43204 41022
rect 43036 41010 43092 41020
rect 43148 40964 43204 41020
rect 42700 40338 42756 40348
rect 42812 40516 42868 40526
rect 41692 39554 41748 39564
rect 41916 40290 41972 40302
rect 41916 40238 41918 40290
rect 41970 40238 41972 40290
rect 41244 39106 41300 39116
rect 41804 39394 41860 39406
rect 41804 39342 41806 39394
rect 41858 39342 41860 39394
rect 41804 39172 41860 39342
rect 41804 39106 41860 39116
rect 41580 39060 41636 39070
rect 41132 38892 41412 38948
rect 40236 38782 40238 38834
rect 40290 38782 40292 38834
rect 40236 38770 40292 38782
rect 40796 38834 40964 38836
rect 40796 38782 40910 38834
rect 40962 38782 40964 38834
rect 40796 38780 40964 38782
rect 40796 38668 40852 38780
rect 40908 38770 40964 38780
rect 40796 38612 41076 38668
rect 39676 38500 39732 38510
rect 39676 38050 39732 38444
rect 39676 37998 39678 38050
rect 39730 37998 39732 38050
rect 39676 37986 39732 37998
rect 39452 37426 39508 37436
rect 39228 37212 39508 37268
rect 37772 36484 37828 36494
rect 37996 36484 38052 36494
rect 37828 36482 38052 36484
rect 37828 36430 37998 36482
rect 38050 36430 38052 36482
rect 37828 36428 38052 36430
rect 37772 36390 37828 36428
rect 37996 36418 38052 36428
rect 37772 35924 37828 35934
rect 37660 35922 37828 35924
rect 37660 35870 37774 35922
rect 37826 35870 37828 35922
rect 37660 35868 37828 35870
rect 38444 35924 38500 37212
rect 38556 37202 38612 37212
rect 39452 37156 39508 37212
rect 39676 37156 39732 37166
rect 39452 37154 39732 37156
rect 39452 37102 39678 37154
rect 39730 37102 39732 37154
rect 39452 37100 39732 37102
rect 39340 37042 39396 37054
rect 39340 36990 39342 37042
rect 39394 36990 39396 37042
rect 38668 36482 38724 36494
rect 38668 36430 38670 36482
rect 38722 36430 38724 36482
rect 38556 35924 38612 35934
rect 38444 35922 38612 35924
rect 38444 35870 38558 35922
rect 38610 35870 38612 35922
rect 38444 35868 38612 35870
rect 37772 35858 37828 35868
rect 38556 35858 38612 35868
rect 37324 34974 37326 35026
rect 37378 34974 37380 35026
rect 37324 34962 37380 34974
rect 38556 35028 38612 35038
rect 35196 34916 35252 34926
rect 35196 34802 35252 34860
rect 37884 34916 37940 34926
rect 37884 34822 37940 34860
rect 35196 34750 35198 34802
rect 35250 34750 35252 34802
rect 35196 34738 35252 34750
rect 36540 34690 36596 34702
rect 36540 34638 36542 34690
rect 36594 34638 36596 34690
rect 36092 34468 36148 34478
rect 33740 34244 33796 34254
rect 33740 34242 34356 34244
rect 33740 34190 33742 34242
rect 33794 34190 34356 34242
rect 33740 34188 34356 34190
rect 33740 34178 33796 34188
rect 33516 34076 33684 34132
rect 32956 33908 33012 33918
rect 32956 33814 33012 33852
rect 31836 32562 31892 32574
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31500 28532 31556 28542
rect 31500 27970 31556 28476
rect 31724 28420 31780 28430
rect 31724 28326 31780 28364
rect 31836 28084 31892 32510
rect 32396 32564 32452 32574
rect 32508 32564 32564 33404
rect 33516 33122 33572 34076
rect 34300 33458 34356 34188
rect 36092 34130 36148 34412
rect 36540 34468 36596 34638
rect 36540 34402 36596 34412
rect 36092 34078 36094 34130
rect 36146 34078 36148 34130
rect 36092 34066 36148 34078
rect 36428 34130 36484 34142
rect 36428 34078 36430 34130
rect 36482 34078 36484 34130
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34300 33406 34302 33458
rect 34354 33406 34356 33458
rect 34300 33394 34356 33406
rect 35084 33460 35140 33470
rect 35084 33366 35140 33404
rect 35644 33460 35700 33470
rect 35644 33366 35700 33404
rect 36428 33460 36484 34078
rect 36428 33394 36484 33404
rect 36764 34130 36820 34142
rect 36764 34078 36766 34130
rect 36818 34078 36820 34130
rect 34524 33346 34580 33358
rect 34524 33294 34526 33346
rect 34578 33294 34580 33346
rect 34524 33236 34580 33294
rect 36092 33346 36148 33358
rect 36092 33294 36094 33346
rect 36146 33294 36148 33346
rect 34524 33170 34580 33180
rect 35868 33234 35924 33246
rect 35868 33182 35870 33234
rect 35922 33182 35924 33234
rect 33516 33070 33518 33122
rect 33570 33070 33572 33122
rect 33516 33058 33572 33070
rect 34076 33122 34132 33134
rect 34076 33070 34078 33122
rect 34130 33070 34132 33122
rect 32396 32562 32564 32564
rect 32396 32510 32398 32562
rect 32450 32510 32564 32562
rect 32396 32508 32564 32510
rect 33740 32674 33796 32686
rect 33740 32622 33742 32674
rect 33794 32622 33796 32674
rect 32396 31948 32452 32508
rect 32172 31892 32452 31948
rect 32956 32338 33012 32350
rect 32956 32286 32958 32338
rect 33010 32286 33012 32338
rect 32956 31948 33012 32286
rect 32956 31892 33124 31948
rect 32172 31780 32228 31892
rect 32060 31554 32116 31566
rect 32060 31502 32062 31554
rect 32114 31502 32116 31554
rect 32060 29652 32116 31502
rect 32172 30884 32228 31724
rect 32956 31778 33012 31790
rect 32956 31726 32958 31778
rect 33010 31726 33012 31778
rect 32732 31556 32788 31566
rect 32172 30790 32228 30828
rect 32284 31554 32788 31556
rect 32284 31502 32734 31554
rect 32786 31502 32788 31554
rect 32284 31500 32788 31502
rect 32172 29988 32228 29998
rect 32172 29894 32228 29932
rect 32060 29586 32116 29596
rect 32060 29428 32116 29438
rect 32060 29334 32116 29372
rect 31836 28018 31892 28028
rect 31500 27918 31502 27970
rect 31554 27918 31556 27970
rect 31500 27906 31556 27918
rect 31388 27122 31444 27132
rect 31836 27746 31892 27758
rect 32172 27748 32228 27758
rect 31836 27694 31838 27746
rect 31890 27694 31892 27746
rect 31836 26964 31892 27694
rect 32060 27746 32228 27748
rect 32060 27694 32174 27746
rect 32226 27694 32228 27746
rect 32060 27692 32228 27694
rect 31948 26964 32004 26974
rect 31836 26962 32004 26964
rect 31836 26910 31950 26962
rect 32002 26910 32004 26962
rect 31836 26908 32004 26910
rect 31948 26898 32004 26908
rect 32060 26514 32116 27692
rect 32172 27682 32228 27692
rect 32060 26462 32062 26514
rect 32114 26462 32116 26514
rect 32060 26450 32116 26462
rect 31388 25508 31444 25518
rect 31388 24836 31444 25452
rect 31388 24770 31444 24780
rect 32060 25506 32116 25518
rect 32060 25454 32062 25506
rect 32114 25454 32116 25506
rect 31612 23714 31668 23726
rect 31612 23662 31614 23714
rect 31666 23662 31668 23714
rect 31612 21588 31668 23662
rect 32060 23716 32116 25454
rect 32060 23650 32116 23660
rect 32060 23378 32116 23390
rect 32060 23326 32062 23378
rect 32114 23326 32116 23378
rect 32060 23268 32116 23326
rect 32060 23202 32116 23212
rect 32284 23044 32340 31500
rect 32732 31490 32788 31500
rect 32956 30994 33012 31726
rect 32956 30942 32958 30994
rect 33010 30942 33012 30994
rect 32956 30210 33012 30942
rect 33068 30324 33124 31892
rect 33740 31892 33796 32622
rect 34076 31948 34132 33070
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34076 31892 35028 31948
rect 33740 31826 33796 31836
rect 33404 31780 33460 31790
rect 33404 31686 33460 31724
rect 33628 30994 33684 31006
rect 33628 30942 33630 30994
rect 33682 30942 33684 30994
rect 33068 30258 33124 30268
rect 33180 30884 33236 30894
rect 32956 30158 32958 30210
rect 33010 30158 33012 30210
rect 32732 29988 32788 29998
rect 32732 29986 32900 29988
rect 32732 29934 32734 29986
rect 32786 29934 32900 29986
rect 32732 29932 32900 29934
rect 32732 29922 32788 29932
rect 32620 29426 32676 29438
rect 32620 29374 32622 29426
rect 32674 29374 32676 29426
rect 32620 29316 32676 29374
rect 32620 29250 32676 29260
rect 32396 28532 32452 28542
rect 32396 27860 32452 28476
rect 32396 27766 32452 27804
rect 32508 28084 32564 28094
rect 32396 23714 32452 23726
rect 32396 23662 32398 23714
rect 32450 23662 32452 23714
rect 32396 23380 32452 23662
rect 32396 23314 32452 23324
rect 32284 22988 32452 23044
rect 31612 21522 31668 21532
rect 32284 22148 32340 22158
rect 31500 21364 31556 21374
rect 31500 21362 31892 21364
rect 31500 21310 31502 21362
rect 31554 21310 31892 21362
rect 31500 21308 31892 21310
rect 31500 21298 31556 21308
rect 31500 20578 31556 20590
rect 31500 20526 31502 20578
rect 31554 20526 31556 20578
rect 31276 20356 31332 20366
rect 31052 19294 31054 19346
rect 31106 19294 31108 19346
rect 31052 19282 31108 19294
rect 31164 20244 31220 20254
rect 30828 18286 30830 18338
rect 30882 18286 30884 18338
rect 30828 18274 30884 18286
rect 30716 16718 30718 16770
rect 30770 16718 30772 16770
rect 30716 16706 30772 16718
rect 31164 15202 31220 20188
rect 31164 15150 31166 15202
rect 31218 15150 31220 15202
rect 31164 15138 31220 15150
rect 30156 14590 30158 14642
rect 30210 14590 30212 14642
rect 30156 14578 30212 14590
rect 26348 14366 26350 14418
rect 26402 14366 26404 14418
rect 26348 14354 26404 14366
rect 31276 14418 31332 20300
rect 31500 17554 31556 20526
rect 31836 18564 31892 21308
rect 32284 20690 32340 22092
rect 32396 21812 32452 22988
rect 32396 21746 32452 21756
rect 32284 20638 32286 20690
rect 32338 20638 32340 20690
rect 32284 20626 32340 20638
rect 32396 21588 32452 21598
rect 31836 18508 32116 18564
rect 31500 17502 31502 17554
rect 31554 17502 31556 17554
rect 31500 17490 31556 17502
rect 31836 18228 31892 18238
rect 31836 16212 31892 18172
rect 31948 16212 32004 16222
rect 31836 16210 32004 16212
rect 31836 16158 31950 16210
rect 32002 16158 32004 16210
rect 31836 16156 32004 16158
rect 31948 16146 32004 16156
rect 32060 15426 32116 18508
rect 32396 17778 32452 21532
rect 32508 21476 32564 28028
rect 32732 26852 32788 26862
rect 32732 26758 32788 26796
rect 32620 26068 32676 26078
rect 32620 26066 32788 26068
rect 32620 26014 32622 26066
rect 32674 26014 32788 26066
rect 32620 26012 32788 26014
rect 32620 26002 32676 26012
rect 32508 21410 32564 21420
rect 32620 22930 32676 22942
rect 32620 22878 32622 22930
rect 32674 22878 32676 22930
rect 32620 20468 32676 22878
rect 32620 20402 32676 20412
rect 32396 17726 32398 17778
rect 32450 17726 32452 17778
rect 32396 17714 32452 17726
rect 32732 16996 32788 26012
rect 32844 22148 32900 29932
rect 32956 29316 33012 30158
rect 33068 29988 33124 29998
rect 33068 29538 33124 29932
rect 33068 29486 33070 29538
rect 33122 29486 33124 29538
rect 33068 29474 33124 29486
rect 33068 29316 33124 29326
rect 32956 29260 33068 29316
rect 33068 29250 33124 29260
rect 33180 28082 33236 30828
rect 33516 30212 33572 30222
rect 33516 30118 33572 30156
rect 33180 28030 33182 28082
rect 33234 28030 33236 28082
rect 33180 28018 33236 28030
rect 33292 29428 33348 29438
rect 33292 27972 33348 29372
rect 33404 29314 33460 29326
rect 33404 29262 33406 29314
rect 33458 29262 33460 29314
rect 33404 28756 33460 29262
rect 33404 28690 33460 28700
rect 33628 28644 33684 30942
rect 33740 29652 33796 29662
rect 33740 29538 33796 29596
rect 33740 29486 33742 29538
rect 33794 29486 33796 29538
rect 33740 29474 33796 29486
rect 33964 29426 34020 29438
rect 33964 29374 33966 29426
rect 34018 29374 34020 29426
rect 33964 28756 34020 29374
rect 33964 28690 34020 28700
rect 34636 29316 34692 29326
rect 33628 28588 33796 28644
rect 33628 28420 33684 28430
rect 33292 27916 33572 27972
rect 32956 26066 33012 26078
rect 32956 26014 32958 26066
rect 33010 26014 33012 26066
rect 32956 23604 33012 26014
rect 32956 23538 33012 23548
rect 33068 23268 33124 23278
rect 33068 23174 33124 23212
rect 33292 23154 33348 23166
rect 33292 23102 33294 23154
rect 33346 23102 33348 23154
rect 33292 23044 33348 23102
rect 33292 22978 33348 22988
rect 33068 22372 33124 22382
rect 33068 22278 33124 22316
rect 33404 22370 33460 22382
rect 33404 22318 33406 22370
rect 33458 22318 33460 22370
rect 32844 22092 33348 22148
rect 33180 20132 33236 20142
rect 33292 20132 33348 22092
rect 33404 21588 33460 22318
rect 33404 21522 33460 21532
rect 33180 20130 33348 20132
rect 33180 20078 33182 20130
rect 33234 20078 33348 20130
rect 33180 20076 33348 20078
rect 33404 21364 33460 21374
rect 33180 20066 33236 20076
rect 32732 16930 32788 16940
rect 33292 15988 33348 15998
rect 33404 15988 33460 21308
rect 33516 19346 33572 27916
rect 33628 27970 33684 28364
rect 33628 27918 33630 27970
rect 33682 27918 33684 27970
rect 33628 27906 33684 27918
rect 33740 27636 33796 28588
rect 34076 28642 34132 28654
rect 34636 28644 34692 29260
rect 34076 28590 34078 28642
rect 34130 28590 34132 28642
rect 33852 27860 33908 27870
rect 33852 27766 33908 27804
rect 33740 27580 33908 27636
rect 33516 19294 33518 19346
rect 33570 19294 33572 19346
rect 33516 19282 33572 19294
rect 33628 26852 33684 26862
rect 33628 18562 33684 26796
rect 33740 26516 33796 26526
rect 33740 26422 33796 26460
rect 33852 23940 33908 27580
rect 33964 27188 34020 27198
rect 34076 27188 34132 28590
rect 34412 28642 34692 28644
rect 34412 28590 34638 28642
rect 34690 28590 34692 28642
rect 34412 28588 34692 28590
rect 34412 27858 34468 28588
rect 34636 28578 34692 28588
rect 34860 28530 34916 28542
rect 34860 28478 34862 28530
rect 34914 28478 34916 28530
rect 34412 27806 34414 27858
rect 34466 27806 34468 27858
rect 34412 27794 34468 27806
rect 34748 27858 34804 27870
rect 34748 27806 34750 27858
rect 34802 27806 34804 27858
rect 34076 27132 34692 27188
rect 33964 27094 34020 27132
rect 34524 26964 34580 26974
rect 34524 25282 34580 26908
rect 34524 25230 34526 25282
rect 34578 25230 34580 25282
rect 34524 25218 34580 25230
rect 34076 24836 34132 24846
rect 34132 24780 34356 24836
rect 34076 24742 34132 24780
rect 34300 23940 34356 24780
rect 34636 24164 34692 27132
rect 34748 26740 34804 27806
rect 34748 26674 34804 26684
rect 34748 26516 34804 26526
rect 34860 26516 34916 28478
rect 34972 26962 35028 31892
rect 35868 31554 35924 33182
rect 36092 33236 36148 33294
rect 36092 33170 36148 33180
rect 36540 33348 36596 33358
rect 36764 33348 36820 34078
rect 37436 34132 37492 34142
rect 37436 34038 37492 34076
rect 36596 33292 36820 33348
rect 38556 33346 38612 34972
rect 38556 33294 38558 33346
rect 38610 33294 38612 33346
rect 36092 32564 36148 32574
rect 36092 32470 36148 32508
rect 36540 32564 36596 33292
rect 37324 33236 37380 33246
rect 36764 32564 36820 32574
rect 36540 32562 36820 32564
rect 36540 32510 36542 32562
rect 36594 32510 36766 32562
rect 36818 32510 36820 32562
rect 36540 32508 36820 32510
rect 36540 32498 36596 32508
rect 36764 32498 36820 32508
rect 36988 31892 37044 31902
rect 36988 31798 37044 31836
rect 36540 31780 36596 31790
rect 36540 31686 36596 31724
rect 37324 31668 37380 33180
rect 37436 32564 37492 32574
rect 37436 32470 37492 32508
rect 38556 31948 38612 33294
rect 38668 32340 38724 36430
rect 38892 36484 38948 36494
rect 38892 35922 38948 36428
rect 38892 35870 38894 35922
rect 38946 35870 38948 35922
rect 38892 35858 38948 35870
rect 39340 33012 39396 36990
rect 39676 36596 39732 37100
rect 39676 36530 39732 36540
rect 40124 37154 40180 37166
rect 40124 37102 40126 37154
rect 40178 37102 40180 37154
rect 40124 36372 40180 37102
rect 40348 37156 40404 37166
rect 40348 37062 40404 37100
rect 41020 36596 41076 38612
rect 41356 37156 41412 38892
rect 41580 38834 41636 39004
rect 41580 38782 41582 38834
rect 41634 38782 41636 38834
rect 41580 38770 41636 38782
rect 41804 38052 41860 38062
rect 41804 37266 41860 37996
rect 41804 37214 41806 37266
rect 41858 37214 41860 37266
rect 41804 37156 41860 37214
rect 41356 37154 41860 37156
rect 41356 37102 41358 37154
rect 41410 37102 41860 37154
rect 41356 37100 41860 37102
rect 41356 37090 41412 37100
rect 41692 36708 41748 36718
rect 41692 36614 41748 36652
rect 40124 36306 40180 36316
rect 40908 36372 40964 36382
rect 40908 36278 40964 36316
rect 41020 35698 41076 36540
rect 41020 35646 41022 35698
rect 41074 35646 41076 35698
rect 39900 34354 39956 34366
rect 39900 34302 39902 34354
rect 39954 34302 39956 34354
rect 39900 33460 39956 34302
rect 41020 34130 41076 35646
rect 41468 35700 41524 35710
rect 41468 35606 41524 35644
rect 41020 34078 41022 34130
rect 41074 34078 41076 34130
rect 41020 34066 41076 34078
rect 41132 35140 41188 35150
rect 41132 34132 41188 35084
rect 41804 34804 41860 37100
rect 41916 36932 41972 40238
rect 42700 39730 42756 39742
rect 42700 39678 42702 39730
rect 42754 39678 42756 39730
rect 42700 38836 42756 39678
rect 42700 38770 42756 38780
rect 42700 38276 42756 38286
rect 42812 38276 42868 40460
rect 42700 38274 42868 38276
rect 42700 38222 42702 38274
rect 42754 38222 42868 38274
rect 42700 38220 42868 38222
rect 42924 40514 42980 40526
rect 42924 40462 42926 40514
rect 42978 40462 42980 40514
rect 42924 38276 42980 40462
rect 42700 38210 42756 38220
rect 42924 38210 42980 38220
rect 43036 38724 43092 38734
rect 42140 37940 42196 37950
rect 42140 37826 42196 37884
rect 42924 37940 42980 37950
rect 42924 37846 42980 37884
rect 42140 37774 42142 37826
rect 42194 37774 42196 37826
rect 42140 37762 42196 37774
rect 41916 36866 41972 36876
rect 43036 36932 43092 38668
rect 43036 36866 43092 36876
rect 43148 38050 43204 40908
rect 43708 40852 43764 41020
rect 43708 40786 43764 40796
rect 43708 40516 43764 40526
rect 43820 40516 43876 41356
rect 43932 41300 43988 42142
rect 44492 41972 44548 41982
rect 44604 41972 44660 43652
rect 44940 43540 44996 45948
rect 45388 45332 45444 46734
rect 46060 46116 46116 50652
rect 46172 49700 46228 49710
rect 46172 49606 46228 49644
rect 46284 47348 46340 52220
rect 48412 52274 48692 52276
rect 48412 52222 48638 52274
rect 48690 52222 48692 52274
rect 48412 52220 48692 52222
rect 47180 52052 47236 52062
rect 47180 52050 47460 52052
rect 47180 51998 47182 52050
rect 47234 51998 47460 52050
rect 47180 51996 47460 51998
rect 47180 51986 47236 51996
rect 47068 50484 47124 50494
rect 47068 50390 47124 50428
rect 46844 49924 46900 49934
rect 46844 49830 46900 49868
rect 46396 49810 46452 49822
rect 46396 49758 46398 49810
rect 46450 49758 46452 49810
rect 46396 49700 46452 49758
rect 46396 48916 46452 49644
rect 47068 49810 47124 49822
rect 47068 49758 47070 49810
rect 47122 49758 47124 49810
rect 47068 49700 47124 49758
rect 47068 49634 47124 49644
rect 46396 48850 46452 48860
rect 45388 45266 45444 45276
rect 45500 46060 46116 46116
rect 46172 47292 46340 47348
rect 46508 48804 46564 48814
rect 45164 45220 45220 45230
rect 45164 44434 45220 45164
rect 45500 45106 45556 46060
rect 45724 45668 45780 45678
rect 45724 45574 45780 45612
rect 46172 45444 46228 47292
rect 46172 45378 46228 45388
rect 46284 47124 46340 47134
rect 46284 45778 46340 47068
rect 46284 45726 46286 45778
rect 46338 45726 46340 45778
rect 45500 45054 45502 45106
rect 45554 45054 45556 45106
rect 45500 45042 45556 45054
rect 45948 45108 46004 45118
rect 46284 45108 46340 45726
rect 46508 45220 46564 48748
rect 45948 45106 46340 45108
rect 45948 45054 45950 45106
rect 46002 45054 46340 45106
rect 45948 45052 46340 45054
rect 46396 45164 46564 45220
rect 46844 46900 46900 46910
rect 46844 45218 46900 46844
rect 47292 45332 47348 45342
rect 47292 45238 47348 45276
rect 46844 45166 46846 45218
rect 46898 45166 46900 45218
rect 45164 44382 45166 44434
rect 45218 44382 45220 44434
rect 45164 44370 45220 44382
rect 45388 44322 45444 44334
rect 45388 44270 45390 44322
rect 45442 44270 45444 44322
rect 45388 44212 45444 44270
rect 45948 44322 46004 45052
rect 45948 44270 45950 44322
rect 46002 44270 46004 44322
rect 45444 44156 45556 44212
rect 45388 44146 45444 44156
rect 45388 43988 45444 43998
rect 45164 43540 45220 43550
rect 44940 43538 45220 43540
rect 44940 43486 45166 43538
rect 45218 43486 45220 43538
rect 44940 43484 45220 43486
rect 44940 42756 44996 42766
rect 44492 41970 44660 41972
rect 44492 41918 44494 41970
rect 44546 41918 44660 41970
rect 44492 41916 44660 41918
rect 44828 41972 44884 41982
rect 44940 41972 44996 42700
rect 44828 41970 44996 41972
rect 44828 41918 44830 41970
rect 44882 41918 44996 41970
rect 44828 41916 44996 41918
rect 44492 41906 44548 41916
rect 44828 41906 44884 41916
rect 43932 41234 43988 41244
rect 44828 41076 44884 41086
rect 43708 40514 43876 40516
rect 43708 40462 43710 40514
rect 43762 40462 43876 40514
rect 43708 40460 43876 40462
rect 43932 41074 44884 41076
rect 43932 41022 44830 41074
rect 44882 41022 44884 41074
rect 43932 41020 44884 41022
rect 43708 40450 43764 40460
rect 43708 39620 43764 39630
rect 43708 38162 43764 39564
rect 43932 39058 43988 41020
rect 44828 41010 44884 41020
rect 44044 40852 44100 40862
rect 44044 40514 44100 40796
rect 44044 40462 44046 40514
rect 44098 40462 44100 40514
rect 44044 40450 44100 40462
rect 44492 40402 44548 40414
rect 44492 40350 44494 40402
rect 44546 40350 44548 40402
rect 44492 39732 44548 40350
rect 44940 40404 44996 40414
rect 44940 40310 44996 40348
rect 44492 39666 44548 39676
rect 44940 39618 44996 39630
rect 44940 39566 44942 39618
rect 44994 39566 44996 39618
rect 44044 39508 44100 39518
rect 44044 39506 44660 39508
rect 44044 39454 44046 39506
rect 44098 39454 44660 39506
rect 44044 39452 44660 39454
rect 44044 39442 44100 39452
rect 43932 39006 43934 39058
rect 43986 39006 43988 39058
rect 43932 38994 43988 39006
rect 44604 39058 44660 39452
rect 44604 39006 44606 39058
rect 44658 39006 44660 39058
rect 44604 38994 44660 39006
rect 43708 38110 43710 38162
rect 43762 38110 43764 38162
rect 43708 38098 43764 38110
rect 44380 38836 44436 38846
rect 43148 37998 43150 38050
rect 43202 37998 43204 38050
rect 43148 37940 43204 37998
rect 43148 37156 43204 37884
rect 43820 38050 43876 38062
rect 43820 37998 43822 38050
rect 43874 37998 43876 38050
rect 43820 37940 43876 37998
rect 43820 37874 43876 37884
rect 42028 36596 42084 36606
rect 42028 36502 42084 36540
rect 42812 36596 42868 36606
rect 42812 36502 42868 36540
rect 43148 36594 43204 37100
rect 43148 36542 43150 36594
rect 43202 36542 43204 36594
rect 43148 36530 43204 36542
rect 44380 36594 44436 38780
rect 44940 38722 44996 39566
rect 45052 38836 45108 43484
rect 45164 43428 45220 43484
rect 45164 43362 45220 43372
rect 45388 42754 45444 43932
rect 45500 43708 45556 44156
rect 45948 43876 46004 44270
rect 46396 43988 46452 45164
rect 46844 45154 46900 45166
rect 46508 44996 46564 45006
rect 46508 44902 46564 44940
rect 47180 44996 47236 45006
rect 47180 44902 47236 44940
rect 46620 44324 46676 44334
rect 46620 44230 46676 44268
rect 46396 43922 46452 43932
rect 45948 43810 46004 43820
rect 45500 43652 45780 43708
rect 45388 42702 45390 42754
rect 45442 42702 45444 42754
rect 45388 42690 45444 42702
rect 45724 43426 45780 43652
rect 47404 43540 47460 51996
rect 48412 49812 48468 52220
rect 48636 52210 48692 52220
rect 48636 52052 48692 52062
rect 48412 49746 48468 49756
rect 48524 51996 48636 52052
rect 47516 49700 47572 49710
rect 47516 49606 47572 49644
rect 47852 49698 47908 49710
rect 47852 49646 47854 49698
rect 47906 49646 47908 49698
rect 47852 48914 47908 49646
rect 47852 48862 47854 48914
rect 47906 48862 47908 48914
rect 47852 48850 47908 48862
rect 47964 49700 48020 49710
rect 47740 48692 47796 48702
rect 47628 47234 47684 47246
rect 47628 47182 47630 47234
rect 47682 47182 47684 47234
rect 47628 46900 47684 47182
rect 47628 46834 47684 46844
rect 47740 46674 47796 48636
rect 47964 48132 48020 49644
rect 48412 48916 48468 48926
rect 47964 48130 48244 48132
rect 47964 48078 47966 48130
rect 48018 48078 48244 48130
rect 47964 48076 48244 48078
rect 47964 48066 48020 48076
rect 47740 46622 47742 46674
rect 47794 46622 47796 46674
rect 47740 46610 47796 46622
rect 48076 47124 48132 47134
rect 48076 46674 48132 47068
rect 48076 46622 48078 46674
rect 48130 46622 48132 46674
rect 48076 46610 48132 46622
rect 48188 45332 48244 48076
rect 48412 47682 48468 48860
rect 48524 48468 48580 51996
rect 48636 51986 48692 51996
rect 48636 50708 48692 50746
rect 48636 50642 48692 50652
rect 48636 50484 48692 50494
rect 48636 49250 48692 50428
rect 48636 49198 48638 49250
rect 48690 49198 48692 49250
rect 48636 49186 48692 49198
rect 48636 48468 48692 48478
rect 48524 48466 48692 48468
rect 48524 48414 48638 48466
rect 48690 48414 48692 48466
rect 48524 48412 48692 48414
rect 48636 48402 48692 48412
rect 48412 47630 48414 47682
rect 48466 47630 48468 47682
rect 48412 47618 48468 47630
rect 48524 47458 48580 47470
rect 48524 47406 48526 47458
rect 48578 47406 48580 47458
rect 48524 47124 48580 47406
rect 49196 47458 49252 52780
rect 50092 52770 50148 52780
rect 51100 52164 51156 53006
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 51100 52098 51156 52108
rect 49868 52050 49924 52062
rect 49868 51998 49870 52050
rect 49922 51998 49924 52050
rect 49756 51266 49812 51278
rect 49756 51214 49758 51266
rect 49810 51214 49812 51266
rect 49644 50484 49700 50494
rect 49196 47406 49198 47458
rect 49250 47406 49252 47458
rect 49196 47394 49252 47406
rect 49308 50482 49700 50484
rect 49308 50430 49646 50482
rect 49698 50430 49700 50482
rect 49308 50428 49700 50430
rect 49308 47236 49364 50428
rect 49644 50418 49700 50428
rect 49420 49700 49476 49710
rect 49644 49700 49700 49710
rect 49420 49606 49476 49644
rect 49532 49698 49700 49700
rect 49532 49646 49646 49698
rect 49698 49646 49700 49698
rect 49532 49644 49700 49646
rect 49420 48468 49476 48478
rect 49532 48468 49588 49644
rect 49644 49634 49700 49644
rect 49756 48692 49812 51214
rect 49868 49588 49924 51998
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50764 51492 50820 51502
rect 50764 51398 50820 51436
rect 53788 51490 53844 51502
rect 53788 51438 53790 51490
rect 53842 51438 53844 51490
rect 52556 51266 52612 51278
rect 52556 51214 52558 51266
rect 52610 51214 52612 51266
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50316 49810 50372 49822
rect 50316 49758 50318 49810
rect 50370 49758 50372 49810
rect 49980 49700 50036 49710
rect 49980 49606 50036 49644
rect 49868 49522 49924 49532
rect 49868 49138 49924 49150
rect 49868 49086 49870 49138
rect 49922 49086 49924 49138
rect 49868 48804 49924 49086
rect 49868 48738 49924 48748
rect 49756 48626 49812 48636
rect 49420 48466 49588 48468
rect 49420 48414 49422 48466
rect 49474 48414 49588 48466
rect 49420 48412 49588 48414
rect 49420 48402 49476 48412
rect 49532 48132 49588 48142
rect 49308 47170 49364 47180
rect 49420 47460 49476 47470
rect 48524 46676 48580 47068
rect 48636 46676 48692 46686
rect 48524 46674 48692 46676
rect 48524 46622 48638 46674
rect 48690 46622 48692 46674
rect 48524 46620 48692 46622
rect 48636 46610 48692 46620
rect 49308 46674 49364 46686
rect 49308 46622 49310 46674
rect 49362 46622 49364 46674
rect 49308 46004 49364 46622
rect 49308 45938 49364 45948
rect 48188 45238 48244 45276
rect 48860 45106 48916 45118
rect 48860 45054 48862 45106
rect 48914 45054 48916 45106
rect 48860 43764 48916 45054
rect 49308 45108 49364 45118
rect 49420 45108 49476 47404
rect 49308 45106 49476 45108
rect 49308 45054 49310 45106
rect 49362 45054 49476 45106
rect 49308 45052 49476 45054
rect 49308 45042 49364 45052
rect 49532 44884 49588 48076
rect 49308 44828 49588 44884
rect 49644 46228 49700 46238
rect 49084 44100 49140 44110
rect 49084 44098 49252 44100
rect 49084 44046 49086 44098
rect 49138 44046 49252 44098
rect 49084 44044 49252 44046
rect 49084 44034 49140 44044
rect 49084 43876 49140 43886
rect 48972 43764 49028 43774
rect 48860 43708 48972 43764
rect 47404 43474 47460 43484
rect 47740 43652 47796 43662
rect 45724 43374 45726 43426
rect 45778 43374 45780 43426
rect 45276 41972 45332 41982
rect 45276 41878 45332 41916
rect 45500 41300 45556 41310
rect 45500 41206 45556 41244
rect 45724 41300 45780 43374
rect 47740 42756 47796 43596
rect 48188 43652 48244 43662
rect 48188 43558 48244 43596
rect 48860 43428 48916 43438
rect 48860 43334 48916 43372
rect 46508 42532 46564 42542
rect 46172 41300 46228 41310
rect 45724 41244 46172 41300
rect 45724 41186 45780 41244
rect 46172 41206 46228 41244
rect 46508 41298 46564 42476
rect 47628 42532 47684 42542
rect 47628 42438 47684 42476
rect 47516 42084 47572 42094
rect 47180 42082 47572 42084
rect 47180 42030 47518 42082
rect 47570 42030 47572 42082
rect 47180 42028 47572 42030
rect 46508 41246 46510 41298
rect 46562 41246 46564 41298
rect 46508 41234 46564 41246
rect 46844 41300 46900 41310
rect 46844 41206 46900 41244
rect 47180 41298 47236 42028
rect 47516 42018 47572 42028
rect 47180 41246 47182 41298
rect 47234 41246 47236 41298
rect 47180 41234 47236 41246
rect 45724 41134 45726 41186
rect 45778 41134 45780 41186
rect 45164 41076 45220 41086
rect 45164 40982 45220 41020
rect 45724 40852 45780 41134
rect 47628 41188 47684 41198
rect 47740 41188 47796 42700
rect 48300 43204 48356 43214
rect 48300 41970 48356 43148
rect 48972 42868 49028 43708
rect 48636 42812 49028 42868
rect 48636 42754 48692 42812
rect 48636 42702 48638 42754
rect 48690 42702 48692 42754
rect 48412 42644 48468 42654
rect 48412 42550 48468 42588
rect 48300 41918 48302 41970
rect 48354 41918 48356 41970
rect 48300 41906 48356 41918
rect 48636 41970 48692 42702
rect 49084 42754 49140 43820
rect 49196 43650 49252 44044
rect 49196 43598 49198 43650
rect 49250 43598 49252 43650
rect 49196 43586 49252 43598
rect 49084 42702 49086 42754
rect 49138 42702 49140 42754
rect 49084 42690 49140 42702
rect 49196 43428 49252 43438
rect 48636 41918 48638 41970
rect 48690 41918 48692 41970
rect 48636 41906 48692 41918
rect 47628 41186 47796 41188
rect 47628 41134 47630 41186
rect 47682 41134 47796 41186
rect 47628 41132 47796 41134
rect 48076 41188 48132 41198
rect 47628 41122 47684 41132
rect 48076 41094 48132 41132
rect 45724 40786 45780 40796
rect 47404 40626 47460 40638
rect 47404 40574 47406 40626
rect 47458 40574 47460 40626
rect 45388 39620 45444 39630
rect 45388 39526 45444 39564
rect 45388 39060 45444 39070
rect 45388 38966 45444 39004
rect 47068 38948 47124 38958
rect 47068 38854 47124 38892
rect 45052 38770 45108 38780
rect 44940 38670 44942 38722
rect 44994 38670 44996 38722
rect 44940 38668 44996 38670
rect 44380 36542 44382 36594
rect 44434 36542 44436 36594
rect 44380 36484 44436 36542
rect 44380 36418 44436 36428
rect 44828 38612 44996 38668
rect 45836 38722 45892 38734
rect 45836 38670 45838 38722
rect 45890 38670 45892 38722
rect 44828 38050 44884 38612
rect 44828 37998 44830 38050
rect 44882 37998 44884 38050
rect 44828 37156 44884 37998
rect 45388 38276 45444 38286
rect 45388 38050 45444 38220
rect 45388 37998 45390 38050
rect 45442 37998 45444 38050
rect 45388 37986 45444 37998
rect 44828 36596 44884 37100
rect 45500 37940 45556 37950
rect 45500 37380 45556 37884
rect 43484 36372 43540 36382
rect 43484 36370 43764 36372
rect 43484 36318 43486 36370
rect 43538 36318 43764 36370
rect 43484 36316 43764 36318
rect 43484 36306 43540 36316
rect 43708 35922 43764 36316
rect 43708 35870 43710 35922
rect 43762 35870 43764 35922
rect 43708 35858 43764 35870
rect 44492 35924 44548 35934
rect 44492 35830 44548 35868
rect 44828 35700 44884 36540
rect 44268 35698 44884 35700
rect 44268 35646 44830 35698
rect 44882 35646 44884 35698
rect 44268 35644 44884 35646
rect 44268 35026 44324 35644
rect 44828 35634 44884 35644
rect 45276 36820 45332 36830
rect 45276 35698 45332 36764
rect 45500 36706 45556 37324
rect 45500 36654 45502 36706
rect 45554 36654 45556 36706
rect 45500 36642 45556 36654
rect 45836 36036 45892 38670
rect 47404 38724 47460 40574
rect 47964 40628 48020 40638
rect 47964 40534 48020 40572
rect 49196 40402 49252 43372
rect 49308 41970 49364 44828
rect 49644 44546 49700 46172
rect 49644 44494 49646 44546
rect 49698 44494 49700 44546
rect 49644 44482 49700 44494
rect 49868 45332 49924 45342
rect 49868 44436 49924 45276
rect 49868 44342 49924 44380
rect 50204 45220 50260 45230
rect 50204 44434 50260 45164
rect 50204 44382 50206 44434
rect 50258 44382 50260 44434
rect 50204 44370 50260 44382
rect 49756 44324 49812 44334
rect 49756 43876 49812 44268
rect 49756 43810 49812 43820
rect 50316 43764 50372 49758
rect 50876 49810 50932 49822
rect 50876 49758 50878 49810
rect 50930 49758 50932 49810
rect 50876 49476 50932 49758
rect 50876 49410 50932 49420
rect 51772 49700 51828 49710
rect 50876 48914 50932 48926
rect 51660 48916 51716 48926
rect 50876 48862 50878 48914
rect 50930 48862 50932 48914
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50876 46788 50932 48862
rect 51548 48914 51716 48916
rect 51548 48862 51662 48914
rect 51714 48862 51716 48914
rect 51548 48860 51716 48862
rect 51548 47234 51604 48860
rect 51660 48850 51716 48860
rect 51772 48242 51828 49644
rect 52556 49700 52612 51214
rect 53788 50596 53844 51438
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 53788 50530 53844 50540
rect 54012 50706 54068 50718
rect 54012 50654 54014 50706
rect 54066 50654 54068 50706
rect 53900 50484 53956 50494
rect 53340 50034 53396 50046
rect 53340 49982 53342 50034
rect 53394 49982 53396 50034
rect 53340 49924 53396 49982
rect 53900 50034 53956 50428
rect 53900 49982 53902 50034
rect 53954 49982 53956 50034
rect 53900 49970 53956 49982
rect 53340 49858 53396 49868
rect 52556 49634 52612 49644
rect 51884 49588 51940 49598
rect 51884 49028 51940 49532
rect 53676 49140 53732 49150
rect 53676 49046 53732 49084
rect 51884 48934 51940 48972
rect 52780 49028 52836 49038
rect 52780 48934 52836 48972
rect 53004 49028 53060 49038
rect 51772 48190 51774 48242
rect 51826 48190 51828 48242
rect 51772 48178 51828 48190
rect 52220 48804 52276 48814
rect 52220 47682 52276 48748
rect 52332 48242 52388 48254
rect 52332 48190 52334 48242
rect 52386 48190 52388 48242
rect 52332 48132 52388 48190
rect 52668 48132 52724 48142
rect 52332 48130 52724 48132
rect 52332 48078 52670 48130
rect 52722 48078 52724 48130
rect 52332 48076 52724 48078
rect 52668 48018 52724 48076
rect 52668 47966 52670 48018
rect 52722 47966 52724 48018
rect 52220 47630 52222 47682
rect 52274 47630 52276 47682
rect 52220 47618 52276 47630
rect 52444 47908 52500 47918
rect 51548 47182 51550 47234
rect 51602 47182 51604 47234
rect 51548 47170 51604 47182
rect 52444 46898 52500 47852
rect 52444 46846 52446 46898
rect 52498 46846 52500 46898
rect 52444 46834 52500 46846
rect 52668 47458 52724 47966
rect 52668 47406 52670 47458
rect 52722 47406 52724 47458
rect 51548 46788 51604 46798
rect 50876 46722 50932 46732
rect 51436 46786 51604 46788
rect 51436 46734 51550 46786
rect 51602 46734 51604 46786
rect 51436 46732 51604 46734
rect 50428 45890 50484 45902
rect 50428 45838 50430 45890
rect 50482 45838 50484 45890
rect 50428 45668 50484 45838
rect 50428 45602 50484 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 51436 44996 51492 46732
rect 51548 46722 51604 46732
rect 52220 46564 52276 46574
rect 51884 45668 51940 45678
rect 51660 45666 51940 45668
rect 51660 45614 51886 45666
rect 51938 45614 51940 45666
rect 51660 45612 51940 45614
rect 51548 45220 51604 45230
rect 51548 45126 51604 45164
rect 51436 44940 51604 44996
rect 51100 44436 51156 44446
rect 51436 44436 51492 44446
rect 51156 44434 51492 44436
rect 51156 44382 51438 44434
rect 51490 44382 51492 44434
rect 51156 44380 51492 44382
rect 51100 44342 51156 44380
rect 50652 44100 50708 44110
rect 50652 44098 50932 44100
rect 50652 44046 50654 44098
rect 50706 44046 50932 44098
rect 50652 44044 50932 44046
rect 50652 44034 50708 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50316 43698 50372 43708
rect 49532 43652 49588 43662
rect 49532 43558 49588 43596
rect 49980 43652 50036 43662
rect 49980 43538 50036 43596
rect 50764 43652 50820 43662
rect 50876 43652 50932 44044
rect 50764 43650 50876 43652
rect 50764 43598 50766 43650
rect 50818 43598 50876 43650
rect 50764 43596 50876 43598
rect 50764 43586 50820 43596
rect 50876 43586 50932 43596
rect 49980 43486 49982 43538
rect 50034 43486 50036 43538
rect 49980 43474 50036 43486
rect 50988 43540 51044 43550
rect 50988 43446 51044 43484
rect 51436 43540 51492 44380
rect 51548 44098 51604 44940
rect 51548 44046 51550 44098
rect 51602 44046 51604 44098
rect 51548 44034 51604 44046
rect 51548 43652 51604 43662
rect 51660 43652 51716 45612
rect 51884 45602 51940 45612
rect 51604 43596 51716 43652
rect 51548 43586 51604 43596
rect 51436 43474 51492 43484
rect 50204 43428 50260 43438
rect 50204 43334 50260 43372
rect 51548 43428 51604 43438
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 51548 42194 51604 43372
rect 51660 42756 51716 43596
rect 51772 43652 51828 43662
rect 51772 43558 51828 43596
rect 52220 42978 52276 46508
rect 52332 46452 52388 46462
rect 52332 46358 52388 46396
rect 52668 45892 52724 47406
rect 52892 47572 52948 47582
rect 52556 45890 52836 45892
rect 52556 45838 52670 45890
rect 52722 45838 52836 45890
rect 52556 45836 52836 45838
rect 52332 45780 52388 45790
rect 52332 45330 52388 45724
rect 52332 45278 52334 45330
rect 52386 45278 52388 45330
rect 52332 45266 52388 45278
rect 52556 45106 52612 45836
rect 52668 45826 52724 45836
rect 52556 45054 52558 45106
rect 52610 45054 52612 45106
rect 52556 45042 52612 45054
rect 52668 45668 52724 45678
rect 52668 44996 52724 45612
rect 52220 42926 52222 42978
rect 52274 42926 52276 42978
rect 52220 42914 52276 42926
rect 52332 44884 52388 44894
rect 51660 42700 51828 42756
rect 51548 42142 51550 42194
rect 51602 42142 51604 42194
rect 51548 42130 51604 42142
rect 51660 42530 51716 42542
rect 51660 42478 51662 42530
rect 51714 42478 51716 42530
rect 49308 41918 49310 41970
rect 49362 41918 49364 41970
rect 49308 41906 49364 41918
rect 51436 41300 51492 41310
rect 51436 41188 51492 41244
rect 51660 41298 51716 42478
rect 51660 41246 51662 41298
rect 51714 41246 51716 41298
rect 51660 41234 51716 41246
rect 51772 41300 51828 42700
rect 52332 41970 52388 44828
rect 52668 44322 52724 44940
rect 52668 44270 52670 44322
rect 52722 44270 52724 44322
rect 52332 41918 52334 41970
rect 52386 41918 52388 41970
rect 52332 41906 52388 41918
rect 52444 41970 52500 41982
rect 52444 41918 52446 41970
rect 52498 41918 52500 41970
rect 52108 41300 52164 41310
rect 51772 41244 52108 41300
rect 51212 41186 51492 41188
rect 51212 41134 51438 41186
rect 51490 41134 51492 41186
rect 51212 41132 51492 41134
rect 49196 40350 49198 40402
rect 49250 40350 49252 40402
rect 49196 40338 49252 40350
rect 50316 40962 50372 40974
rect 50316 40910 50318 40962
rect 50370 40910 50372 40962
rect 50316 40180 50372 40910
rect 51100 40964 51156 40974
rect 51100 40870 51156 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 51100 40292 51156 40302
rect 51212 40292 51268 41132
rect 51436 41122 51492 41132
rect 51996 40404 52052 41244
rect 52108 41206 52164 41244
rect 51100 40290 51268 40292
rect 51100 40238 51102 40290
rect 51154 40238 51268 40290
rect 51100 40236 51268 40238
rect 51772 40402 52052 40404
rect 51772 40350 51998 40402
rect 52050 40350 52052 40402
rect 51772 40348 52052 40350
rect 51100 40226 51156 40236
rect 50316 40114 50372 40124
rect 51436 40180 51492 40190
rect 50204 40068 50260 40078
rect 48412 39956 48468 39966
rect 48412 39842 48468 39900
rect 48412 39790 48414 39842
rect 48466 39790 48468 39842
rect 48412 39778 48468 39790
rect 49196 39732 49252 39742
rect 49252 39676 49588 39732
rect 49196 39638 49252 39676
rect 47852 39394 47908 39406
rect 47852 39342 47854 39394
rect 47906 39342 47908 39394
rect 47404 38658 47460 38668
rect 47740 38722 47796 38734
rect 47740 38670 47742 38722
rect 47794 38670 47796 38722
rect 47628 37826 47684 37838
rect 47628 37774 47630 37826
rect 47682 37774 47684 37826
rect 47292 37380 47348 37390
rect 47292 37286 47348 37324
rect 47628 37378 47684 37774
rect 47628 37326 47630 37378
rect 47682 37326 47684 37378
rect 47628 37314 47684 37326
rect 46732 37156 46788 37166
rect 45836 35970 45892 35980
rect 46396 36596 46452 36606
rect 45276 35646 45278 35698
rect 45330 35646 45332 35698
rect 45276 35634 45332 35646
rect 44268 34974 44270 35026
rect 44322 34974 44324 35026
rect 44268 34962 44324 34974
rect 46060 34914 46116 34926
rect 46060 34862 46062 34914
rect 46114 34862 46116 34914
rect 41804 34738 41860 34748
rect 42924 34804 42980 34814
rect 42924 34710 42980 34748
rect 43596 34804 43652 34814
rect 43596 34690 43652 34748
rect 43596 34638 43598 34690
rect 43650 34638 43652 34690
rect 40460 33908 40516 33918
rect 40460 33814 40516 33852
rect 39900 33394 39956 33404
rect 40348 33348 40404 33358
rect 40348 33234 40404 33292
rect 40348 33182 40350 33234
rect 40402 33182 40404 33234
rect 40348 33170 40404 33182
rect 39340 32946 39396 32956
rect 39900 33124 39956 33134
rect 39900 32786 39956 33068
rect 39900 32734 39902 32786
rect 39954 32734 39956 32786
rect 39900 32722 39956 32734
rect 41132 32786 41188 34076
rect 41468 34132 41524 34142
rect 41468 34038 41524 34076
rect 41916 33572 41972 33582
rect 41132 32734 41134 32786
rect 41186 32734 41188 32786
rect 41132 32722 41188 32734
rect 41244 33348 41300 33358
rect 41244 32562 41300 33292
rect 41244 32510 41246 32562
rect 41298 32510 41300 32562
rect 38668 32274 38724 32284
rect 40460 32338 40516 32350
rect 40460 32286 40462 32338
rect 40514 32286 40516 32338
rect 38444 31892 38612 31948
rect 40460 32004 40516 32286
rect 40460 31938 40516 31948
rect 37324 31574 37380 31612
rect 38220 31778 38276 31790
rect 38220 31726 38222 31778
rect 38274 31726 38276 31778
rect 35868 31502 35870 31554
rect 35922 31502 35924 31554
rect 35868 31490 35924 31502
rect 37772 31554 37828 31566
rect 37772 31502 37774 31554
rect 37826 31502 37828 31554
rect 37324 31332 37380 31342
rect 36092 31220 36148 31230
rect 36092 31126 36148 31164
rect 37324 30994 37380 31276
rect 37772 31332 37828 31502
rect 37772 31266 37828 31276
rect 37324 30942 37326 30994
rect 37378 30942 37380 30994
rect 37324 30930 37380 30942
rect 36652 30772 36708 30782
rect 36652 30678 36708 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35644 30324 35700 30334
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28642 35140 28654
rect 35084 28590 35086 28642
rect 35138 28590 35140 28642
rect 35084 27860 35140 28590
rect 35084 27794 35140 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34972 26910 34974 26962
rect 35026 26910 35028 26962
rect 34972 26898 35028 26910
rect 35644 26964 35700 30268
rect 37100 30210 37156 30222
rect 37100 30158 37102 30210
rect 37154 30158 37156 30210
rect 35980 29986 36036 29998
rect 35980 29934 35982 29986
rect 36034 29934 36036 29986
rect 35980 28756 36036 29934
rect 36540 29988 36596 29998
rect 36540 29986 36820 29988
rect 36540 29934 36542 29986
rect 36594 29934 36820 29986
rect 36540 29932 36820 29934
rect 36540 29922 36596 29932
rect 36204 29428 36260 29438
rect 36204 29334 36260 29372
rect 36092 28756 36148 28766
rect 35980 28754 36148 28756
rect 35980 28702 36094 28754
rect 36146 28702 36148 28754
rect 35980 28700 36148 28702
rect 36092 28690 36148 28700
rect 36316 28756 36372 28766
rect 36316 28642 36372 28700
rect 36316 28590 36318 28642
rect 36370 28590 36372 28642
rect 36316 28578 36372 28590
rect 35756 27860 35812 27870
rect 35756 27186 35812 27804
rect 36764 27300 36820 29932
rect 37100 29316 37156 30158
rect 37100 29250 37156 29260
rect 37548 30210 37604 30222
rect 37548 30158 37550 30210
rect 37602 30158 37604 30210
rect 36876 28644 36932 28654
rect 36876 28642 37044 28644
rect 36876 28590 36878 28642
rect 36930 28590 37044 28642
rect 36876 28588 37044 28590
rect 36876 28578 36932 28588
rect 36988 27412 37044 28588
rect 37548 28196 37604 30158
rect 38220 30212 38276 31726
rect 38220 30146 38276 30156
rect 38332 31668 38388 31678
rect 38332 30996 38388 31612
rect 38332 30770 38388 30940
rect 38332 30718 38334 30770
rect 38386 30718 38388 30770
rect 38332 28756 38388 30718
rect 38444 29428 38500 31892
rect 38668 31778 38724 31790
rect 38668 31726 38670 31778
rect 38722 31726 38724 31778
rect 38668 30884 38724 31726
rect 41132 31668 41188 31678
rect 41132 31554 41188 31612
rect 41132 31502 41134 31554
rect 41186 31502 41188 31554
rect 41132 31490 41188 31502
rect 39900 31220 39956 31230
rect 39900 31126 39956 31164
rect 39788 30996 39844 31006
rect 39788 30902 39844 30940
rect 41020 30996 41076 31006
rect 41244 30996 41300 32510
rect 41916 32562 41972 33516
rect 42924 33460 42980 33470
rect 42924 33366 42980 33404
rect 43260 33460 43316 33470
rect 41916 32510 41918 32562
rect 41970 32510 41972 32562
rect 41916 32498 41972 32510
rect 42924 32900 42980 32910
rect 42924 31890 42980 32844
rect 43260 31892 43316 33404
rect 42924 31838 42926 31890
rect 42978 31838 42980 31890
rect 42924 31826 42980 31838
rect 43036 31890 43316 31892
rect 43036 31838 43262 31890
rect 43314 31838 43316 31890
rect 43036 31836 43316 31838
rect 42252 31780 42308 31790
rect 42700 31780 42756 31790
rect 42252 31778 42756 31780
rect 42252 31726 42254 31778
rect 42306 31726 42702 31778
rect 42754 31726 42756 31778
rect 42252 31724 42756 31726
rect 42252 31714 42308 31724
rect 41692 31666 41748 31678
rect 41692 31614 41694 31666
rect 41746 31614 41748 31666
rect 41692 31556 41748 31614
rect 41916 31668 41972 31678
rect 42700 31668 42756 31724
rect 43036 31668 43092 31836
rect 43260 31826 43316 31836
rect 42700 31612 43092 31668
rect 41916 31574 41972 31612
rect 41692 31490 41748 31500
rect 43372 31556 43428 31566
rect 43372 31462 43428 31500
rect 41020 30994 41300 30996
rect 41020 30942 41022 30994
rect 41074 30942 41300 30994
rect 41020 30940 41300 30942
rect 41468 30996 41524 31006
rect 41020 30930 41076 30940
rect 41468 30902 41524 30940
rect 38668 30818 38724 30828
rect 40684 30212 40740 30222
rect 41244 30212 41300 30222
rect 40012 29988 40068 29998
rect 40012 29894 40068 29932
rect 40572 29986 40628 29998
rect 40572 29934 40574 29986
rect 40626 29934 40628 29986
rect 38444 29362 38500 29372
rect 38892 29428 38948 29438
rect 37660 28420 37716 28430
rect 37660 28326 37716 28364
rect 37548 28130 37604 28140
rect 37324 28082 37380 28094
rect 37324 28030 37326 28082
rect 37378 28030 37380 28082
rect 37324 27972 37380 28030
rect 38108 27972 38164 27982
rect 37324 27970 38164 27972
rect 37324 27918 38110 27970
rect 38162 27918 38164 27970
rect 37324 27916 38164 27918
rect 38108 27906 38164 27916
rect 38332 27858 38388 28700
rect 38332 27806 38334 27858
rect 38386 27806 38388 27858
rect 38332 27794 38388 27806
rect 38556 29316 38612 29326
rect 37884 27636 37940 27646
rect 37884 27634 38500 27636
rect 37884 27582 37886 27634
rect 37938 27582 38500 27634
rect 37884 27580 38500 27582
rect 37884 27570 37940 27580
rect 36988 27356 37380 27412
rect 36764 27244 37268 27300
rect 35756 27134 35758 27186
rect 35810 27134 35812 27186
rect 35756 27122 35812 27134
rect 37100 27076 37156 27086
rect 37100 26982 37156 27020
rect 36092 26964 36148 26974
rect 35644 26908 35812 26964
rect 35756 26852 35924 26908
rect 36092 26870 36148 26908
rect 34804 26460 34916 26516
rect 34748 26450 34804 26460
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35084 25284 35140 25294
rect 34860 25282 35140 25284
rect 34860 25230 35086 25282
rect 35138 25230 35140 25282
rect 34860 25228 35140 25230
rect 34636 24108 34804 24164
rect 33852 23884 34244 23940
rect 34076 23716 34132 23726
rect 33740 23380 33796 23390
rect 33740 23266 33796 23324
rect 33740 23214 33742 23266
rect 33794 23214 33796 23266
rect 33740 23202 33796 23214
rect 33964 23154 34020 23166
rect 33964 23102 33966 23154
rect 34018 23102 34020 23154
rect 33964 23044 34020 23102
rect 33964 22978 34020 22988
rect 34076 21924 34132 23660
rect 34188 22036 34244 23884
rect 34300 23154 34356 23884
rect 34636 23938 34692 23950
rect 34636 23886 34638 23938
rect 34690 23886 34692 23938
rect 34300 23102 34302 23154
rect 34354 23102 34356 23154
rect 34300 22372 34356 23102
rect 34300 22306 34356 22316
rect 34412 23604 34468 23614
rect 34188 21980 34356 22036
rect 34076 21868 34244 21924
rect 34076 21476 34132 21486
rect 34076 21382 34132 21420
rect 33740 20468 33796 20478
rect 33740 19460 33796 20412
rect 33740 19404 34020 19460
rect 33628 18510 33630 18562
rect 33682 18510 33684 18562
rect 33628 18498 33684 18510
rect 33292 15986 33460 15988
rect 33292 15934 33294 15986
rect 33346 15934 33460 15986
rect 33292 15932 33460 15934
rect 33964 15986 34020 19404
rect 34188 16770 34244 21868
rect 34300 19906 34356 21980
rect 34300 19854 34302 19906
rect 34354 19854 34356 19906
rect 34300 19842 34356 19854
rect 34412 17554 34468 23548
rect 34636 21924 34692 23886
rect 34636 21858 34692 21868
rect 34524 21812 34580 21822
rect 34524 19122 34580 21756
rect 34524 19070 34526 19122
rect 34578 19070 34580 19122
rect 34524 19058 34580 19070
rect 34636 20802 34692 20814
rect 34636 20750 34638 20802
rect 34690 20750 34692 20802
rect 34636 18564 34692 20750
rect 34636 18498 34692 18508
rect 34748 18338 34804 24108
rect 34860 21812 34916 25228
rect 35084 25218 35140 25228
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 23940 35140 23950
rect 35084 23846 35140 23884
rect 35756 23938 35812 23950
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35532 23826 35588 23838
rect 35532 23774 35534 23826
rect 35586 23774 35588 23826
rect 34972 23156 35028 23166
rect 34972 23154 35140 23156
rect 34972 23102 34974 23154
rect 35026 23102 35140 23154
rect 34972 23100 35140 23102
rect 34972 23090 35028 23100
rect 34860 21746 34916 21756
rect 34972 22372 35028 22382
rect 34972 20802 35028 22316
rect 35084 22036 35140 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22148 35588 23774
rect 35756 23044 35812 23886
rect 35756 22978 35812 22988
rect 35532 22082 35588 22092
rect 35084 21980 35364 22036
rect 35308 21812 35364 21980
rect 35756 21924 35812 21934
rect 35308 21756 35588 21812
rect 35196 21700 35252 21710
rect 35196 21606 35252 21644
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34972 20750 34974 20802
rect 35026 20750 35028 20802
rect 34972 20738 35028 20750
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34748 18286 34750 18338
rect 34802 18286 34804 18338
rect 34748 18274 34804 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17780 35476 17790
rect 35532 17780 35588 21756
rect 35756 21700 35812 21868
rect 35420 17778 35588 17780
rect 35420 17726 35422 17778
rect 35474 17726 35588 17778
rect 35420 17724 35588 17726
rect 35644 21644 35812 21700
rect 35868 21700 35924 26852
rect 36876 26740 36932 26750
rect 36092 26290 36148 26302
rect 36092 26238 36094 26290
rect 36146 26238 36148 26290
rect 36092 23604 36148 26238
rect 36428 26292 36484 26302
rect 36764 26292 36820 26302
rect 36428 26290 36820 26292
rect 36428 26238 36430 26290
rect 36482 26238 36766 26290
rect 36818 26238 36820 26290
rect 36428 26236 36820 26238
rect 36428 25508 36484 26236
rect 36764 26226 36820 26236
rect 36428 23940 36484 25452
rect 36428 23874 36484 23884
rect 36092 23538 36148 23548
rect 36876 22372 36932 26684
rect 37100 23940 37156 23950
rect 37100 23846 37156 23884
rect 37100 23604 37156 23614
rect 36876 22316 37044 22372
rect 35420 17714 35476 17724
rect 34412 17502 34414 17554
rect 34466 17502 34468 17554
rect 34412 17490 34468 17502
rect 35308 16996 35364 17006
rect 35308 16902 35364 16940
rect 34188 16718 34190 16770
rect 34242 16718 34244 16770
rect 34188 16706 34244 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 16212 35364 16222
rect 35644 16212 35700 21644
rect 35868 21634 35924 21644
rect 35980 22146 36036 22158
rect 35980 22094 35982 22146
rect 36034 22094 36036 22146
rect 35756 21364 35812 21374
rect 35756 21270 35812 21308
rect 35980 20916 36036 22094
rect 36540 22148 36596 22158
rect 36876 22148 36932 22158
rect 36540 22146 36708 22148
rect 36540 22094 36542 22146
rect 36594 22094 36708 22146
rect 36540 22092 36708 22094
rect 36540 22082 36596 22092
rect 36540 21924 36596 21934
rect 36540 21810 36596 21868
rect 36540 21758 36542 21810
rect 36594 21758 36596 21810
rect 36540 21746 36596 21758
rect 35980 20850 36036 20860
rect 36652 20244 36708 22092
rect 36652 20178 36708 20188
rect 36764 22146 36932 22148
rect 36764 22094 36878 22146
rect 36930 22094 36932 22146
rect 36764 22092 36932 22094
rect 35308 16210 35700 16212
rect 35308 16158 35310 16210
rect 35362 16158 35700 16210
rect 35308 16156 35700 16158
rect 35756 18564 35812 18574
rect 35308 16146 35364 16156
rect 33964 15934 33966 15986
rect 34018 15934 34020 15986
rect 33292 15922 33348 15932
rect 33964 15922 34020 15934
rect 32060 15374 32062 15426
rect 32114 15374 32116 15426
rect 32060 15362 32116 15374
rect 35756 15202 35812 18508
rect 36764 15426 36820 22092
rect 36876 22082 36932 22092
rect 36988 21924 37044 22316
rect 36876 21868 37044 21924
rect 36876 19906 36932 21868
rect 36988 20916 37044 20926
rect 36988 20822 37044 20860
rect 36876 19854 36878 19906
rect 36930 19854 36932 19906
rect 36876 19842 36932 19854
rect 37100 18340 37156 23548
rect 37212 20132 37268 27244
rect 37324 25284 37380 27356
rect 37548 27076 37604 27086
rect 37548 27074 37716 27076
rect 37548 27022 37550 27074
rect 37602 27022 37716 27074
rect 37548 27020 37716 27022
rect 37548 27010 37604 27020
rect 37660 26908 37716 27020
rect 37660 26852 38388 26908
rect 37324 25218 37380 25228
rect 37436 26290 37492 26302
rect 37436 26238 37438 26290
rect 37490 26238 37492 26290
rect 37436 24276 37492 26238
rect 38108 25506 38164 25518
rect 38108 25454 38110 25506
rect 38162 25454 38164 25506
rect 37884 25396 37940 25406
rect 37436 24210 37492 24220
rect 37548 25394 37940 25396
rect 37548 25342 37886 25394
rect 37938 25342 37940 25394
rect 37548 25340 37940 25342
rect 37436 23940 37492 23950
rect 37324 23938 37492 23940
rect 37324 23886 37438 23938
rect 37490 23886 37492 23938
rect 37324 23884 37492 23886
rect 37324 23156 37380 23884
rect 37436 23874 37492 23884
rect 37436 23380 37492 23390
rect 37548 23380 37604 25340
rect 37884 25330 37940 25340
rect 37436 23378 37604 23380
rect 37436 23326 37438 23378
rect 37490 23326 37604 23378
rect 37436 23324 37604 23326
rect 37436 23314 37492 23324
rect 38108 23156 38164 25454
rect 37324 23100 37492 23156
rect 37324 22932 37380 22942
rect 37324 20914 37380 22876
rect 37324 20862 37326 20914
rect 37378 20862 37380 20914
rect 37324 20850 37380 20862
rect 37436 20468 37492 23100
rect 38108 23090 38164 23100
rect 37660 23044 37716 23054
rect 37660 22258 37716 22988
rect 38220 23042 38276 23054
rect 38220 22990 38222 23042
rect 38274 22990 38276 23042
rect 37660 22206 37662 22258
rect 37714 22206 37716 22258
rect 37660 22194 37716 22206
rect 37996 22930 38052 22942
rect 37996 22878 37998 22930
rect 38050 22878 38052 22930
rect 37996 20692 38052 22878
rect 38220 21924 38276 22990
rect 38220 21858 38276 21868
rect 37996 20626 38052 20636
rect 37436 20412 38164 20468
rect 37996 20244 38052 20254
rect 37884 20132 37940 20142
rect 37212 20130 37940 20132
rect 37212 20078 37886 20130
rect 37938 20078 37940 20130
rect 37212 20076 37940 20078
rect 37884 20066 37940 20076
rect 37324 18340 37380 18350
rect 37100 18338 37380 18340
rect 37100 18286 37326 18338
rect 37378 18286 37380 18338
rect 37100 18284 37380 18286
rect 37324 18274 37380 18284
rect 37996 15986 38052 20188
rect 38108 16770 38164 20412
rect 38332 19346 38388 26852
rect 38444 25844 38500 27580
rect 38556 27076 38612 29260
rect 38556 27010 38612 27020
rect 38780 28196 38836 28206
rect 38444 25778 38500 25788
rect 38444 25508 38500 25518
rect 38444 25414 38500 25452
rect 38444 23156 38500 23166
rect 38444 23062 38500 23100
rect 38332 19294 38334 19346
rect 38386 19294 38388 19346
rect 38332 19282 38388 19294
rect 38444 21812 38500 21822
rect 38444 18562 38500 21756
rect 38780 20916 38836 28140
rect 38892 28082 38948 29372
rect 40572 28868 40628 29934
rect 40572 28802 40628 28812
rect 40684 29428 40740 30156
rect 41132 30210 41300 30212
rect 41132 30158 41246 30210
rect 41298 30158 41300 30210
rect 41132 30156 41300 30158
rect 40908 29988 40964 29998
rect 40908 29538 40964 29932
rect 40908 29486 40910 29538
rect 40962 29486 40964 29538
rect 40908 29474 40964 29486
rect 40012 28642 40068 28654
rect 40012 28590 40014 28642
rect 40066 28590 40068 28642
rect 39900 28420 39956 28430
rect 38892 28030 38894 28082
rect 38946 28030 38948 28082
rect 38892 26908 38948 28030
rect 39452 28084 39508 28094
rect 39452 28082 39844 28084
rect 39452 28030 39454 28082
rect 39506 28030 39844 28082
rect 39452 28028 39844 28030
rect 39452 28018 39508 28028
rect 39676 27860 39732 27870
rect 39564 27804 39676 27860
rect 39564 27746 39620 27804
rect 39676 27794 39732 27804
rect 39564 27694 39566 27746
rect 39618 27694 39620 27746
rect 39564 27682 39620 27694
rect 39788 26962 39844 28028
rect 39900 27970 39956 28364
rect 39900 27918 39902 27970
rect 39954 27918 39956 27970
rect 39900 27906 39956 27918
rect 40012 27748 40068 28590
rect 40572 28644 40628 28654
rect 40684 28644 40740 29372
rect 40572 28642 41076 28644
rect 40572 28590 40574 28642
rect 40626 28590 41076 28642
rect 40572 28588 41076 28590
rect 40572 28578 40628 28588
rect 40684 28420 40740 28430
rect 40684 28418 40964 28420
rect 40684 28366 40686 28418
rect 40738 28366 40964 28418
rect 40684 28364 40964 28366
rect 40684 28354 40740 28364
rect 40236 27972 40292 27982
rect 40236 27878 40292 27916
rect 40012 27682 40068 27692
rect 40796 27634 40852 27646
rect 40796 27582 40798 27634
rect 40850 27582 40852 27634
rect 40684 27076 40740 27086
rect 40684 26982 40740 27020
rect 39788 26910 39790 26962
rect 39842 26910 39844 26962
rect 38892 26852 39172 26908
rect 39788 26898 39844 26910
rect 39004 25508 39060 25518
rect 38892 25506 39060 25508
rect 38892 25454 39006 25506
rect 39058 25454 39060 25506
rect 38892 25452 39060 25454
rect 38892 23716 38948 25452
rect 39004 25442 39060 25452
rect 39004 25284 39060 25294
rect 39004 24388 39060 25228
rect 39116 24722 39172 26852
rect 40572 26850 40628 26862
rect 40572 26798 40574 26850
rect 40626 26798 40628 26850
rect 39676 26402 39732 26414
rect 39676 26350 39678 26402
rect 39730 26350 39732 26402
rect 39564 25620 39620 25630
rect 39564 24834 39620 25564
rect 39676 24946 39732 26350
rect 40460 26066 40516 26078
rect 40460 26014 40462 26066
rect 40514 26014 40516 26066
rect 39676 24894 39678 24946
rect 39730 24894 39732 24946
rect 39676 24882 39732 24894
rect 39900 25844 39956 25854
rect 39564 24782 39566 24834
rect 39618 24782 39620 24834
rect 39564 24770 39620 24782
rect 39116 24670 39118 24722
rect 39170 24670 39172 24722
rect 39116 24612 39172 24670
rect 39116 24546 39172 24556
rect 39004 24332 39172 24388
rect 39004 23716 39060 23726
rect 38892 23660 39004 23716
rect 39004 23650 39060 23660
rect 38892 23156 38948 23166
rect 38892 23062 38948 23100
rect 38892 21588 38948 21598
rect 38892 21586 39060 21588
rect 38892 21534 38894 21586
rect 38946 21534 39060 21586
rect 38892 21532 39060 21534
rect 38892 21522 38948 21532
rect 38892 20916 38948 20926
rect 38780 20914 38948 20916
rect 38780 20862 38894 20914
rect 38946 20862 38948 20914
rect 38780 20860 38948 20862
rect 38892 20850 38948 20860
rect 38444 18510 38446 18562
rect 38498 18510 38500 18562
rect 38444 18498 38500 18510
rect 38892 20692 38948 20702
rect 38892 16994 38948 20636
rect 38892 16942 38894 16994
rect 38946 16942 38948 16994
rect 38892 16930 38948 16942
rect 38108 16718 38110 16770
rect 38162 16718 38164 16770
rect 38108 16706 38164 16718
rect 39004 16212 39060 21532
rect 39116 19124 39172 24332
rect 39788 23716 39844 23726
rect 39228 23714 39844 23716
rect 39228 23662 39790 23714
rect 39842 23662 39844 23714
rect 39228 23660 39844 23662
rect 39228 23266 39284 23660
rect 39788 23650 39844 23660
rect 39228 23214 39230 23266
rect 39282 23214 39284 23266
rect 39228 23202 39284 23214
rect 39564 23156 39620 23166
rect 39564 23062 39620 23100
rect 39788 23044 39844 23054
rect 39788 22950 39844 22988
rect 39452 21588 39508 21598
rect 39452 21494 39508 21532
rect 39788 21588 39844 21598
rect 39788 21494 39844 21532
rect 39900 20690 39956 25788
rect 40348 24612 40404 24622
rect 40348 24518 40404 24556
rect 40124 24276 40180 24286
rect 39900 20638 39902 20690
rect 39954 20638 39956 20690
rect 39900 20626 39956 20638
rect 40012 22370 40068 22382
rect 40012 22318 40014 22370
rect 40066 22318 40068 22370
rect 40012 20356 40068 22318
rect 40012 20290 40068 20300
rect 39340 19124 39396 19134
rect 39116 19122 39396 19124
rect 39116 19070 39342 19122
rect 39394 19070 39396 19122
rect 39116 19068 39396 19070
rect 39340 19058 39396 19068
rect 40124 17778 40180 24220
rect 40348 23828 40404 23838
rect 40348 23378 40404 23772
rect 40460 23604 40516 26014
rect 40572 24388 40628 26798
rect 40684 24388 40740 24398
rect 40572 24332 40684 24388
rect 40684 24322 40740 24332
rect 40796 24052 40852 27582
rect 40908 25060 40964 28364
rect 41020 26514 41076 28588
rect 41020 26462 41022 26514
rect 41074 26462 41076 26514
rect 41020 26450 41076 26462
rect 40908 24994 40964 25004
rect 41132 24948 41188 30156
rect 41244 30146 41300 30156
rect 43596 30212 43652 34638
rect 45164 34802 45220 34814
rect 45164 34750 45166 34802
rect 45218 34750 45220 34802
rect 43708 34242 43764 34254
rect 43708 34190 43710 34242
rect 43762 34190 43764 34242
rect 43708 32900 43764 34190
rect 44492 34020 44548 34030
rect 44716 34020 44772 34030
rect 44492 33926 44548 33964
rect 44604 34018 44772 34020
rect 44604 33966 44718 34018
rect 44770 33966 44772 34018
rect 44604 33964 44772 33966
rect 43932 33796 43988 33806
rect 43932 33460 43988 33740
rect 43932 33366 43988 33404
rect 44604 33348 44660 33964
rect 44716 33954 44772 33964
rect 45052 34018 45108 34030
rect 45052 33966 45054 34018
rect 45106 33966 45108 34018
rect 45052 33796 45108 33966
rect 45052 33730 45108 33740
rect 44380 33292 44660 33348
rect 44716 33346 44772 33358
rect 44716 33294 44718 33346
rect 44770 33294 44772 33346
rect 43820 33124 43876 33134
rect 43820 33030 43876 33068
rect 43708 32834 43764 32844
rect 44380 32786 44436 33292
rect 44380 32734 44382 32786
rect 44434 32734 44436 32786
rect 44380 32722 44436 32734
rect 44716 32452 44772 33294
rect 44940 32788 44996 32798
rect 44940 32694 44996 32732
rect 44156 31778 44212 31790
rect 44156 31726 44158 31778
rect 44210 31726 44212 31778
rect 43932 31666 43988 31678
rect 43932 31614 43934 31666
rect 43986 31614 43988 31666
rect 43708 31556 43764 31566
rect 43708 31218 43764 31500
rect 43708 31166 43710 31218
rect 43762 31166 43764 31218
rect 43708 31154 43764 31166
rect 43596 30146 43652 30156
rect 43596 29986 43652 29998
rect 43596 29934 43598 29986
rect 43650 29934 43652 29986
rect 41692 29764 41748 29774
rect 41580 29652 41636 29662
rect 41244 29596 41580 29652
rect 41244 29538 41300 29596
rect 41580 29586 41636 29596
rect 41244 29486 41246 29538
rect 41298 29486 41300 29538
rect 41244 29474 41300 29486
rect 41580 29314 41636 29326
rect 41580 29262 41582 29314
rect 41634 29262 41636 29314
rect 41468 28532 41524 28542
rect 41580 28532 41636 29262
rect 41468 28530 41636 28532
rect 41468 28478 41470 28530
rect 41522 28478 41636 28530
rect 41468 28476 41636 28478
rect 41468 28466 41524 28476
rect 41580 28084 41636 28094
rect 41692 28084 41748 29708
rect 41580 28082 41748 28084
rect 41580 28030 41582 28082
rect 41634 28030 41748 28082
rect 41580 28028 41748 28030
rect 41916 29652 41972 29662
rect 41916 29538 41972 29596
rect 41916 29486 41918 29538
rect 41970 29486 41972 29538
rect 41580 28018 41636 28028
rect 41916 27972 41972 29486
rect 42252 29428 42308 29438
rect 42252 29334 42308 29372
rect 42924 29426 42980 29438
rect 42924 29374 42926 29426
rect 42978 29374 42980 29426
rect 41468 27748 41524 27758
rect 41356 27076 41412 27086
rect 41356 26982 41412 27020
rect 41356 26292 41412 26302
rect 41132 24882 41188 24892
rect 41244 26290 41412 26292
rect 41244 26238 41358 26290
rect 41410 26238 41412 26290
rect 41244 26236 41412 26238
rect 41020 24724 41076 24734
rect 41244 24724 41300 26236
rect 41356 26226 41412 26236
rect 41020 24722 41300 24724
rect 41020 24670 41022 24722
rect 41074 24670 41300 24722
rect 41020 24668 41300 24670
rect 41356 24722 41412 24734
rect 41356 24670 41358 24722
rect 41410 24670 41412 24722
rect 40796 23996 40964 24052
rect 40684 23938 40740 23950
rect 40684 23886 40686 23938
rect 40738 23886 40740 23938
rect 40684 23828 40740 23886
rect 40796 23828 40852 23838
rect 40684 23772 40796 23828
rect 40796 23762 40852 23772
rect 40460 23538 40516 23548
rect 40572 23714 40628 23726
rect 40572 23662 40574 23714
rect 40626 23662 40628 23714
rect 40348 23326 40350 23378
rect 40402 23326 40404 23378
rect 40348 22370 40404 23326
rect 40572 22596 40628 23662
rect 40908 23156 40964 23996
rect 40572 22530 40628 22540
rect 40796 23100 40964 23156
rect 41020 23828 41076 24668
rect 40348 22318 40350 22370
rect 40402 22318 40404 22370
rect 40348 22306 40404 22318
rect 40796 19124 40852 23100
rect 41020 23042 41076 23772
rect 41020 22990 41022 23042
rect 41074 22990 41076 23042
rect 40908 22372 40964 22382
rect 41020 22372 41076 22990
rect 40908 22370 41076 22372
rect 40908 22318 40910 22370
rect 40962 22318 41076 22370
rect 40908 22316 41076 22318
rect 40908 22306 40964 22316
rect 41020 21588 41076 22316
rect 41020 21474 41076 21532
rect 41020 21422 41022 21474
rect 41074 21422 41076 21474
rect 41020 20244 41076 21422
rect 41020 20178 41076 20188
rect 41132 24388 41188 24398
rect 40796 19058 40852 19068
rect 40124 17726 40126 17778
rect 40178 17726 40180 17778
rect 40124 17714 40180 17726
rect 41132 17554 41188 24332
rect 41244 23938 41300 23950
rect 41244 23886 41246 23938
rect 41298 23886 41300 23938
rect 41244 19012 41300 23886
rect 41356 22820 41412 24670
rect 41356 22754 41412 22764
rect 41244 18946 41300 18956
rect 41356 22370 41412 22382
rect 41356 22318 41358 22370
rect 41410 22318 41412 22370
rect 41356 18452 41412 22318
rect 41468 19348 41524 27692
rect 41916 25620 41972 27916
rect 42028 26292 42084 26302
rect 42028 26290 42532 26292
rect 42028 26238 42030 26290
rect 42082 26238 42532 26290
rect 42028 26236 42532 26238
rect 42028 26226 42084 26236
rect 41916 25554 41972 25564
rect 41580 25396 41636 25406
rect 41580 25282 41636 25340
rect 42364 25396 42420 25406
rect 42364 25302 42420 25340
rect 41580 25230 41582 25282
rect 41634 25230 41636 25282
rect 41580 25218 41636 25230
rect 42140 25284 42196 25294
rect 42140 25282 42308 25284
rect 42140 25230 42142 25282
rect 42194 25230 42308 25282
rect 42140 25228 42308 25230
rect 42140 25218 42196 25228
rect 42140 24948 42196 24958
rect 41692 24612 41748 24622
rect 41580 23716 41636 23726
rect 41580 22708 41636 23660
rect 41692 23156 41748 24556
rect 42028 23156 42084 23166
rect 41692 23154 42084 23156
rect 41692 23102 41694 23154
rect 41746 23102 42030 23154
rect 42082 23102 42084 23154
rect 41692 23100 42084 23102
rect 41692 23090 41748 23100
rect 42028 23090 42084 23100
rect 41580 22652 41972 22708
rect 41580 21364 41636 21374
rect 41580 21362 41748 21364
rect 41580 21310 41582 21362
rect 41634 21310 41748 21362
rect 41580 21308 41748 21310
rect 41580 21298 41636 21308
rect 41580 19348 41636 19358
rect 41468 19346 41636 19348
rect 41468 19294 41582 19346
rect 41634 19294 41636 19346
rect 41468 19292 41636 19294
rect 41580 19282 41636 19292
rect 41356 18386 41412 18396
rect 41132 17502 41134 17554
rect 41186 17502 41188 17554
rect 41132 17490 41188 17502
rect 39116 16212 39172 16222
rect 39004 16210 39172 16212
rect 39004 16158 39118 16210
rect 39170 16158 39172 16210
rect 39004 16156 39172 16158
rect 39116 16146 39172 16156
rect 37996 15934 37998 15986
rect 38050 15934 38052 15986
rect 37996 15922 38052 15934
rect 41692 15988 41748 21308
rect 41804 20356 41860 20366
rect 41804 16772 41860 20300
rect 41916 18338 41972 22652
rect 42140 20914 42196 24892
rect 42252 21588 42308 25228
rect 42364 24612 42420 24622
rect 42364 21810 42420 24556
rect 42364 21758 42366 21810
rect 42418 21758 42420 21810
rect 42364 21746 42420 21758
rect 42252 21522 42308 21532
rect 42476 21476 42532 26236
rect 42700 25620 42756 25630
rect 42700 25526 42756 25564
rect 42924 24052 42980 29374
rect 43596 26908 43652 29934
rect 43932 29764 43988 31614
rect 43932 29698 43988 29708
rect 44156 29652 44212 31726
rect 44716 31778 44772 32396
rect 44716 31726 44718 31778
rect 44770 31726 44772 31778
rect 44716 30994 44772 31726
rect 45164 31556 45220 34750
rect 45500 34804 45556 34814
rect 46060 34804 46116 34862
rect 45500 34802 46116 34804
rect 45500 34750 45502 34802
rect 45554 34750 46116 34802
rect 45500 34748 46116 34750
rect 45500 34738 45556 34748
rect 45612 34130 45668 34142
rect 45612 34078 45614 34130
rect 45666 34078 45668 34130
rect 45388 33348 45444 33358
rect 45388 33254 45444 33292
rect 45388 32564 45444 32574
rect 45388 32228 45444 32508
rect 45388 32162 45444 32172
rect 45612 32564 45668 34078
rect 46060 33796 46116 34748
rect 46060 33730 46116 33740
rect 46284 34802 46340 34814
rect 46284 34750 46286 34802
rect 46338 34750 46340 34802
rect 46284 33236 46340 34750
rect 46284 33170 46340 33180
rect 46396 32788 46452 36540
rect 46732 35028 46788 37100
rect 47068 36484 47124 36494
rect 47068 36390 47124 36428
rect 47740 35922 47796 38670
rect 47852 37492 47908 39342
rect 48748 39396 48804 39406
rect 48748 39394 48916 39396
rect 48748 39342 48750 39394
rect 48802 39342 48916 39394
rect 48748 39340 48916 39342
rect 48748 39330 48804 39340
rect 47852 37426 47908 37436
rect 47964 38722 48020 38734
rect 48748 38724 48804 38734
rect 47964 38670 47966 38722
rect 48018 38670 48020 38722
rect 47964 38668 48020 38670
rect 48636 38722 48804 38724
rect 48636 38670 48750 38722
rect 48802 38670 48804 38722
rect 48636 38668 48804 38670
rect 47964 38612 48692 38668
rect 48748 38658 48804 38668
rect 47964 37380 48020 38612
rect 48748 38052 48804 38062
rect 48860 38052 48916 39340
rect 49532 38834 49588 39676
rect 49532 38782 49534 38834
rect 49586 38782 49588 38834
rect 48972 38724 49028 38734
rect 48972 38630 49028 38668
rect 47964 37314 48020 37324
rect 48188 38050 48916 38052
rect 48188 37998 48750 38050
rect 48802 37998 48916 38050
rect 48188 37996 48916 37998
rect 48188 37490 48244 37996
rect 48748 37986 48804 37996
rect 48412 37828 48468 37838
rect 48412 37734 48468 37772
rect 48188 37438 48190 37490
rect 48242 37438 48244 37490
rect 48188 37156 48244 37438
rect 48524 37380 48580 37390
rect 48748 37380 48804 37390
rect 48580 37378 48804 37380
rect 48580 37326 48750 37378
rect 48802 37326 48804 37378
rect 48580 37324 48804 37326
rect 48524 37314 48580 37324
rect 48748 37314 48804 37324
rect 48860 37380 48916 37996
rect 49196 38388 49252 38398
rect 49196 38050 49252 38332
rect 49196 37998 49198 38050
rect 49250 37998 49252 38050
rect 49196 37986 49252 37998
rect 49532 37604 49588 38782
rect 49644 39730 49700 39742
rect 49644 39678 49646 39730
rect 49698 39678 49700 39730
rect 49644 38500 49700 39678
rect 50204 38834 50260 40012
rect 51436 39730 51492 40124
rect 51436 39678 51438 39730
rect 51490 39678 51492 39730
rect 51436 39666 51492 39678
rect 51772 39730 51828 40348
rect 51996 40338 52052 40348
rect 52444 41188 52500 41918
rect 52556 41188 52612 41198
rect 52444 41186 52612 41188
rect 52444 41134 52558 41186
rect 52610 41134 52612 41186
rect 52444 41132 52612 41134
rect 52444 40402 52500 41132
rect 52556 41122 52612 41132
rect 52444 40350 52446 40402
rect 52498 40350 52500 40402
rect 52220 40292 52276 40302
rect 52220 40290 52388 40292
rect 52220 40238 52222 40290
rect 52274 40238 52388 40290
rect 52220 40236 52388 40238
rect 52220 40226 52276 40236
rect 51772 39678 51774 39730
rect 51826 39678 51828 39730
rect 51772 39666 51828 39678
rect 50876 39506 50932 39518
rect 50876 39454 50878 39506
rect 50930 39454 50932 39506
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50204 38782 50206 38834
rect 50258 38782 50260 38834
rect 50204 38770 50260 38782
rect 49644 38434 49700 38444
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 49532 37548 50036 37604
rect 50556 37594 50820 37604
rect 48188 37090 48244 37100
rect 48412 37044 48468 37054
rect 48076 36484 48132 36494
rect 48300 36484 48356 36494
rect 48132 36482 48356 36484
rect 48132 36430 48302 36482
rect 48354 36430 48356 36482
rect 48132 36428 48356 36430
rect 48076 36390 48132 36428
rect 48300 36418 48356 36428
rect 47740 35870 47742 35922
rect 47794 35870 47796 35922
rect 47740 35858 47796 35870
rect 48300 35924 48356 35934
rect 48412 35924 48468 36988
rect 48300 35922 48468 35924
rect 48300 35870 48302 35922
rect 48354 35870 48468 35922
rect 48300 35868 48468 35870
rect 48860 35924 48916 37324
rect 48972 37492 49028 37502
rect 48972 37154 49028 37436
rect 49532 37380 49588 37390
rect 49532 37286 49588 37324
rect 49980 37268 50036 37548
rect 49980 37266 50372 37268
rect 49980 37214 49982 37266
rect 50034 37214 50372 37266
rect 49980 37212 50372 37214
rect 49980 37202 50036 37212
rect 48972 37102 48974 37154
rect 49026 37102 49028 37154
rect 48972 37090 49028 37102
rect 50316 36932 50372 37212
rect 50652 37266 50708 37278
rect 50652 37214 50654 37266
rect 50706 37214 50708 37266
rect 50652 37156 50708 37214
rect 50652 37090 50708 37100
rect 50316 36876 50484 36932
rect 50316 36594 50372 36606
rect 50316 36542 50318 36594
rect 50370 36542 50372 36594
rect 49308 35924 49364 35934
rect 48860 35922 49364 35924
rect 48860 35870 48862 35922
rect 48914 35870 49310 35922
rect 49362 35870 49364 35922
rect 48860 35868 49364 35870
rect 48300 35858 48356 35868
rect 48860 35858 48916 35868
rect 49308 35858 49364 35868
rect 50316 35810 50372 36542
rect 50316 35758 50318 35810
rect 50370 35758 50372 35810
rect 47628 35588 47684 35598
rect 46732 35026 47012 35028
rect 46732 34974 46734 35026
rect 46786 34974 47012 35026
rect 46732 34972 47012 34974
rect 46732 34962 46788 34972
rect 46956 34914 47012 34972
rect 46956 34862 46958 34914
rect 47010 34862 47012 34914
rect 46956 34850 47012 34862
rect 47628 34914 47684 35532
rect 47628 34862 47630 34914
rect 47682 34862 47684 34914
rect 47628 34850 47684 34862
rect 49980 35586 50036 35598
rect 49980 35534 49982 35586
rect 50034 35534 50036 35586
rect 49980 34690 50036 35534
rect 50316 35588 50372 35758
rect 50428 36484 50484 36876
rect 50876 36708 50932 39454
rect 52332 39060 52388 40236
rect 52444 39732 52500 40350
rect 52444 39666 52500 39676
rect 52668 39396 52724 44270
rect 52780 43764 52836 45836
rect 52892 45108 52948 47516
rect 53004 47460 53060 48972
rect 53116 48244 53172 48254
rect 53452 48244 53508 48254
rect 53116 48242 53452 48244
rect 53116 48190 53118 48242
rect 53170 48190 53452 48242
rect 53116 48188 53452 48190
rect 53116 48018 53172 48188
rect 53452 48178 53508 48188
rect 53564 48132 53620 48142
rect 53564 48038 53620 48076
rect 53116 47966 53118 48018
rect 53170 47966 53172 48018
rect 53116 47954 53172 47966
rect 53228 48020 53284 48030
rect 53116 47460 53172 47470
rect 53004 47458 53172 47460
rect 53004 47406 53118 47458
rect 53170 47406 53172 47458
rect 53004 47404 53172 47406
rect 53116 47394 53172 47404
rect 53228 47236 53284 47964
rect 54012 48020 54068 50654
rect 56812 50706 56868 50718
rect 56812 50654 56814 50706
rect 56866 50654 56868 50706
rect 55132 50482 55188 50494
rect 55132 50430 55134 50482
rect 55186 50430 55188 50482
rect 54124 49924 54180 49934
rect 54124 49830 54180 49868
rect 54348 49810 54404 49822
rect 54348 49758 54350 49810
rect 54402 49758 54404 49810
rect 54348 49588 54404 49758
rect 54348 49522 54404 49532
rect 55020 49698 55076 49710
rect 55020 49646 55022 49698
rect 55074 49646 55076 49698
rect 55020 49588 55076 49646
rect 55020 49522 55076 49532
rect 54684 48916 54740 48926
rect 54684 48822 54740 48860
rect 54012 47954 54068 47964
rect 54572 48354 54628 48366
rect 54572 48302 54574 48354
rect 54626 48302 54628 48354
rect 53116 47180 53284 47236
rect 53116 45890 53172 47180
rect 53228 46788 53284 46798
rect 53228 46694 53284 46732
rect 54572 46228 54628 48302
rect 55132 47908 55188 50430
rect 56252 49924 56308 49934
rect 55468 49698 55524 49710
rect 55468 49646 55470 49698
rect 55522 49646 55524 49698
rect 55356 49588 55412 49598
rect 55356 49250 55412 49532
rect 55356 49198 55358 49250
rect 55410 49198 55412 49250
rect 55356 48354 55412 49198
rect 55356 48302 55358 48354
rect 55410 48302 55412 48354
rect 55356 48290 55412 48302
rect 55468 48244 55524 49646
rect 55580 49250 55636 49262
rect 55580 49198 55582 49250
rect 55634 49198 55636 49250
rect 55580 49138 55636 49198
rect 55580 49086 55582 49138
rect 55634 49086 55636 49138
rect 55580 49074 55636 49086
rect 55468 48178 55524 48188
rect 55692 48356 55748 48366
rect 55132 47842 55188 47852
rect 55580 48130 55636 48142
rect 55580 48078 55582 48130
rect 55634 48078 55636 48130
rect 55580 47234 55636 48078
rect 55580 47182 55582 47234
rect 55634 47182 55636 47234
rect 55580 47170 55636 47182
rect 55580 46676 55636 46686
rect 55692 46676 55748 48300
rect 56252 47682 56308 49868
rect 56476 49476 56532 49486
rect 56476 49138 56532 49420
rect 56476 49086 56478 49138
rect 56530 49086 56532 49138
rect 56476 49074 56532 49086
rect 56812 49028 56868 50654
rect 57820 50484 57876 50494
rect 57820 50390 57876 50428
rect 58828 49924 58884 49934
rect 58828 49830 58884 49868
rect 56812 48962 56868 48972
rect 57596 49698 57652 49710
rect 57596 49646 57598 49698
rect 57650 49646 57652 49698
rect 57484 48916 57540 48926
rect 57484 48822 57540 48860
rect 57596 48356 57652 49646
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 57596 48290 57652 48300
rect 58828 48354 58884 48366
rect 58828 48302 58830 48354
rect 58882 48302 58884 48354
rect 57596 48130 57652 48142
rect 57596 48078 57598 48130
rect 57650 48078 57652 48130
rect 57596 47796 57652 48078
rect 57596 47730 57652 47740
rect 56252 47630 56254 47682
rect 56306 47630 56308 47682
rect 56252 47618 56308 47630
rect 57484 47572 57540 47582
rect 57484 47478 57540 47516
rect 56140 47348 56196 47358
rect 55580 46674 55748 46676
rect 55580 46622 55582 46674
rect 55634 46622 55748 46674
rect 55580 46620 55748 46622
rect 56028 47292 56140 47348
rect 55580 46610 55636 46620
rect 54572 46162 54628 46172
rect 53116 45838 53118 45890
rect 53170 45838 53172 45890
rect 53116 45826 53172 45838
rect 55692 45892 55748 45902
rect 55692 45666 55748 45836
rect 55692 45614 55694 45666
rect 55746 45614 55748 45666
rect 55692 45602 55748 45614
rect 53116 45332 53172 45342
rect 56028 45332 56084 47292
rect 56140 47282 56196 47292
rect 58492 47348 58548 47358
rect 58492 47254 58548 47292
rect 56588 47236 56644 47246
rect 56588 47234 56756 47236
rect 56588 47182 56590 47234
rect 56642 47182 56756 47234
rect 56588 47180 56756 47182
rect 56588 47170 56644 47180
rect 56252 47124 56308 47134
rect 56140 46674 56196 46686
rect 56140 46622 56142 46674
rect 56194 46622 56196 46674
rect 56140 45668 56196 46622
rect 56252 46114 56308 47068
rect 56252 46062 56254 46114
rect 56306 46062 56308 46114
rect 56252 46050 56308 46062
rect 56700 46562 56756 47180
rect 58828 47124 58884 48302
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 59388 47236 59444 47246
rect 59388 47234 59556 47236
rect 59388 47182 59390 47234
rect 59442 47182 59556 47234
rect 59388 47180 59556 47182
rect 59388 47170 59444 47180
rect 58828 47058 58884 47068
rect 58828 46788 58884 46798
rect 58828 46694 58884 46732
rect 59388 46788 59444 46798
rect 59388 46694 59444 46732
rect 59500 46676 59556 47180
rect 59612 46676 59668 46686
rect 59500 46674 59668 46676
rect 59500 46622 59614 46674
rect 59666 46622 59668 46674
rect 59500 46620 59668 46622
rect 56700 46510 56702 46562
rect 56754 46510 56756 46562
rect 56588 45668 56644 45678
rect 56700 45668 56756 46510
rect 57148 46562 57204 46574
rect 57148 46510 57150 46562
rect 57202 46510 57204 46562
rect 57036 45668 57092 45678
rect 57148 45668 57204 46510
rect 57596 46562 57652 46574
rect 57596 46510 57598 46562
rect 57650 46510 57652 46562
rect 57484 46004 57540 46014
rect 57484 45910 57540 45948
rect 56140 45666 57204 45668
rect 56140 45614 56590 45666
rect 56642 45614 57038 45666
rect 57090 45614 57204 45666
rect 56140 45612 57204 45614
rect 56588 45602 56644 45612
rect 57036 45602 57092 45612
rect 56140 45332 56196 45342
rect 56028 45330 56196 45332
rect 56028 45278 56142 45330
rect 56194 45278 56196 45330
rect 56028 45276 56196 45278
rect 53004 45108 53060 45118
rect 52892 45106 53060 45108
rect 52892 45054 53006 45106
rect 53058 45054 53060 45106
rect 52892 45052 53060 45054
rect 53004 45042 53060 45052
rect 52780 43540 52836 43708
rect 52780 42754 52836 43484
rect 52780 42702 52782 42754
rect 52834 42702 52836 42754
rect 52780 42690 52836 42702
rect 53004 44436 53060 44446
rect 53004 41970 53060 44380
rect 53116 42754 53172 45276
rect 56140 45266 56196 45276
rect 55356 45220 55412 45230
rect 55356 45126 55412 45164
rect 56700 44996 56756 45006
rect 56700 44902 56756 44940
rect 57148 44994 57204 45612
rect 57596 45332 57652 46510
rect 59276 45892 59332 45902
rect 59276 45798 59332 45836
rect 59500 45890 59556 46620
rect 59612 46610 59668 46620
rect 59500 45838 59502 45890
rect 59554 45838 59556 45890
rect 58492 45780 58548 45790
rect 58492 45686 58548 45724
rect 57596 45266 57652 45276
rect 59500 45668 59556 45838
rect 61404 46452 61460 46462
rect 58828 45218 58884 45230
rect 58828 45166 58830 45218
rect 58882 45166 58884 45218
rect 57148 44942 57150 44994
rect 57202 44942 57204 44994
rect 54124 44772 54180 44782
rect 54124 43538 54180 44716
rect 57148 44436 57204 44942
rect 56700 44434 57204 44436
rect 56700 44382 57150 44434
rect 57202 44382 57204 44434
rect 56700 44380 57204 44382
rect 55468 44212 55524 44222
rect 54908 43652 54964 43662
rect 54908 43558 54964 43596
rect 54124 43486 54126 43538
rect 54178 43486 54180 43538
rect 54124 43474 54180 43486
rect 54684 43540 54740 43550
rect 54684 43446 54740 43484
rect 55132 43538 55188 43550
rect 55132 43486 55134 43538
rect 55186 43486 55188 43538
rect 55132 43428 55188 43486
rect 55132 43362 55188 43372
rect 53116 42702 53118 42754
rect 53170 42702 53172 42754
rect 53116 42690 53172 42702
rect 53228 43316 53284 43326
rect 53004 41918 53006 41970
rect 53058 41918 53060 41970
rect 53004 41906 53060 41918
rect 53228 41186 53284 43260
rect 55468 42642 55524 44156
rect 56028 43764 56084 43774
rect 55916 43652 56084 43708
rect 56140 43652 56196 43662
rect 55916 43538 55972 43652
rect 55916 43486 55918 43538
rect 55970 43486 55972 43538
rect 55916 43474 55972 43486
rect 55468 42590 55470 42642
rect 55522 42590 55524 42642
rect 55468 42578 55524 42590
rect 55692 43426 55748 43438
rect 55692 43374 55694 43426
rect 55746 43374 55748 43426
rect 55356 42196 55412 42206
rect 55356 42102 55412 42140
rect 53228 41134 53230 41186
rect 53282 41134 53284 41186
rect 53228 41122 53284 41134
rect 55580 41300 55636 41310
rect 55356 40516 55412 40526
rect 54908 40514 55412 40516
rect 54908 40462 55358 40514
rect 55410 40462 55412 40514
rect 54908 40460 55412 40462
rect 53116 40404 53172 40414
rect 53116 40310 53172 40348
rect 53676 40180 53732 40190
rect 53004 39732 53060 39742
rect 53004 39618 53060 39676
rect 53004 39566 53006 39618
rect 53058 39566 53060 39618
rect 53004 39554 53060 39566
rect 53676 39618 53732 40124
rect 53676 39566 53678 39618
rect 53730 39566 53732 39618
rect 53676 39554 53732 39566
rect 53788 39732 53844 39742
rect 52780 39396 52836 39406
rect 52668 39394 52836 39396
rect 52668 39342 52782 39394
rect 52834 39342 52836 39394
rect 52668 39340 52836 39342
rect 52444 39060 52500 39070
rect 52332 39058 52500 39060
rect 52332 39006 52446 39058
rect 52498 39006 52500 39058
rect 52332 39004 52500 39006
rect 52444 38994 52500 39004
rect 52780 38052 52836 39340
rect 53788 39058 53844 39676
rect 53788 39006 53790 39058
rect 53842 39006 53844 39058
rect 53228 38948 53284 38958
rect 53228 38854 53284 38892
rect 53788 38836 53844 39006
rect 53788 38770 53844 38780
rect 54460 38724 54516 38734
rect 54348 38722 54516 38724
rect 54348 38670 54462 38722
rect 54514 38670 54516 38722
rect 54348 38668 54516 38670
rect 52780 37958 52836 37996
rect 53340 38164 53396 38174
rect 50876 36642 50932 36652
rect 51436 37826 51492 37838
rect 51436 37774 51438 37826
rect 51490 37774 51492 37826
rect 51436 36594 51492 37774
rect 52220 37828 52276 37838
rect 52220 37734 52276 37772
rect 53116 37490 53172 37502
rect 53116 37438 53118 37490
rect 53170 37438 53172 37490
rect 53116 37380 53172 37438
rect 53116 37314 53172 37324
rect 51436 36542 51438 36594
rect 51490 36542 51492 36594
rect 51436 36530 51492 36542
rect 53228 36596 53284 36606
rect 50428 35700 50484 36428
rect 51324 36482 51380 36494
rect 51324 36430 51326 36482
rect 51378 36430 51380 36482
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50540 35700 50596 35710
rect 50428 35698 50596 35700
rect 50428 35646 50542 35698
rect 50594 35646 50596 35698
rect 50428 35644 50596 35646
rect 50540 35634 50596 35644
rect 51100 35698 51156 35710
rect 51100 35646 51102 35698
rect 51154 35646 51156 35698
rect 50316 35532 50484 35588
rect 50428 35252 50484 35532
rect 50428 35186 50484 35196
rect 50988 35252 51044 35262
rect 50988 34914 51044 35196
rect 50988 34862 50990 34914
rect 51042 34862 51044 34914
rect 50988 34850 51044 34862
rect 49980 34638 49982 34690
rect 50034 34638 50036 34690
rect 49980 34626 50036 34638
rect 50652 34692 50708 34730
rect 50652 34626 50708 34636
rect 50556 34524 50820 34534
rect 48748 34468 48804 34478
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 47068 33908 47124 33918
rect 47068 33572 47124 33852
rect 47964 33906 48020 33918
rect 47964 33854 47966 33906
rect 48018 33854 48020 33906
rect 47964 33796 48020 33854
rect 47964 33730 48020 33740
rect 47068 33506 47124 33516
rect 48524 33346 48580 33358
rect 48524 33294 48526 33346
rect 48578 33294 48580 33346
rect 47628 33236 47684 33246
rect 47628 33142 47684 33180
rect 48412 33122 48468 33134
rect 48412 33070 48414 33122
rect 48466 33070 48468 33122
rect 46396 32722 46452 32732
rect 47180 33012 47236 33022
rect 47180 32674 47236 32956
rect 48412 32788 48468 33070
rect 48412 32722 48468 32732
rect 47180 32622 47182 32674
rect 47234 32622 47236 32674
rect 47180 32610 47236 32622
rect 45388 31778 45444 31790
rect 45388 31726 45390 31778
rect 45442 31726 45444 31778
rect 45164 31500 45332 31556
rect 44716 30942 44718 30994
rect 44770 30942 44772 30994
rect 44492 30772 44548 30782
rect 44492 30678 44548 30716
rect 44156 29586 44212 29596
rect 44380 29986 44436 29998
rect 44380 29934 44382 29986
rect 44434 29934 44436 29986
rect 44156 29428 44212 29438
rect 43372 26852 43652 26908
rect 43708 28642 43764 28654
rect 43708 28590 43710 28642
rect 43762 28590 43764 28642
rect 43148 25620 43204 25630
rect 43148 25506 43204 25564
rect 43372 25618 43428 26852
rect 43372 25566 43374 25618
rect 43426 25566 43428 25618
rect 43372 25554 43428 25566
rect 43148 25454 43150 25506
rect 43202 25454 43204 25506
rect 43148 25442 43204 25454
rect 42924 23986 42980 23996
rect 43148 25060 43204 25070
rect 42700 23604 42756 23614
rect 42588 21476 42644 21486
rect 42476 21420 42588 21476
rect 42588 21410 42644 21420
rect 42140 20862 42142 20914
rect 42194 20862 42196 20914
rect 42140 20850 42196 20862
rect 42364 20244 42420 20254
rect 42700 20244 42756 23548
rect 42924 22596 42980 22606
rect 42980 22540 43092 22596
rect 42924 22530 42980 22540
rect 42700 20188 42980 20244
rect 42364 20018 42420 20188
rect 42364 19966 42366 20018
rect 42418 19966 42420 20018
rect 42364 19348 42420 19966
rect 42364 19282 42420 19292
rect 42812 20018 42868 20030
rect 42812 19966 42814 20018
rect 42866 19966 42868 20018
rect 42588 19124 42644 19134
rect 42588 19030 42644 19068
rect 41916 18286 41918 18338
rect 41970 18286 41972 18338
rect 41916 18274 41972 18286
rect 42588 18452 42644 18462
rect 41916 16772 41972 16782
rect 41804 16770 41972 16772
rect 41804 16718 41918 16770
rect 41970 16718 41972 16770
rect 41804 16716 41972 16718
rect 41916 16706 41972 16716
rect 42588 16210 42644 18396
rect 42812 18116 42868 19966
rect 42924 18562 42980 20188
rect 42924 18510 42926 18562
rect 42978 18510 42980 18562
rect 42924 18498 42980 18510
rect 42812 18050 42868 18060
rect 43036 16994 43092 22540
rect 43148 20690 43204 25004
rect 43708 24164 43764 28590
rect 44156 28642 44212 29372
rect 44156 28590 44158 28642
rect 44210 28590 44212 28642
rect 43932 27858 43988 27870
rect 43932 27806 43934 27858
rect 43986 27806 43988 27858
rect 43932 27300 43988 27806
rect 44156 27860 44212 28590
rect 44380 28420 44436 29934
rect 44380 28354 44436 28364
rect 44716 29652 44772 30942
rect 45164 30994 45220 31006
rect 45164 30942 45166 30994
rect 45218 30942 45220 30994
rect 45164 30660 45220 30942
rect 45164 30594 45220 30604
rect 44716 28644 44772 29596
rect 45276 29650 45332 31500
rect 45276 29598 45278 29650
rect 45330 29598 45332 29650
rect 45276 29586 45332 29598
rect 45388 29540 45444 31726
rect 45612 31332 45668 32508
rect 48076 32564 48132 32574
rect 45724 32452 45780 32462
rect 45724 32358 45780 32396
rect 46172 32450 46228 32462
rect 46172 32398 46174 32450
rect 46226 32398 46228 32450
rect 46172 32340 46228 32398
rect 46172 32274 46228 32284
rect 47068 32340 47124 32350
rect 47068 31780 47124 32284
rect 47068 31714 47124 31724
rect 47852 31556 47908 31566
rect 47852 31462 47908 31500
rect 45612 31266 45668 31276
rect 47740 31218 47796 31230
rect 47740 31166 47742 31218
rect 47794 31166 47796 31218
rect 45388 29474 45444 29484
rect 46060 30772 46116 30782
rect 45948 29204 46004 29214
rect 45948 29110 46004 29148
rect 45612 28868 45668 28878
rect 44828 28644 44884 28654
rect 44716 28642 44884 28644
rect 44716 28590 44830 28642
rect 44882 28590 44884 28642
rect 44716 28588 44884 28590
rect 44268 27860 44324 27870
rect 44716 27860 44772 28588
rect 44828 28578 44884 28588
rect 45500 28644 45556 28654
rect 45500 28550 45556 28588
rect 44156 27858 44772 27860
rect 44156 27806 44270 27858
rect 44322 27806 44772 27858
rect 44156 27804 44772 27806
rect 44268 27794 44324 27804
rect 43932 27234 43988 27244
rect 44156 27076 44212 27086
rect 43820 26850 43876 26862
rect 43820 26798 43822 26850
rect 43874 26798 43876 26850
rect 43820 25618 43876 26798
rect 43820 25566 43822 25618
rect 43874 25566 43876 25618
rect 43820 25554 43876 25566
rect 44044 26068 44100 26078
rect 44044 25620 44100 26012
rect 44044 25526 44100 25564
rect 43708 24098 43764 24108
rect 43932 24946 43988 24958
rect 43932 24894 43934 24946
rect 43986 24894 43988 24946
rect 43820 23714 43876 23726
rect 43820 23662 43822 23714
rect 43874 23662 43876 23714
rect 43148 20638 43150 20690
rect 43202 20638 43204 20690
rect 43148 20626 43204 20638
rect 43596 22146 43652 22158
rect 43596 22094 43598 22146
rect 43650 22094 43652 22146
rect 43596 19010 43652 22094
rect 43820 20916 43876 23662
rect 43932 22260 43988 24894
rect 43932 22194 43988 22204
rect 43932 20916 43988 20926
rect 43820 20914 43988 20916
rect 43820 20862 43934 20914
rect 43986 20862 43988 20914
rect 43820 20860 43988 20862
rect 43932 20850 43988 20860
rect 43708 19684 43764 19694
rect 43708 19346 43764 19628
rect 43708 19294 43710 19346
rect 43762 19294 43764 19346
rect 43708 19282 43764 19294
rect 43596 18958 43598 19010
rect 43650 18958 43652 19010
rect 43596 18946 43652 18958
rect 44156 18340 44212 27020
rect 44716 27074 44772 27804
rect 44828 27860 44884 27870
rect 44828 27766 44884 27804
rect 45276 27860 45332 27870
rect 45276 27858 45556 27860
rect 45276 27806 45278 27858
rect 45330 27806 45556 27858
rect 45276 27804 45556 27806
rect 45276 27794 45332 27804
rect 44716 27022 44718 27074
rect 44770 27022 44772 27074
rect 44716 26908 44772 27022
rect 45388 27076 45444 27086
rect 45388 26982 45444 27020
rect 44380 26852 44436 26862
rect 44716 26852 44996 26908
rect 44268 26850 44436 26852
rect 44268 26798 44382 26850
rect 44434 26798 44436 26850
rect 44268 26796 44436 26798
rect 44268 21924 44324 26796
rect 44380 26786 44436 26796
rect 44492 26516 44548 26526
rect 44492 26422 44548 26460
rect 44940 25620 44996 26852
rect 45052 26852 45108 26862
rect 45052 26514 45108 26796
rect 45052 26462 45054 26514
rect 45106 26462 45108 26514
rect 45052 26450 45108 26462
rect 45388 26290 45444 26302
rect 45388 26238 45390 26290
rect 45442 26238 45444 26290
rect 45388 25732 45444 26238
rect 45500 26180 45556 27804
rect 45500 26114 45556 26124
rect 44940 25618 45332 25620
rect 44940 25566 44942 25618
rect 44994 25566 45332 25618
rect 44940 25564 45332 25566
rect 44940 25554 44996 25564
rect 45276 25506 45332 25564
rect 45276 25454 45278 25506
rect 45330 25454 45332 25506
rect 45276 25442 45332 25454
rect 45388 25284 45444 25676
rect 45276 25228 45444 25284
rect 45612 25284 45668 28812
rect 45276 25172 45332 25228
rect 45612 25218 45668 25228
rect 45948 25506 46004 25518
rect 45948 25454 45950 25506
rect 46002 25454 46004 25506
rect 45164 25116 45332 25172
rect 44828 24724 44884 24734
rect 44828 24722 44996 24724
rect 44828 24670 44830 24722
rect 44882 24670 44996 24722
rect 44828 24668 44996 24670
rect 44828 24658 44884 24668
rect 44492 24500 44548 24510
rect 44492 24498 44884 24500
rect 44492 24446 44494 24498
rect 44546 24446 44884 24498
rect 44492 24444 44884 24446
rect 44492 24434 44548 24444
rect 44380 23714 44436 23726
rect 44380 23662 44382 23714
rect 44434 23662 44436 23714
rect 44380 23492 44436 23662
rect 44380 23426 44436 23436
rect 44828 22708 44884 24444
rect 44828 22642 44884 22652
rect 44940 22484 44996 24668
rect 45052 24052 45108 24062
rect 45164 24052 45220 25116
rect 45276 24722 45332 24734
rect 45276 24670 45278 24722
rect 45330 24670 45332 24722
rect 45276 24276 45332 24670
rect 45276 24210 45332 24220
rect 45052 24050 45220 24052
rect 45052 23998 45054 24050
rect 45106 23998 45220 24050
rect 45052 23996 45220 23998
rect 45052 23986 45108 23996
rect 44828 22428 44996 22484
rect 45276 23938 45332 23950
rect 45276 23886 45278 23938
rect 45330 23886 45332 23938
rect 44828 22370 44884 22428
rect 44828 22318 44830 22370
rect 44882 22318 44884 22370
rect 44828 22260 44884 22318
rect 44828 22204 44996 22260
rect 44380 22148 44436 22158
rect 44940 22148 44996 22204
rect 44380 22146 44660 22148
rect 44380 22094 44382 22146
rect 44434 22094 44660 22146
rect 44380 22092 44660 22094
rect 44380 22082 44436 22092
rect 44268 21868 44548 21924
rect 44268 20690 44324 20702
rect 44268 20638 44270 20690
rect 44322 20638 44324 20690
rect 44268 19684 44324 20638
rect 44268 19618 44324 19628
rect 44380 19348 44436 19358
rect 44380 19254 44436 19292
rect 44492 19124 44548 21868
rect 44492 19058 44548 19068
rect 44604 18676 44660 22092
rect 44716 21586 44772 21598
rect 44716 21534 44718 21586
rect 44770 21534 44772 21586
rect 44716 20020 44772 21534
rect 44940 20802 44996 22092
rect 45276 21812 45332 23886
rect 45836 23938 45892 23950
rect 45836 23886 45838 23938
rect 45890 23886 45892 23938
rect 45836 22708 45892 23886
rect 45836 22642 45892 22652
rect 45388 22370 45444 22382
rect 45388 22318 45390 22370
rect 45442 22318 45444 22370
rect 45388 22036 45444 22318
rect 45388 21970 45444 21980
rect 45612 21924 45668 21934
rect 45612 21812 45668 21868
rect 45276 21810 45668 21812
rect 45276 21758 45614 21810
rect 45666 21758 45668 21810
rect 45276 21756 45668 21758
rect 45276 21586 45332 21756
rect 45276 21534 45278 21586
rect 45330 21534 45332 21586
rect 45276 21522 45332 21534
rect 44940 20750 44942 20802
rect 44994 20750 44996 20802
rect 44940 20738 44996 20750
rect 45388 20802 45444 20814
rect 45388 20750 45390 20802
rect 45442 20750 45444 20802
rect 45052 20132 45108 20142
rect 45052 20038 45108 20076
rect 44716 19954 44772 19964
rect 45388 19908 45444 20750
rect 45388 19842 45444 19852
rect 45052 19348 45108 19358
rect 45500 19348 45556 21756
rect 45612 21746 45668 21756
rect 45108 19346 45556 19348
rect 45108 19294 45502 19346
rect 45554 19294 45556 19346
rect 45108 19292 45556 19294
rect 45052 19254 45108 19292
rect 45500 19282 45556 19292
rect 45724 21588 45780 21598
rect 44604 18610 44660 18620
rect 45724 18562 45780 21532
rect 45948 21588 46004 25454
rect 46060 23828 46116 30716
rect 46284 30212 46340 30222
rect 46284 30118 46340 30156
rect 46732 30212 46788 30222
rect 46284 29652 46340 29662
rect 46284 29558 46340 29596
rect 46732 29650 46788 30156
rect 46732 29598 46734 29650
rect 46786 29598 46788 29650
rect 46732 29586 46788 29598
rect 46844 30098 46900 30110
rect 46844 30046 46846 30098
rect 46898 30046 46900 30098
rect 46844 29652 46900 30046
rect 47740 30100 47796 31166
rect 48076 30324 48132 32508
rect 48524 32452 48580 33294
rect 48748 33236 48804 34412
rect 49308 34356 49364 34366
rect 48860 34132 48916 34142
rect 48860 34038 48916 34076
rect 49308 34130 49364 34300
rect 49308 34078 49310 34130
rect 49362 34078 49364 34130
rect 49308 34066 49364 34078
rect 49196 33348 49252 33358
rect 49196 33254 49252 33292
rect 48748 33170 48804 33180
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51100 32788 51156 35646
rect 51324 35252 51380 36430
rect 52556 36484 52612 36494
rect 52612 36428 52724 36484
rect 52556 36390 52612 36428
rect 51324 35186 51380 35196
rect 52108 35252 52164 35262
rect 52108 35026 52164 35196
rect 52108 34974 52110 35026
rect 52162 34974 52164 35026
rect 52108 34962 52164 34974
rect 52668 34914 52724 36428
rect 53228 36482 53284 36540
rect 53228 36430 53230 36482
rect 53282 36430 53284 36482
rect 53228 36418 53284 36430
rect 52668 34862 52670 34914
rect 52722 34862 52724 34914
rect 52668 34850 52724 34862
rect 53340 34914 53396 38108
rect 53900 37380 53956 37390
rect 53900 37286 53956 37324
rect 54236 37268 54292 37278
rect 54236 37174 54292 37212
rect 53676 37042 53732 37054
rect 53676 36990 53678 37042
rect 53730 36990 53732 37042
rect 53676 36372 53732 36990
rect 53676 36306 53732 36316
rect 53676 35924 53732 35934
rect 53676 35830 53732 35868
rect 54348 35700 54404 38668
rect 54460 38658 54516 38668
rect 54684 37380 54740 37390
rect 54684 37266 54740 37324
rect 54908 37378 54964 40460
rect 55356 40450 55412 40460
rect 55468 40516 55524 40526
rect 55468 38946 55524 40460
rect 55468 38894 55470 38946
rect 55522 38894 55524 38946
rect 55468 38882 55524 38894
rect 54908 37326 54910 37378
rect 54962 37326 54964 37378
rect 54908 37314 54964 37326
rect 55580 37380 55636 41244
rect 55692 40962 55748 43374
rect 56140 41970 56196 43596
rect 56700 43540 56756 44380
rect 57148 44370 57204 44380
rect 57596 44994 57652 45006
rect 57596 44942 57598 44994
rect 57650 44942 57652 44994
rect 57596 44324 57652 44942
rect 58828 44884 58884 45166
rect 58828 44818 58884 44828
rect 58940 45220 58996 45230
rect 58940 44434 58996 45164
rect 58940 44382 58942 44434
rect 58994 44382 58996 44434
rect 58940 44370 58996 44382
rect 59500 44994 59556 45612
rect 60620 45668 60676 45678
rect 60620 45574 60676 45612
rect 61404 45218 61460 46396
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 61404 45166 61406 45218
rect 61458 45166 61460 45218
rect 61404 45154 61460 45166
rect 59500 44942 59502 44994
rect 59554 44942 59556 44994
rect 57596 44258 57652 44268
rect 58492 44322 58548 44334
rect 58492 44270 58494 44322
rect 58546 44270 58548 44322
rect 58268 44212 58324 44222
rect 58268 44118 58324 44156
rect 57596 44100 57652 44110
rect 56700 43426 56756 43484
rect 56700 43374 56702 43426
rect 56754 43374 56756 43426
rect 56588 42756 56644 42766
rect 56700 42756 56756 43374
rect 56588 42754 56756 42756
rect 56588 42702 56590 42754
rect 56642 42702 56756 42754
rect 56588 42700 56756 42702
rect 56588 42690 56644 42700
rect 56252 42644 56308 42654
rect 56252 42550 56308 42588
rect 56140 41918 56142 41970
rect 56194 41918 56196 41970
rect 56140 41906 56196 41918
rect 56252 42084 56308 42094
rect 56252 41410 56308 42028
rect 56252 41358 56254 41410
rect 56306 41358 56308 41410
rect 56252 41346 56308 41358
rect 56700 41972 56756 42700
rect 56700 41298 56756 41916
rect 56700 41246 56702 41298
rect 56754 41246 56756 41298
rect 56700 41234 56756 41246
rect 56812 43764 56868 43774
rect 56812 41300 56868 43708
rect 57148 43428 57204 43438
rect 57148 43334 57204 43372
rect 57596 43426 57652 44044
rect 58492 43764 58548 44270
rect 58492 43698 58548 43708
rect 59276 44212 59332 44222
rect 59500 44212 59556 44942
rect 60396 44996 60452 45006
rect 60396 44902 60452 44940
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 61516 44436 61572 44446
rect 61516 44342 61572 44380
rect 59276 44210 59556 44212
rect 59276 44158 59278 44210
rect 59330 44158 59556 44210
rect 59276 44156 59556 44158
rect 60060 44212 60116 44222
rect 57596 43374 57598 43426
rect 57650 43374 57652 43426
rect 57596 43362 57652 43374
rect 58828 43650 58884 43662
rect 58828 43598 58830 43650
rect 58882 43598 58884 43650
rect 58828 43204 58884 43598
rect 59276 43428 59332 44156
rect 59724 44098 59780 44110
rect 59724 44046 59726 44098
rect 59778 44046 59780 44098
rect 59500 43764 59556 43802
rect 59724 43764 59780 44046
rect 59556 43708 59780 43764
rect 59500 43698 59556 43708
rect 59276 43362 59332 43372
rect 58828 43138 58884 43148
rect 57036 42868 57092 42878
rect 57036 42754 57092 42812
rect 57036 42702 57038 42754
rect 57090 42702 57092 42754
rect 57036 42690 57092 42702
rect 59388 42530 59444 42542
rect 59388 42478 59390 42530
rect 59442 42478 59444 42530
rect 58828 42420 58884 42430
rect 58828 42082 58884 42364
rect 58828 42030 58830 42082
rect 58882 42030 58884 42082
rect 58828 42018 58884 42030
rect 59276 42196 59332 42206
rect 57148 41858 57204 41870
rect 57148 41806 57150 41858
rect 57202 41806 57204 41858
rect 55692 40910 55694 40962
rect 55746 40910 55748 40962
rect 55692 40898 55748 40910
rect 56140 40740 56196 40750
rect 56140 40626 56196 40684
rect 56140 40574 56142 40626
rect 56194 40574 56196 40626
rect 56140 40562 56196 40574
rect 56700 40628 56756 40638
rect 56812 40628 56868 41244
rect 57036 41300 57092 41310
rect 57148 41300 57204 41806
rect 57596 41860 57652 41870
rect 57596 41766 57652 41804
rect 57036 41298 57204 41300
rect 57036 41246 57038 41298
rect 57090 41246 57204 41298
rect 57036 41244 57204 41246
rect 57036 41234 57092 41244
rect 57148 40628 57204 41244
rect 56700 40626 56868 40628
rect 56700 40574 56702 40626
rect 56754 40574 56868 40626
rect 56700 40572 56868 40574
rect 57036 40626 57204 40628
rect 57036 40574 57150 40626
rect 57202 40574 57204 40626
rect 57036 40572 57204 40574
rect 56700 40562 56756 40572
rect 57036 39732 57092 40572
rect 57148 40562 57204 40572
rect 57484 41298 57540 41310
rect 57484 41246 57486 41298
rect 57538 41246 57540 41298
rect 56812 39730 57092 39732
rect 56812 39678 57038 39730
rect 57090 39678 57092 39730
rect 56812 39676 57092 39678
rect 55916 39396 55972 39406
rect 55580 37314 55636 37324
rect 55804 39394 55972 39396
rect 55804 39342 55918 39394
rect 55970 39342 55972 39394
rect 55804 39340 55972 39342
rect 55804 37378 55860 39340
rect 55916 39330 55972 39340
rect 56700 39396 56756 39406
rect 56700 39302 56756 39340
rect 56700 39060 56756 39070
rect 56812 39060 56868 39676
rect 57036 39666 57092 39676
rect 56700 39058 56868 39060
rect 56700 39006 56702 39058
rect 56754 39006 56868 39058
rect 56700 39004 56868 39006
rect 57484 39060 57540 41246
rect 59276 41298 59332 42140
rect 59388 41860 59444 42478
rect 59500 41972 59556 41982
rect 59500 41878 59556 41916
rect 59388 41794 59444 41804
rect 59612 41748 59668 43708
rect 60060 42978 60116 44156
rect 62524 44212 62580 44222
rect 62524 44118 62580 44156
rect 61404 43652 61460 43662
rect 61404 43558 61460 43596
rect 60396 43428 60452 43438
rect 60396 43334 60452 43372
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 60060 42926 60062 42978
rect 60114 42926 60116 42978
rect 60060 42914 60116 42926
rect 61516 42868 61572 42878
rect 61516 42774 61572 42812
rect 62524 42644 62580 42654
rect 62524 42550 62580 42588
rect 61404 42084 61460 42094
rect 61404 41990 61460 42028
rect 62412 41970 62468 41982
rect 62412 41918 62414 41970
rect 62466 41918 62468 41970
rect 59612 41300 59668 41692
rect 59276 41246 59278 41298
rect 59330 41246 59332 41298
rect 59276 41234 59332 41246
rect 59500 41298 59668 41300
rect 59500 41246 59614 41298
rect 59666 41246 59668 41298
rect 59500 41244 59668 41246
rect 58492 41076 58548 41086
rect 58492 40982 58548 41020
rect 59500 40626 59556 41244
rect 59612 41234 59668 41244
rect 60396 41858 60452 41870
rect 60396 41806 60398 41858
rect 60450 41806 60452 41858
rect 60396 41188 60452 41806
rect 62188 41860 62244 41870
rect 62188 41766 62244 41804
rect 62412 41748 62468 41918
rect 62412 41682 62468 41692
rect 62972 41858 63028 41870
rect 62972 41806 62974 41858
rect 63026 41806 63028 41858
rect 62972 41748 63028 41806
rect 62972 41682 63028 41692
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 60396 41122 60452 41132
rect 61740 41298 61796 41310
rect 61740 41246 61742 41298
rect 61794 41246 61796 41298
rect 59500 40574 59502 40626
rect 59554 40574 59556 40626
rect 59500 40562 59556 40574
rect 61404 40964 61460 40974
rect 58828 40516 58884 40526
rect 58828 40422 58884 40460
rect 61404 40514 61460 40908
rect 61404 40462 61406 40514
rect 61458 40462 61460 40514
rect 61404 40450 61460 40462
rect 61516 40404 61572 40414
rect 57596 40290 57652 40302
rect 57596 40238 57598 40290
rect 57650 40238 57652 40290
rect 57596 39844 57652 40238
rect 60396 40290 60452 40302
rect 60396 40238 60398 40290
rect 60450 40238 60452 40290
rect 60396 40068 60452 40238
rect 60396 40002 60452 40012
rect 57596 39778 57652 39788
rect 58940 39956 58996 39966
rect 57932 39732 57988 39742
rect 57932 39638 57988 39676
rect 56700 38836 56756 39004
rect 57484 38994 57540 39004
rect 57596 39620 57652 39630
rect 56700 38162 56756 38780
rect 57596 38722 57652 39564
rect 58940 39506 58996 39900
rect 61516 39730 61572 40348
rect 61740 40180 61796 41246
rect 62524 41074 62580 41086
rect 62524 41022 62526 41074
rect 62578 41022 62580 41074
rect 62524 40740 62580 41022
rect 62524 40674 62580 40684
rect 61740 40114 61796 40124
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 61516 39678 61518 39730
rect 61570 39678 61572 39730
rect 61516 39666 61572 39678
rect 58940 39454 58942 39506
rect 58994 39454 58996 39506
rect 58940 39442 58996 39454
rect 62524 39506 62580 39518
rect 62524 39454 62526 39506
rect 62578 39454 62580 39506
rect 61404 39396 61460 39406
rect 57596 38670 57598 38722
rect 57650 38670 57652 38722
rect 57596 38658 57652 38670
rect 58828 38946 58884 38958
rect 58828 38894 58830 38946
rect 58882 38894 58884 38946
rect 56700 38110 56702 38162
rect 56754 38110 56756 38162
rect 56700 38098 56756 38110
rect 57596 38276 57652 38286
rect 55804 37326 55806 37378
rect 55858 37326 55860 37378
rect 55804 37314 55860 37326
rect 56700 37380 56756 37390
rect 56700 37286 56756 37324
rect 54684 37214 54686 37266
rect 54738 37214 54740 37266
rect 54684 37202 54740 37214
rect 55468 37268 55524 37278
rect 55468 37156 55524 37212
rect 55468 37154 55636 37156
rect 55468 37102 55470 37154
rect 55522 37102 55636 37154
rect 55468 37100 55636 37102
rect 55468 37090 55524 37100
rect 55468 36260 55524 36270
rect 55132 36258 55524 36260
rect 55132 36206 55470 36258
rect 55522 36206 55524 36258
rect 55132 36204 55524 36206
rect 54348 35634 54404 35644
rect 54460 35924 54516 35934
rect 53340 34862 53342 34914
rect 53394 34862 53396 34914
rect 53340 34850 53396 34862
rect 54236 35474 54292 35486
rect 54236 35422 54238 35474
rect 54290 35422 54292 35474
rect 51212 34804 51268 34814
rect 51212 34802 51604 34804
rect 51212 34750 51214 34802
rect 51266 34750 51604 34802
rect 51212 34748 51604 34750
rect 51212 34738 51268 34748
rect 51548 34354 51604 34748
rect 51548 34302 51550 34354
rect 51602 34302 51604 34354
rect 51548 34290 51604 34302
rect 51772 34802 51828 34814
rect 51772 34750 51774 34802
rect 51826 34750 51828 34802
rect 51436 33796 51492 33806
rect 51212 32788 51268 32798
rect 51100 32732 51212 32788
rect 51212 32722 51268 32732
rect 50764 32674 50820 32686
rect 50764 32622 50766 32674
rect 50818 32622 50820 32674
rect 48860 32452 48916 32462
rect 49308 32452 49364 32462
rect 48580 32450 48916 32452
rect 48580 32398 48862 32450
rect 48914 32398 48916 32450
rect 48580 32396 48916 32398
rect 48524 32386 48580 32396
rect 48300 31892 48356 31902
rect 48300 31218 48356 31836
rect 48300 31166 48302 31218
rect 48354 31166 48356 31218
rect 48300 31154 48356 31166
rect 48412 31554 48468 31566
rect 48412 31502 48414 31554
rect 48466 31502 48468 31554
rect 48076 30258 48132 30268
rect 47740 30034 47796 30044
rect 47180 29652 47236 29662
rect 46900 29650 47236 29652
rect 46900 29598 47182 29650
rect 47234 29598 47236 29650
rect 46900 29596 47236 29598
rect 46844 29586 46900 29596
rect 47180 29586 47236 29596
rect 47964 29314 48020 29326
rect 47964 29262 47966 29314
rect 48018 29262 48020 29314
rect 47740 28756 47796 28766
rect 47740 28082 47796 28700
rect 47740 28030 47742 28082
rect 47794 28030 47796 28082
rect 47740 28018 47796 28030
rect 47852 28418 47908 28430
rect 47852 28366 47854 28418
rect 47906 28366 47908 28418
rect 47852 27748 47908 28366
rect 47852 27682 47908 27692
rect 47964 26908 48020 29262
rect 48188 29314 48244 29326
rect 48188 29262 48190 29314
rect 48242 29262 48244 29314
rect 48188 28980 48244 29262
rect 48188 28914 48244 28924
rect 48412 27972 48468 31502
rect 48748 31554 48804 32396
rect 48860 32386 48916 32396
rect 49196 32450 49364 32452
rect 49196 32398 49310 32450
rect 49362 32398 49364 32450
rect 49196 32396 49364 32398
rect 49196 31556 49252 32396
rect 49308 32386 49364 32396
rect 49756 32452 49812 32462
rect 49756 32358 49812 32396
rect 50764 32340 50820 32622
rect 50764 32274 50820 32284
rect 48748 31502 48750 31554
rect 48802 31502 48804 31554
rect 48748 30996 48804 31502
rect 49084 31554 49252 31556
rect 49084 31502 49198 31554
rect 49250 31502 49252 31554
rect 49084 31500 49252 31502
rect 49084 30996 49140 31500
rect 49196 31490 49252 31500
rect 49644 31890 49700 31902
rect 51436 31892 51492 33740
rect 51660 33124 51716 33134
rect 51772 33124 51828 34750
rect 53676 34468 53732 34478
rect 52332 34356 52388 34366
rect 52332 34262 52388 34300
rect 52444 34132 52500 34142
rect 52500 34076 52836 34132
rect 52444 34038 52500 34076
rect 52780 33458 52836 34076
rect 53116 34130 53172 34142
rect 53116 34078 53118 34130
rect 53170 34078 53172 34130
rect 53116 33684 53172 34078
rect 53116 33618 53172 33628
rect 52780 33406 52782 33458
rect 52834 33406 52836 33458
rect 51660 33122 51828 33124
rect 51660 33070 51662 33122
rect 51714 33070 51828 33122
rect 51660 33068 51828 33070
rect 52220 33124 52276 33134
rect 51660 33058 51716 33068
rect 52220 33030 52276 33068
rect 49644 31838 49646 31890
rect 49698 31838 49700 31890
rect 48748 30994 49140 30996
rect 48748 30942 48750 30994
rect 48802 30942 49140 30994
rect 48748 30940 49140 30942
rect 49308 30996 49364 31006
rect 48748 30930 48804 30940
rect 48748 30324 48804 30334
rect 48524 28868 48580 28878
rect 48524 28774 48580 28812
rect 48748 28642 48804 30268
rect 48748 28590 48750 28642
rect 48802 28590 48804 28642
rect 48748 28532 48804 28590
rect 48412 27906 48468 27916
rect 48636 28476 48804 28532
rect 48860 29426 48916 29438
rect 48860 29374 48862 29426
rect 48914 29374 48916 29426
rect 48300 27634 48356 27646
rect 48300 27582 48302 27634
rect 48354 27582 48356 27634
rect 47852 26850 47908 26862
rect 47964 26852 48244 26908
rect 47852 26798 47854 26850
rect 47906 26798 47908 26850
rect 46956 26178 47012 26190
rect 46956 26126 46958 26178
rect 47010 26126 47012 26178
rect 46956 26068 47012 26126
rect 46956 26002 47012 26012
rect 47628 25284 47684 25294
rect 47628 24724 47684 25228
rect 47740 24948 47796 24958
rect 47740 24854 47796 24892
rect 47628 24668 47796 24724
rect 46060 23762 46116 23772
rect 46508 24164 46564 24174
rect 46060 23492 46116 23502
rect 46116 23436 46228 23492
rect 46060 23426 46116 23436
rect 46060 23156 46116 23166
rect 46060 21924 46116 23100
rect 46060 21810 46116 21868
rect 46060 21758 46062 21810
rect 46114 21758 46116 21810
rect 46060 21746 46116 21758
rect 45948 21522 46004 21532
rect 46060 21476 46116 21486
rect 45836 19796 45892 19806
rect 45836 19794 46004 19796
rect 45836 19742 45838 19794
rect 45890 19742 46004 19794
rect 45836 19740 46004 19742
rect 45836 19730 45892 19740
rect 45724 18510 45726 18562
rect 45778 18510 45780 18562
rect 45724 18498 45780 18510
rect 45836 19012 45892 19022
rect 44716 18340 44772 18350
rect 44156 18338 44772 18340
rect 44156 18286 44718 18338
rect 44770 18286 44772 18338
rect 44156 18284 44772 18286
rect 44716 18274 44772 18284
rect 43036 16942 43038 16994
rect 43090 16942 43092 16994
rect 43036 16930 43092 16942
rect 44716 18116 44772 18126
rect 44716 16770 44772 18060
rect 45836 17778 45892 18956
rect 45836 17726 45838 17778
rect 45890 17726 45892 17778
rect 45836 17714 45892 17726
rect 45948 17556 46004 19740
rect 46060 19346 46116 21420
rect 46060 19294 46062 19346
rect 46114 19294 46116 19346
rect 46060 19282 46116 19294
rect 45948 17490 46004 17500
rect 46060 16996 46116 17006
rect 46172 16996 46228 23436
rect 46284 22260 46340 22270
rect 46284 20242 46340 22204
rect 46508 21474 46564 24108
rect 46956 23156 47012 23166
rect 46956 23042 47012 23100
rect 46956 22990 46958 23042
rect 47010 22990 47012 23042
rect 46956 22978 47012 22990
rect 47628 22148 47684 22158
rect 46508 21422 46510 21474
rect 46562 21422 46564 21474
rect 46508 21410 46564 21422
rect 47180 22146 47684 22148
rect 47180 22094 47630 22146
rect 47682 22094 47684 22146
rect 47180 22092 47684 22094
rect 46284 20190 46286 20242
rect 46338 20190 46340 20242
rect 46284 20178 46340 20190
rect 46732 20132 46788 20142
rect 46732 20038 46788 20076
rect 47068 20132 47124 20142
rect 46396 19908 46452 19918
rect 47068 19908 47124 20076
rect 46396 19906 47124 19908
rect 46396 19854 46398 19906
rect 46450 19854 47124 19906
rect 46396 19852 47124 19854
rect 46396 19684 46452 19852
rect 46396 19618 46452 19628
rect 46844 18564 46900 19852
rect 47068 19124 47124 19134
rect 47068 19030 47124 19068
rect 46844 18470 46900 18508
rect 47068 18452 47124 18462
rect 47068 17554 47124 18396
rect 47180 18450 47236 22092
rect 47628 22082 47684 22092
rect 47740 21698 47796 24668
rect 47852 23378 47908 26798
rect 48188 25394 48244 26852
rect 48188 25342 48190 25394
rect 48242 25342 48244 25394
rect 48188 25330 48244 25342
rect 48300 24724 48356 27582
rect 48636 27636 48692 28476
rect 48860 28420 48916 29374
rect 48748 28364 48916 28420
rect 48748 27860 48804 28364
rect 48860 28084 48916 28094
rect 48972 28084 49028 30940
rect 49308 30902 49364 30940
rect 49644 29988 49700 31838
rect 50988 31890 51492 31892
rect 50988 31838 51438 31890
rect 51490 31838 51492 31890
rect 50988 31836 51492 31838
rect 50876 31666 50932 31678
rect 50876 31614 50878 31666
rect 50930 31614 50932 31666
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50876 30548 50932 31614
rect 50876 30482 50932 30492
rect 50764 30324 50820 30334
rect 50988 30324 51044 31836
rect 51436 31826 51492 31836
rect 52220 32450 52276 32462
rect 52220 32398 52222 32450
rect 52274 32398 52276 32450
rect 51548 31556 51604 31566
rect 51548 31462 51604 31500
rect 50764 30322 51044 30324
rect 50764 30270 50766 30322
rect 50818 30270 51044 30322
rect 50764 30268 51044 30270
rect 51548 31106 51604 31118
rect 51548 31054 51550 31106
rect 51602 31054 51604 31106
rect 50764 30258 50820 30268
rect 50428 30100 50484 30110
rect 50428 30006 50484 30044
rect 49644 29922 49700 29932
rect 51212 29986 51268 29998
rect 51212 29934 51214 29986
rect 51266 29934 51268 29986
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 49308 29428 49364 29438
rect 49308 29334 49364 29372
rect 49756 28980 49812 28990
rect 49644 28084 49700 28094
rect 48860 28082 49644 28084
rect 48860 28030 48862 28082
rect 48914 28030 49644 28082
rect 48860 28028 49644 28030
rect 48860 28018 48916 28028
rect 48748 27794 48804 27804
rect 49196 27748 49252 27758
rect 49196 27654 49252 27692
rect 49532 27748 49588 27758
rect 49532 27654 49588 27692
rect 48636 27580 49140 27636
rect 49084 27076 49140 27580
rect 49084 26908 49140 27020
rect 48412 26850 48468 26862
rect 49084 26852 49252 26908
rect 48412 26798 48414 26850
rect 48466 26798 48468 26850
rect 48412 25620 48468 26798
rect 49084 26516 49140 26526
rect 48860 26290 48916 26302
rect 48860 26238 48862 26290
rect 48914 26238 48916 26290
rect 48412 25554 48468 25564
rect 48748 26068 48804 26078
rect 48748 24834 48804 26012
rect 48748 24782 48750 24834
rect 48802 24782 48804 24834
rect 48748 24770 48804 24782
rect 48860 24724 48916 26238
rect 48972 25508 49028 25518
rect 48972 25414 49028 25452
rect 49084 24834 49140 26460
rect 49084 24782 49086 24834
rect 49138 24782 49140 24834
rect 49084 24770 49140 24782
rect 49196 25732 49252 26852
rect 49196 25506 49252 25676
rect 49196 25454 49198 25506
rect 49250 25454 49252 25506
rect 49196 24836 49252 25454
rect 49308 26290 49364 26302
rect 49308 26238 49310 26290
rect 49362 26238 49364 26290
rect 49308 25396 49364 26238
rect 49308 25330 49364 25340
rect 48300 24668 48580 24724
rect 48300 24498 48356 24510
rect 48300 24446 48302 24498
rect 48354 24446 48356 24498
rect 48076 23714 48132 23726
rect 48076 23662 48078 23714
rect 48130 23662 48132 23714
rect 47852 23326 47854 23378
rect 47906 23326 47908 23378
rect 47852 23314 47908 23326
rect 47964 23604 48020 23614
rect 47740 21646 47742 21698
rect 47794 21646 47796 21698
rect 47740 21634 47796 21646
rect 47964 23266 48020 23548
rect 47964 23214 47966 23266
rect 48018 23214 48020 23266
rect 47964 21364 48020 23214
rect 47516 21308 48020 21364
rect 47516 20132 47572 21308
rect 47516 20018 47572 20076
rect 47740 20578 47796 20590
rect 47740 20526 47742 20578
rect 47794 20526 47796 20578
rect 47740 20130 47796 20526
rect 47740 20078 47742 20130
rect 47794 20078 47796 20130
rect 47740 20066 47796 20078
rect 47516 19966 47518 20018
rect 47570 19966 47572 20018
rect 47516 19954 47572 19966
rect 47852 18564 47908 18574
rect 47852 18470 47908 18508
rect 47180 18398 47182 18450
rect 47234 18398 47236 18450
rect 47180 18386 47236 18398
rect 48076 18338 48132 23662
rect 48300 22596 48356 24446
rect 48300 22530 48356 22540
rect 48412 22260 48468 22270
rect 48412 22166 48468 22204
rect 48524 22148 48580 24668
rect 48860 23940 48916 24668
rect 49196 24052 49252 24780
rect 49420 24612 49476 24622
rect 49420 24518 49476 24556
rect 49308 24052 49364 24062
rect 49644 24052 49700 28028
rect 49756 27748 49812 28924
rect 51100 28980 51156 28990
rect 51100 28754 51156 28924
rect 51100 28702 51102 28754
rect 51154 28702 51156 28754
rect 49980 28644 50036 28654
rect 49980 27860 50036 28588
rect 49980 27766 50036 27804
rect 50316 28420 50372 28430
rect 49756 27682 49812 27692
rect 49196 24050 49364 24052
rect 49196 23998 49310 24050
rect 49362 23998 49364 24050
rect 49196 23996 49364 23998
rect 49308 23986 49364 23996
rect 49420 24050 49700 24052
rect 49420 23998 49646 24050
rect 49698 23998 49700 24050
rect 49420 23996 49700 23998
rect 48748 23884 48916 23940
rect 48636 22372 48692 22382
rect 48748 22372 48804 23884
rect 48860 23714 48916 23726
rect 48860 23662 48862 23714
rect 48914 23662 48916 23714
rect 48860 23380 48916 23662
rect 48860 23314 48916 23324
rect 48860 23156 48916 23166
rect 49308 23156 49364 23166
rect 48916 23100 49028 23156
rect 48860 23062 48916 23100
rect 48636 22370 48916 22372
rect 48636 22318 48638 22370
rect 48690 22318 48916 22370
rect 48636 22316 48916 22318
rect 48636 22306 48692 22316
rect 48860 22148 48916 22316
rect 48524 22092 48692 22148
rect 48524 21812 48580 21822
rect 48412 21028 48468 21038
rect 48412 20934 48468 20972
rect 48188 20132 48244 20142
rect 48188 20038 48244 20076
rect 48076 18286 48078 18338
rect 48130 18286 48132 18338
rect 48076 18274 48132 18286
rect 48524 17780 48580 21756
rect 48636 20244 48692 22092
rect 48860 21586 48916 22092
rect 48860 21534 48862 21586
rect 48914 21534 48916 21586
rect 48860 21522 48916 21534
rect 48636 20178 48692 20188
rect 48860 20132 48916 20142
rect 48972 20132 49028 23100
rect 49308 23062 49364 23100
rect 49420 22932 49476 23996
rect 49644 23986 49700 23996
rect 49756 27186 49812 27198
rect 49756 27134 49758 27186
rect 49810 27134 49812 27186
rect 49756 24836 49812 27134
rect 50316 26404 50372 28364
rect 51100 28420 51156 28702
rect 51100 28354 51156 28364
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 51212 28084 51268 29934
rect 51212 28018 51268 28028
rect 50652 27858 50708 27870
rect 50652 27806 50654 27858
rect 50706 27806 50708 27858
rect 50652 27412 50708 27806
rect 50652 27346 50708 27356
rect 51548 27186 51604 31054
rect 52220 30212 52276 32398
rect 52556 32450 52612 32462
rect 52556 32398 52558 32450
rect 52610 32398 52612 32450
rect 52556 30884 52612 32398
rect 52780 31780 52836 33406
rect 53676 33458 53732 34412
rect 53676 33406 53678 33458
rect 53730 33406 53732 33458
rect 53676 33394 53732 33406
rect 53900 32900 53956 32910
rect 53788 32674 53844 32686
rect 53788 32622 53790 32674
rect 53842 32622 53844 32674
rect 53788 32004 53844 32622
rect 53900 32564 53956 32844
rect 54236 32900 54292 35422
rect 54236 32834 54292 32844
rect 53900 32498 53956 32508
rect 54460 32450 54516 35868
rect 55132 35810 55188 36204
rect 55468 36194 55524 36204
rect 55132 35758 55134 35810
rect 55186 35758 55188 35810
rect 55132 35746 55188 35758
rect 54908 35698 54964 35710
rect 54908 35646 54910 35698
rect 54962 35646 54964 35698
rect 54908 35476 54964 35646
rect 54908 35410 54964 35420
rect 55580 35698 55636 37100
rect 57596 37154 57652 38220
rect 58828 38052 58884 38894
rect 61404 38946 61460 39340
rect 61404 38894 61406 38946
rect 61458 38894 61460 38946
rect 61404 38882 61460 38894
rect 62524 38948 62580 39454
rect 62524 38882 62580 38892
rect 60396 38722 60452 38734
rect 60396 38670 60398 38722
rect 60450 38670 60452 38722
rect 60396 38388 60452 38670
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 60396 38322 60452 38332
rect 61516 38164 61572 38174
rect 61516 38070 61572 38108
rect 58828 37986 58884 37996
rect 62524 37938 62580 37950
rect 62524 37886 62526 37938
rect 62578 37886 62580 37938
rect 61404 37828 61460 37838
rect 57596 37102 57598 37154
rect 57650 37102 57652 37154
rect 57596 37090 57652 37102
rect 58828 37378 58884 37390
rect 58828 37326 58830 37378
rect 58882 37326 58884 37378
rect 58828 37044 58884 37326
rect 61404 37378 61460 37772
rect 61404 37326 61406 37378
rect 61458 37326 61460 37378
rect 61404 37314 61460 37326
rect 60396 37156 60452 37166
rect 60396 37062 60452 37100
rect 58828 36978 58884 36988
rect 57596 36932 57652 36942
rect 56252 36820 56308 36830
rect 56252 36706 56308 36764
rect 56252 36654 56254 36706
rect 56306 36654 56308 36706
rect 56252 36642 56308 36654
rect 56588 36484 56644 36494
rect 56588 35924 56644 36428
rect 56700 35924 56756 35934
rect 56588 35922 56756 35924
rect 56588 35870 56702 35922
rect 56754 35870 56756 35922
rect 56588 35868 56756 35870
rect 55580 35646 55582 35698
rect 55634 35646 55636 35698
rect 55580 35476 55636 35646
rect 55580 35410 55636 35420
rect 55692 35586 55748 35598
rect 55692 35534 55694 35586
rect 55746 35534 55748 35586
rect 54572 35252 54628 35262
rect 54572 32562 54628 35196
rect 55356 34692 55412 34702
rect 55356 34354 55412 34636
rect 55692 34690 55748 35534
rect 56364 35140 56420 35150
rect 56364 35046 56420 35084
rect 56700 35028 56756 35868
rect 57596 35586 57652 36876
rect 58492 36708 58548 36718
rect 57596 35534 57598 35586
rect 57650 35534 57652 35586
rect 57596 35522 57652 35534
rect 57708 36594 57764 36606
rect 57708 36542 57710 36594
rect 57762 36542 57764 36594
rect 56812 35028 56868 35038
rect 56700 35026 56868 35028
rect 56700 34974 56814 35026
rect 56866 34974 56868 35026
rect 56700 34972 56868 34974
rect 56812 34962 56868 34972
rect 57596 35028 57652 35038
rect 57596 34934 57652 34972
rect 55692 34638 55694 34690
rect 55746 34638 55748 34690
rect 55692 34626 55748 34638
rect 56140 34804 56196 34814
rect 55356 34302 55358 34354
rect 55410 34302 55412 34354
rect 55356 34290 55412 34302
rect 56140 34354 56196 34748
rect 56140 34302 56142 34354
rect 56194 34302 56196 34354
rect 56140 34290 56196 34302
rect 56812 34018 56868 34030
rect 56812 33966 56814 34018
rect 56866 33966 56868 34018
rect 54684 33460 54740 33470
rect 54684 33234 54740 33404
rect 54684 33182 54686 33234
rect 54738 33182 54740 33234
rect 54684 33170 54740 33182
rect 56476 33458 56532 33470
rect 56476 33406 56478 33458
rect 56530 33406 56532 33458
rect 56476 33012 56532 33406
rect 56476 32946 56532 32956
rect 54572 32510 54574 32562
rect 54626 32510 54628 32562
rect 54572 32498 54628 32510
rect 54460 32398 54462 32450
rect 54514 32398 54516 32450
rect 54460 32386 54516 32398
rect 53788 31938 53844 31948
rect 52556 30818 52612 30828
rect 52668 31778 52836 31780
rect 52668 31726 52782 31778
rect 52834 31726 52836 31778
rect 52668 31724 52836 31726
rect 52668 30994 52724 31724
rect 52780 31714 52836 31724
rect 53228 31892 53284 31902
rect 53228 31778 53284 31836
rect 53228 31726 53230 31778
rect 53282 31726 53284 31778
rect 53228 31714 53284 31726
rect 55692 31554 55748 31566
rect 55692 31502 55694 31554
rect 55746 31502 55748 31554
rect 55356 31108 55412 31118
rect 54572 31106 55412 31108
rect 54572 31054 55358 31106
rect 55410 31054 55412 31106
rect 54572 31052 55412 31054
rect 52668 30942 52670 30994
rect 52722 30942 52724 30994
rect 52332 30772 52388 30782
rect 52332 30678 52388 30716
rect 52220 30146 52276 30156
rect 52668 30324 52724 30942
rect 53116 30996 53172 31006
rect 53116 30994 53284 30996
rect 53116 30942 53118 30994
rect 53170 30942 53284 30994
rect 53116 30940 53284 30942
rect 53116 30930 53172 30940
rect 51660 30098 51716 30110
rect 51660 30046 51662 30098
rect 51714 30046 51716 30098
rect 51660 29650 51716 30046
rect 51660 29598 51662 29650
rect 51714 29598 51716 29650
rect 51660 29586 51716 29598
rect 51996 30100 52052 30110
rect 51660 28756 51716 28766
rect 51660 28662 51716 28700
rect 51996 28756 52052 30044
rect 52332 29204 52388 29214
rect 52332 29110 52388 29148
rect 52444 29202 52500 29214
rect 52444 29150 52446 29202
rect 52498 29150 52500 29202
rect 51996 28420 52052 28700
rect 51548 27134 51550 27186
rect 51602 27134 51604 27186
rect 51548 27122 51604 27134
rect 51884 27188 51940 27198
rect 51996 27188 52052 28364
rect 52444 28420 52500 29150
rect 52444 28354 52500 28364
rect 52668 28644 52724 30268
rect 52780 30100 52836 30110
rect 52780 30006 52836 30044
rect 53116 30098 53172 30110
rect 53116 30046 53118 30098
rect 53170 30046 53172 30098
rect 53116 29650 53172 30046
rect 53228 29876 53284 30940
rect 53228 29810 53284 29820
rect 53900 30212 53956 30222
rect 53116 29598 53118 29650
rect 53170 29598 53172 29650
rect 53116 29586 53172 29598
rect 51884 27186 52052 27188
rect 51884 27134 51886 27186
rect 51938 27134 52052 27186
rect 51884 27132 52052 27134
rect 51884 27122 51940 27132
rect 50764 27076 50820 27086
rect 50764 26982 50820 27020
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50316 26338 50372 26348
rect 51772 26514 51828 26526
rect 51772 26462 51774 26514
rect 51826 26462 51828 26514
rect 51548 25618 51604 25630
rect 51548 25566 51550 25618
rect 51602 25566 51604 25618
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50204 24948 50260 24958
rect 50204 24854 50260 24892
rect 50092 24836 50148 24846
rect 49756 24834 50148 24836
rect 49756 24782 49758 24834
rect 49810 24782 50094 24834
rect 50146 24782 50148 24834
rect 49756 24780 50148 24782
rect 49756 23604 49812 24780
rect 50092 24770 50148 24780
rect 50876 24836 50932 24846
rect 50876 24742 50932 24780
rect 51212 24724 51268 24734
rect 51212 24630 51268 24668
rect 50092 24052 50148 24062
rect 50092 23958 50148 23996
rect 51100 23828 51156 23838
rect 51100 23734 51156 23772
rect 49756 23538 49812 23548
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 49196 22876 49476 22932
rect 49644 23380 49700 23390
rect 49084 22372 49140 22382
rect 49084 22278 49140 22316
rect 49196 20914 49252 22876
rect 49644 22148 49700 23324
rect 49644 22082 49700 22092
rect 50204 23156 50260 23166
rect 49644 21700 49700 21710
rect 49532 21586 49588 21598
rect 49532 21534 49534 21586
rect 49586 21534 49588 21586
rect 49532 21252 49588 21534
rect 49532 21186 49588 21196
rect 49196 20862 49198 20914
rect 49250 20862 49252 20914
rect 49196 20850 49252 20862
rect 49644 20914 49700 21644
rect 49644 20862 49646 20914
rect 49698 20862 49700 20914
rect 49644 20850 49700 20862
rect 49756 21588 49812 21598
rect 48916 20076 49028 20132
rect 48860 20038 48916 20076
rect 48636 20020 48692 20030
rect 48636 19346 48692 19964
rect 49756 19906 49812 21532
rect 49756 19854 49758 19906
rect 49810 19854 49812 19906
rect 49756 19842 49812 19854
rect 48636 19294 48638 19346
rect 48690 19294 48692 19346
rect 48636 19282 48692 19294
rect 49644 19796 49700 19806
rect 49644 19122 49700 19740
rect 49644 19070 49646 19122
rect 49698 19070 49700 19122
rect 49644 19058 49700 19070
rect 50204 18338 50260 23100
rect 50428 22596 50484 22606
rect 50428 21812 50484 22540
rect 51436 22148 51492 22158
rect 50876 22146 51492 22148
rect 50876 22094 51438 22146
rect 51490 22094 51492 22146
rect 50876 22092 51492 22094
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50428 21756 50708 21812
rect 50652 20690 50708 21756
rect 50652 20638 50654 20690
rect 50706 20638 50708 20690
rect 50652 20626 50708 20638
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50764 20132 50820 20142
rect 50764 20038 50820 20076
rect 50876 19346 50932 22092
rect 51436 22082 51492 22092
rect 51548 20804 51604 25566
rect 51772 25172 51828 26462
rect 52668 26516 52724 28588
rect 53228 28642 53284 28654
rect 53228 28590 53230 28642
rect 53282 28590 53284 28642
rect 53004 28084 53060 28094
rect 52780 27076 52836 27086
rect 52780 27074 52948 27076
rect 52780 27022 52782 27074
rect 52834 27022 52948 27074
rect 52780 27020 52948 27022
rect 52780 27010 52836 27020
rect 52780 26516 52836 26526
rect 52668 26514 52836 26516
rect 52668 26462 52782 26514
rect 52834 26462 52836 26514
rect 52668 26460 52836 26462
rect 52780 26450 52836 26460
rect 52332 26068 52388 26078
rect 52332 25974 52388 26012
rect 51772 25106 51828 25116
rect 52892 25506 52948 27020
rect 53004 26516 53060 28028
rect 53116 28082 53172 28094
rect 53116 28030 53118 28082
rect 53170 28030 53172 28082
rect 53116 27972 53172 28030
rect 53116 27906 53172 27916
rect 53228 27748 53284 28590
rect 53228 27682 53284 27692
rect 53676 27634 53732 27646
rect 53676 27582 53678 27634
rect 53730 27582 53732 27634
rect 53564 27300 53620 27310
rect 53228 27076 53284 27086
rect 53228 26982 53284 27020
rect 53116 26516 53172 26526
rect 53004 26514 53172 26516
rect 53004 26462 53118 26514
rect 53170 26462 53172 26514
rect 53004 26460 53172 26462
rect 53116 26450 53172 26460
rect 53564 26178 53620 27244
rect 53676 26516 53732 27582
rect 53676 26450 53732 26460
rect 53564 26126 53566 26178
rect 53618 26126 53620 26178
rect 53564 26114 53620 26126
rect 52892 25454 52894 25506
rect 52946 25454 52948 25506
rect 51996 24836 52052 24846
rect 51884 24722 51940 24734
rect 51884 24670 51886 24722
rect 51938 24670 51940 24722
rect 51772 23828 51828 23838
rect 51660 23378 51716 23390
rect 51660 23326 51662 23378
rect 51714 23326 51716 23378
rect 51660 20914 51716 23326
rect 51772 21810 51828 23772
rect 51884 23044 51940 24670
rect 51996 24050 52052 24780
rect 51996 23998 51998 24050
rect 52050 23998 52052 24050
rect 51996 23986 52052 23998
rect 52444 24724 52500 24734
rect 52444 23156 52500 24668
rect 52892 24724 52948 25454
rect 53452 25506 53508 25518
rect 53452 25454 53454 25506
rect 53506 25454 53508 25506
rect 53452 24948 53508 25454
rect 53452 24882 53508 24892
rect 52892 24050 52948 24668
rect 52892 23998 52894 24050
rect 52946 23998 52948 24050
rect 52892 23986 52948 23998
rect 53116 23940 53172 23950
rect 53004 23156 53060 23166
rect 52444 23154 52612 23156
rect 52444 23102 52446 23154
rect 52498 23102 52612 23154
rect 52444 23100 52612 23102
rect 52444 23090 52500 23100
rect 51884 22978 51940 22988
rect 52332 22932 52388 22942
rect 52332 22838 52388 22876
rect 52556 22370 52612 23100
rect 52556 22318 52558 22370
rect 52610 22318 52612 22370
rect 52556 22306 52612 22318
rect 52892 23154 53060 23156
rect 52892 23102 53006 23154
rect 53058 23102 53060 23154
rect 52892 23100 53060 23102
rect 51772 21758 51774 21810
rect 51826 21758 51828 21810
rect 51772 21746 51828 21758
rect 51884 22148 51940 22158
rect 51660 20862 51662 20914
rect 51714 20862 51716 20914
rect 51660 20850 51716 20862
rect 51436 20802 51604 20804
rect 51436 20750 51550 20802
rect 51602 20750 51604 20802
rect 51436 20748 51604 20750
rect 51436 20020 51492 20748
rect 51548 20738 51604 20748
rect 50876 19294 50878 19346
rect 50930 19294 50932 19346
rect 50876 19282 50932 19294
rect 51100 19964 51436 20020
rect 51100 19346 51156 19964
rect 51436 19954 51492 19964
rect 51100 19294 51102 19346
rect 51154 19294 51156 19346
rect 51100 19282 51156 19294
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 51548 18564 51604 18574
rect 51884 18564 51940 22092
rect 52220 22146 52276 22158
rect 52220 22094 52222 22146
rect 52274 22094 52276 22146
rect 52220 20692 52276 22094
rect 52892 21700 52948 23100
rect 53004 23090 53060 23100
rect 53116 22932 53172 23884
rect 53900 23940 53956 30156
rect 54348 28756 54404 28766
rect 54348 28084 54404 28700
rect 54348 27858 54404 28028
rect 54572 27970 54628 31052
rect 55356 31042 55412 31052
rect 55468 30324 55524 30334
rect 55468 30230 55524 30268
rect 55580 30100 55636 30110
rect 55580 29426 55636 30044
rect 55580 29374 55582 29426
rect 55634 29374 55636 29426
rect 55580 29362 55636 29374
rect 55580 28418 55636 28430
rect 55580 28366 55582 28418
rect 55634 28366 55636 28418
rect 54572 27918 54574 27970
rect 54626 27918 54628 27970
rect 54572 27906 54628 27918
rect 54908 27972 54964 27982
rect 54908 27878 54964 27916
rect 55244 27972 55300 27982
rect 55244 27878 55300 27916
rect 54348 27806 54350 27858
rect 54402 27806 54404 27858
rect 54348 27794 54404 27806
rect 55580 27636 55636 28366
rect 55692 27970 55748 31502
rect 56252 31556 56308 31566
rect 56252 31462 56308 31500
rect 56588 31556 56644 31566
rect 56812 31556 56868 33966
rect 57596 34020 57652 34030
rect 57596 33926 57652 33964
rect 57484 33236 57540 33246
rect 57036 33234 57540 33236
rect 57036 33182 57486 33234
rect 57538 33182 57540 33234
rect 57036 33180 57540 33182
rect 57036 31780 57092 33180
rect 57484 33170 57540 33180
rect 57708 32564 57764 36542
rect 58492 36370 58548 36652
rect 62524 36708 62580 37886
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 62524 36642 62580 36652
rect 61516 36596 61572 36606
rect 61516 36502 61572 36540
rect 58492 36318 58494 36370
rect 58546 36318 58548 36370
rect 58492 36306 58548 36318
rect 62524 36372 62580 36382
rect 62524 36278 62580 36316
rect 58828 35812 58884 35822
rect 58828 35718 58884 35756
rect 61404 35810 61460 35822
rect 61404 35758 61406 35810
rect 61458 35758 61460 35810
rect 60396 35588 60452 35598
rect 60396 35494 60452 35532
rect 59388 35476 59444 35486
rect 59388 35026 59444 35420
rect 61404 35140 61460 35758
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 61404 35074 61460 35084
rect 59388 34974 59390 35026
rect 59442 34974 59444 35026
rect 59388 34962 59444 34974
rect 61516 35026 61572 35038
rect 61516 34974 61518 35026
rect 61570 34974 61572 35026
rect 58828 34804 58884 34814
rect 58828 34710 58884 34748
rect 59500 34692 59556 34702
rect 59500 34598 59556 34636
rect 61516 34468 61572 34974
rect 62524 34804 62580 34814
rect 62524 34710 62580 34748
rect 61516 34402 61572 34412
rect 61404 34356 61460 34366
rect 58828 34244 58884 34254
rect 58828 34150 58884 34188
rect 61404 34242 61460 34300
rect 61404 34190 61406 34242
rect 61458 34190 61460 34242
rect 61404 34178 61460 34190
rect 60396 34018 60452 34030
rect 60396 33966 60398 34018
rect 60450 33966 60452 34018
rect 60396 33348 60452 33966
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 61516 33572 61572 33582
rect 61516 33458 61572 33516
rect 61516 33406 61518 33458
rect 61570 33406 61572 33458
rect 61516 33394 61572 33406
rect 60396 33282 60452 33292
rect 62524 33236 62580 33246
rect 62524 33142 62580 33180
rect 61404 33124 61460 33134
rect 60396 32788 60452 32798
rect 58828 32676 58884 32686
rect 58828 32582 58884 32620
rect 57708 32498 57764 32508
rect 57596 32452 57652 32462
rect 57596 32358 57652 32396
rect 60396 32450 60452 32732
rect 61404 32674 61460 33068
rect 61404 32622 61406 32674
rect 61458 32622 61460 32674
rect 61404 32610 61460 32622
rect 60396 32398 60398 32450
rect 60450 32398 60452 32450
rect 60396 32386 60452 32398
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 57036 31714 57092 31724
rect 57484 31890 57540 31902
rect 57484 31838 57486 31890
rect 57538 31838 57540 31890
rect 57036 31556 57092 31566
rect 56588 31554 57092 31556
rect 56588 31502 56590 31554
rect 56642 31502 57038 31554
rect 57090 31502 57092 31554
rect 56588 31500 57092 31502
rect 56140 31332 56196 31342
rect 56140 31218 56196 31276
rect 56140 31166 56142 31218
rect 56194 31166 56196 31218
rect 56140 31154 56196 31166
rect 56476 30996 56532 31006
rect 56588 30996 56644 31500
rect 57036 31220 57092 31500
rect 57036 31154 57092 31164
rect 57148 31444 57204 31454
rect 56476 30994 56644 30996
rect 56476 30942 56478 30994
rect 56530 30942 56644 30994
rect 56476 30940 56644 30942
rect 57148 30994 57204 31388
rect 57484 31108 57540 31838
rect 61516 31892 61572 31902
rect 61516 31798 61572 31836
rect 64316 31890 64372 31902
rect 64316 31838 64318 31890
rect 64370 31838 64372 31890
rect 58492 31668 58548 31678
rect 58492 31574 58548 31612
rect 62524 31666 62580 31678
rect 62524 31614 62526 31666
rect 62578 31614 62580 31666
rect 62524 31332 62580 31614
rect 64316 31444 64372 31838
rect 65548 31666 65604 31678
rect 65548 31614 65550 31666
rect 65602 31614 65604 31666
rect 65548 31556 65604 31614
rect 65548 31490 65604 31500
rect 64316 31378 64372 31388
rect 62524 31266 62580 31276
rect 57484 31042 57540 31052
rect 59500 31218 59556 31230
rect 59500 31166 59502 31218
rect 59554 31166 59556 31218
rect 57148 30942 57150 30994
rect 57202 30942 57204 30994
rect 55916 30324 55972 30334
rect 55916 29426 55972 30268
rect 56476 30324 56532 30940
rect 57148 30930 57204 30942
rect 57484 30660 57540 30670
rect 56532 30268 56644 30324
rect 56476 30258 56532 30268
rect 55916 29374 55918 29426
rect 55970 29374 55972 29426
rect 55916 29362 55972 29374
rect 56588 29652 56644 30268
rect 56700 29652 56756 29662
rect 57148 29652 57204 29662
rect 56588 29650 57204 29652
rect 56588 29598 56702 29650
rect 56754 29598 57150 29650
rect 57202 29598 57204 29650
rect 56588 29596 57204 29598
rect 56588 28754 56644 29596
rect 56700 29586 56756 29596
rect 57148 29586 57204 29596
rect 56588 28702 56590 28754
rect 56642 28702 56644 28754
rect 55692 27918 55694 27970
rect 55746 27918 55748 27970
rect 55692 27906 55748 27918
rect 56028 28644 56084 28654
rect 56028 27972 56084 28588
rect 56252 28420 56308 28430
rect 56252 28418 56420 28420
rect 56252 28366 56254 28418
rect 56306 28366 56420 28418
rect 56252 28364 56420 28366
rect 56252 28354 56308 28364
rect 56028 27878 56084 27916
rect 56252 27972 56308 27982
rect 55580 27570 55636 27580
rect 56252 27298 56308 27916
rect 56252 27246 56254 27298
rect 56306 27246 56308 27298
rect 56252 27234 56308 27246
rect 55468 26850 55524 26862
rect 55468 26798 55470 26850
rect 55522 26798 55524 26850
rect 55468 26514 55524 26798
rect 56364 26740 56420 28364
rect 56588 28084 56644 28702
rect 57484 28754 57540 30604
rect 57596 29540 57652 29550
rect 57596 29314 57652 29484
rect 57596 29262 57598 29314
rect 57650 29262 57652 29314
rect 57596 29250 57652 29262
rect 58828 29538 58884 29550
rect 58828 29486 58830 29538
rect 58882 29486 58884 29538
rect 58828 29092 58884 29486
rect 58828 29026 58884 29036
rect 57484 28702 57486 28754
rect 57538 28702 57540 28754
rect 57484 28690 57540 28702
rect 59500 28754 59556 31166
rect 60508 31220 60564 31230
rect 60508 31126 60564 31164
rect 62412 31106 62468 31118
rect 62412 31054 62414 31106
rect 62466 31054 62468 31106
rect 60172 30996 60228 31006
rect 60172 30902 60228 30940
rect 61404 30882 61460 30894
rect 61404 30830 61406 30882
rect 61458 30830 61460 30882
rect 61404 30100 61460 30830
rect 61516 30884 61572 30894
rect 61516 30322 61572 30828
rect 62412 30772 62468 31054
rect 64988 30996 65044 31006
rect 64988 30902 65044 30940
rect 66108 30996 66164 31006
rect 66108 30902 66164 30940
rect 62412 30706 62468 30716
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 61516 30270 61518 30322
rect 61570 30270 61572 30322
rect 61516 30258 61572 30270
rect 61404 30034 61460 30044
rect 62524 30098 62580 30110
rect 62524 30046 62526 30098
rect 62578 30046 62580 30098
rect 61516 29876 61572 29886
rect 61404 29538 61460 29550
rect 61404 29486 61406 29538
rect 61458 29486 61460 29538
rect 60396 29316 60452 29326
rect 60396 29222 60452 29260
rect 61404 28868 61460 29486
rect 61404 28802 61460 28812
rect 59500 28702 59502 28754
rect 59554 28702 59556 28754
rect 59500 28690 59556 28702
rect 61516 28754 61572 29820
rect 62524 28980 62580 30046
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 62524 28914 62580 28924
rect 61516 28702 61518 28754
rect 61570 28702 61572 28754
rect 61516 28690 61572 28702
rect 59276 28644 59332 28654
rect 59276 28550 59332 28588
rect 57596 28532 57652 28542
rect 56700 28084 56756 28094
rect 56588 28082 56756 28084
rect 56588 28030 56702 28082
rect 56754 28030 56756 28082
rect 56588 28028 56756 28030
rect 56700 28018 56756 28028
rect 57596 27746 57652 28476
rect 58492 28530 58548 28542
rect 58492 28478 58494 28530
rect 58546 28478 58548 28530
rect 58492 27860 58548 28478
rect 62524 28532 62580 28542
rect 62524 28438 62580 28476
rect 58492 27794 58548 27804
rect 58940 27970 58996 27982
rect 58940 27918 58942 27970
rect 58994 27918 58996 27970
rect 57596 27694 57598 27746
rect 57650 27694 57652 27746
rect 57596 27682 57652 27694
rect 57484 27188 57540 27198
rect 57484 27094 57540 27132
rect 58492 26962 58548 26974
rect 58492 26910 58494 26962
rect 58546 26910 58548 26962
rect 58492 26852 58548 26910
rect 58492 26786 58548 26796
rect 56364 26674 56420 26684
rect 55468 26462 55470 26514
rect 55522 26462 55524 26514
rect 55468 26450 55524 26462
rect 54572 26404 54628 26414
rect 54572 26310 54628 26348
rect 58828 26404 58884 26414
rect 58828 26310 58884 26348
rect 55356 26178 55412 26190
rect 55356 26126 55358 26178
rect 55410 26126 55412 26178
rect 55132 25172 55188 25182
rect 53900 23874 53956 23884
rect 54348 24946 54404 24958
rect 54348 24894 54350 24946
rect 54402 24894 54404 24946
rect 53004 22876 53172 22932
rect 53004 21810 53060 22876
rect 53676 22708 53732 22718
rect 53004 21758 53006 21810
rect 53058 21758 53060 21810
rect 53004 21746 53060 21758
rect 53228 22370 53284 22382
rect 53228 22318 53230 22370
rect 53282 22318 53284 22370
rect 52892 21634 52948 21644
rect 53228 21476 53284 22318
rect 53676 21476 53732 22652
rect 54348 22596 54404 24894
rect 55132 24834 55188 25116
rect 55132 24782 55134 24834
rect 55186 24782 55188 24834
rect 55132 24770 55188 24782
rect 55356 24836 55412 26126
rect 57596 26180 57652 26190
rect 57596 26086 57652 26124
rect 57708 25618 57764 25630
rect 57708 25566 57710 25618
rect 57762 25566 57764 25618
rect 57596 25396 57652 25406
rect 55916 25284 55972 25294
rect 55916 25190 55972 25228
rect 56476 25282 56532 25294
rect 56476 25230 56478 25282
rect 56530 25230 56532 25282
rect 56476 24836 56532 25230
rect 55356 24780 55524 24836
rect 55468 24610 55524 24780
rect 56476 24770 56532 24780
rect 55468 24558 55470 24610
rect 55522 24558 55524 24610
rect 54908 24500 54964 24510
rect 54908 24406 54964 24444
rect 55468 24052 55524 24558
rect 57596 24610 57652 25340
rect 57596 24558 57598 24610
rect 57650 24558 57652 24610
rect 57596 24546 57652 24558
rect 57708 24276 57764 25566
rect 58716 25620 58772 25630
rect 58772 25564 58884 25620
rect 58716 25554 58772 25564
rect 58828 25394 58884 25564
rect 58940 25508 58996 27918
rect 61404 27972 61460 27982
rect 61404 27878 61460 27916
rect 60396 27748 60452 27758
rect 60396 27654 60452 27692
rect 59276 27636 59332 27646
rect 59276 27186 59332 27580
rect 65916 27468 66180 27478
rect 59276 27134 59278 27186
rect 59330 27134 59332 27186
rect 59276 27122 59332 27134
rect 60284 27412 60340 27422
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 58940 25442 58996 25452
rect 59500 27074 59556 27086
rect 59500 27022 59502 27074
rect 59554 27022 59556 27074
rect 59500 25618 59556 27022
rect 60284 26180 60340 27356
rect 61516 27186 61572 27198
rect 61516 27134 61518 27186
rect 61570 27134 61572 27186
rect 61516 27076 61572 27134
rect 61516 27010 61572 27020
rect 62524 26962 62580 26974
rect 62524 26910 62526 26962
rect 62578 26910 62580 26962
rect 61404 26740 61460 26750
rect 61404 26402 61460 26684
rect 61404 26350 61406 26402
rect 61458 26350 61460 26402
rect 61404 26338 61460 26350
rect 60396 26180 60452 26190
rect 60284 26178 60452 26180
rect 60284 26126 60398 26178
rect 60450 26126 60452 26178
rect 60284 26124 60452 26126
rect 60396 26114 60452 26124
rect 62524 26068 62580 26910
rect 62524 26002 62580 26012
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 59500 25566 59502 25618
rect 59554 25566 59556 25618
rect 58828 25342 58830 25394
rect 58882 25342 58884 25394
rect 58828 25330 58884 25342
rect 58828 24836 58884 24846
rect 58828 24742 58884 24780
rect 57708 24210 57764 24220
rect 55468 23986 55524 23996
rect 55916 24052 55972 24062
rect 55356 23268 55412 23278
rect 54348 22530 54404 22540
rect 54908 23266 55412 23268
rect 54908 23214 55358 23266
rect 55410 23214 55412 23266
rect 54908 23212 55412 23214
rect 53900 22260 53956 22270
rect 53788 21476 53844 21486
rect 53676 21474 53844 21476
rect 53676 21422 53790 21474
rect 53842 21422 53844 21474
rect 53676 21420 53844 21422
rect 53228 21410 53284 21420
rect 53788 21410 53844 21420
rect 52220 20626 52276 20636
rect 52556 21362 52612 21374
rect 52556 21310 52558 21362
rect 52610 21310 52612 21362
rect 52556 20188 52612 21310
rect 53676 21252 53732 21262
rect 53676 20914 53732 21196
rect 53676 20862 53678 20914
rect 53730 20862 53732 20914
rect 53676 20850 53732 20862
rect 52556 20132 52724 20188
rect 52556 19908 52612 19918
rect 52556 19814 52612 19852
rect 52668 19124 52724 20132
rect 53900 20130 53956 22204
rect 53900 20078 53902 20130
rect 53954 20078 53956 20130
rect 53900 20066 53956 20078
rect 54012 21700 54068 21710
rect 54012 19346 54068 21644
rect 54796 21698 54852 21710
rect 54796 21646 54798 21698
rect 54850 21646 54852 21698
rect 54796 21028 54852 21646
rect 54796 20962 54852 20972
rect 54684 20692 54740 20702
rect 54684 20598 54740 20636
rect 54908 20188 54964 23212
rect 55356 23202 55412 23212
rect 55580 22596 55636 22606
rect 55580 21698 55636 22540
rect 55692 22260 55748 22270
rect 55692 22146 55748 22204
rect 55692 22094 55694 22146
rect 55746 22094 55748 22146
rect 55692 22082 55748 22094
rect 55580 21646 55582 21698
rect 55634 21646 55636 21698
rect 55580 21634 55636 21646
rect 55916 21698 55972 23996
rect 58604 24052 58660 24062
rect 58604 23958 58660 23996
rect 59500 24052 59556 25566
rect 59612 25284 59668 25294
rect 59612 25190 59668 25228
rect 60396 24948 60452 24958
rect 60396 24610 60452 24892
rect 60396 24558 60398 24610
rect 60450 24558 60452 24610
rect 60396 24546 60452 24558
rect 61404 24834 61460 24846
rect 61404 24782 61406 24834
rect 61458 24782 61460 24834
rect 61404 24500 61460 24782
rect 61404 24434 61460 24444
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 56476 23940 56532 23950
rect 56476 23846 56532 23884
rect 58268 23828 58324 23838
rect 58268 23734 58324 23772
rect 56252 23268 56308 23278
rect 55916 21646 55918 21698
rect 55970 21646 55972 21698
rect 54684 20132 54964 20188
rect 55916 20132 55972 21646
rect 56140 22930 56196 22942
rect 56140 22878 56142 22930
rect 56194 22878 56196 22930
rect 56140 21700 56196 22878
rect 56252 22594 56308 23212
rect 58828 23268 58884 23278
rect 58828 23174 58884 23212
rect 59500 23154 59556 23996
rect 59500 23102 59502 23154
rect 59554 23102 59556 23154
rect 59500 23090 59556 23102
rect 57596 23044 57652 23054
rect 57596 22950 57652 22988
rect 59612 23042 59668 23054
rect 59612 22990 59614 23042
rect 59666 22990 59668 23042
rect 56252 22542 56254 22594
rect 56306 22542 56308 22594
rect 56252 22530 56308 22542
rect 58492 22932 58548 22942
rect 57484 22484 57540 22494
rect 57484 22390 57540 22428
rect 58492 22258 58548 22876
rect 58492 22206 58494 22258
rect 58546 22206 58548 22258
rect 58492 22194 58548 22206
rect 59612 22260 59668 22990
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 59612 22194 59668 22204
rect 56140 21634 56196 21644
rect 58828 21700 58884 21710
rect 58828 21606 58884 21644
rect 57596 21476 57652 21486
rect 57596 21382 57652 21420
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 54684 20130 54740 20132
rect 54684 20078 54686 20130
rect 54738 20078 54740 20130
rect 54684 20066 54740 20078
rect 55916 20066 55972 20076
rect 54460 20020 54516 20030
rect 54460 19926 54516 19964
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 54012 19294 54014 19346
rect 54066 19294 54068 19346
rect 54012 19282 54068 19294
rect 52668 19058 52724 19068
rect 55020 19124 55076 19134
rect 55020 19030 55076 19068
rect 51548 18562 51940 18564
rect 51548 18510 51550 18562
rect 51602 18510 51940 18562
rect 51548 18508 51940 18510
rect 51548 18498 51604 18508
rect 50204 18286 50206 18338
rect 50258 18286 50260 18338
rect 50204 18274 50260 18286
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 48636 17780 48692 17790
rect 48524 17778 48692 17780
rect 48524 17726 48638 17778
rect 48690 17726 48692 17778
rect 48524 17724 48692 17726
rect 48636 17714 48692 17724
rect 47068 17502 47070 17554
rect 47122 17502 47124 17554
rect 47068 17490 47124 17502
rect 49644 17556 49700 17566
rect 49644 17462 49700 17500
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 46060 16994 46228 16996
rect 46060 16942 46062 16994
rect 46114 16942 46228 16994
rect 46060 16940 46228 16942
rect 46060 16930 46116 16940
rect 44716 16718 44718 16770
rect 44770 16718 44772 16770
rect 44716 16706 44772 16718
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 42588 16158 42590 16210
rect 42642 16158 42644 16210
rect 42588 16146 42644 16158
rect 41692 15922 41748 15932
rect 43708 15988 43764 15998
rect 43708 15894 43764 15932
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 36764 15374 36766 15426
rect 36818 15374 36820 15426
rect 36764 15362 36820 15374
rect 35756 15150 35758 15202
rect 35810 15150 35812 15202
rect 35756 15138 35812 15150
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 31276 14366 31278 14418
rect 31330 14366 31332 14418
rect 31276 14354 31332 14366
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 40572 3332 40628 3342
rect 41244 3332 41300 3342
rect 43932 3332 43988 3342
rect 44604 3332 44660 3342
rect 48636 3332 48692 3342
rect 55020 3332 55076 3342
rect 40348 3330 40628 3332
rect 40348 3278 40574 3330
rect 40626 3278 40628 3330
rect 40348 3276 40628 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 40348 800 40404 3276
rect 40572 3266 40628 3276
rect 41020 3330 41300 3332
rect 41020 3278 41246 3330
rect 41298 3278 41300 3330
rect 41020 3276 41300 3278
rect 41020 800 41076 3276
rect 41244 3266 41300 3276
rect 43708 3330 43988 3332
rect 43708 3278 43934 3330
rect 43986 3278 43988 3330
rect 43708 3276 43988 3278
rect 43708 800 43764 3276
rect 43932 3266 43988 3276
rect 44380 3330 44660 3332
rect 44380 3278 44606 3330
rect 44658 3278 44660 3330
rect 44380 3276 44660 3278
rect 44380 800 44436 3276
rect 44604 3266 44660 3276
rect 48412 3330 48692 3332
rect 48412 3278 48638 3330
rect 48690 3278 48692 3330
rect 48412 3276 48692 3278
rect 48412 800 48468 3276
rect 48636 3266 48692 3276
rect 54460 3330 55076 3332
rect 54460 3278 55022 3330
rect 55074 3278 55076 3330
rect 54460 3276 55076 3278
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 54460 800 54516 3276
rect 55020 3266 55076 3276
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 40320 0 40432 800
rect 40992 0 41104 800
rect 43680 0 43792 800
rect 44352 0 44464 800
rect 48384 0 48496 800
rect 54432 0 54544 800
<< via2 >>
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 66220 62524 66276 62580
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 41468 54348 41524 54404
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 28588 53788 28644 53844
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 10892 47628 10948 47684
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 10780 40572 10836 40628
rect 9996 40348 10052 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 9100 39730 9156 39732
rect 9100 39678 9102 39730
rect 9102 39678 9154 39730
rect 9154 39678 9156 39730
rect 9100 39676 9156 39678
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 7980 38332 8036 38388
rect 6972 38108 7028 38164
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 2044 35868 2100 35924
rect 3052 35644 3108 35700
rect 3052 34860 3108 34916
rect 3836 33292 3892 33348
rect 3052 33068 3108 33124
rect 3052 31666 3108 31668
rect 3052 31614 3054 31666
rect 3054 31614 3106 31666
rect 3106 31614 3108 31666
rect 3052 31612 3108 31614
rect 4172 35810 4228 35812
rect 4172 35758 4174 35810
rect 4174 35758 4226 35810
rect 4226 35758 4228 35810
rect 4172 35756 4228 35758
rect 4172 34076 4228 34132
rect 6972 37378 7028 37380
rect 6972 37326 6974 37378
rect 6974 37326 7026 37378
rect 7026 37326 7028 37378
rect 6972 37324 7028 37326
rect 5180 37212 5236 37268
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 7084 36652 7140 36708
rect 10780 39340 10836 39396
rect 9884 38332 9940 38388
rect 8092 37772 8148 37828
rect 8652 37212 8708 37268
rect 7980 37154 8036 37156
rect 7980 37102 7982 37154
rect 7982 37102 8034 37154
rect 8034 37102 8036 37154
rect 7980 37100 8036 37102
rect 8092 36594 8148 36596
rect 8092 36542 8094 36594
rect 8094 36542 8146 36594
rect 8146 36542 8148 36594
rect 8092 36540 8148 36542
rect 7980 36428 8036 36484
rect 7084 36092 7140 36148
rect 6972 35420 7028 35476
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 5180 35308 5236 35364
rect 4684 35252 4740 35254
rect 7308 35026 7364 35028
rect 7308 34974 7310 35026
rect 7310 34974 7362 35026
rect 7362 34974 7364 35026
rect 7308 34972 7364 34974
rect 6300 34802 6356 34804
rect 6300 34750 6302 34802
rect 6302 34750 6354 34802
rect 6354 34750 6356 34802
rect 6300 34748 6356 34750
rect 9324 37212 9380 37268
rect 10220 36764 10276 36820
rect 9884 36482 9940 36484
rect 9884 36430 9886 36482
rect 9886 36430 9938 36482
rect 9938 36430 9940 36482
rect 9884 36428 9940 36430
rect 17164 47180 17220 47236
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20300 48524 20356 48580
rect 19740 48076 19796 48132
rect 18508 47180 18564 47236
rect 17164 45612 17220 45668
rect 16940 44828 16996 44884
rect 11676 40626 11732 40628
rect 11676 40574 11678 40626
rect 11678 40574 11730 40626
rect 11730 40574 11732 40626
rect 11676 40572 11732 40574
rect 12012 40572 12068 40628
rect 12236 40348 12292 40404
rect 11900 39900 11956 39956
rect 11900 39564 11956 39620
rect 12012 39004 12068 39060
rect 11004 38946 11060 38948
rect 11004 38894 11006 38946
rect 11006 38894 11058 38946
rect 11058 38894 11060 38946
rect 11004 38892 11060 38894
rect 13916 39900 13972 39956
rect 13020 38780 13076 38836
rect 13804 38834 13860 38836
rect 13804 38782 13806 38834
rect 13806 38782 13858 38834
rect 13858 38782 13860 38834
rect 13804 38780 13860 38782
rect 13468 38668 13524 38724
rect 12908 38108 12964 38164
rect 11004 37436 11060 37492
rect 11900 37324 11956 37380
rect 10892 36204 10948 36260
rect 11116 36652 11172 36708
rect 9884 35532 9940 35588
rect 7980 34300 8036 34356
rect 6972 34242 7028 34244
rect 6972 34190 6974 34242
rect 6974 34190 7026 34242
rect 7026 34190 7028 34242
rect 6972 34188 7028 34190
rect 9100 34076 9156 34132
rect 7980 34018 8036 34020
rect 7980 33966 7982 34018
rect 7982 33966 8034 34018
rect 8034 33966 8036 34018
rect 7980 33964 8036 33966
rect 5180 33852 5236 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 7868 33740 7924 33796
rect 4284 33516 4340 33572
rect 4060 33458 4116 33460
rect 4060 33406 4062 33458
rect 4062 33406 4114 33458
rect 4114 33406 4116 33458
rect 4060 33404 4116 33406
rect 8316 33516 8372 33572
rect 4172 32956 4228 33012
rect 6636 32732 6692 32788
rect 6972 32674 7028 32676
rect 6972 32622 6974 32674
rect 6974 32622 7026 32674
rect 7026 32622 7028 32674
rect 6972 32620 7028 32622
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 5180 32172 5236 32228
rect 4684 32116 4740 32118
rect 4060 31890 4116 31892
rect 4060 31838 4062 31890
rect 4062 31838 4114 31890
rect 4114 31838 4116 31890
rect 4060 31836 4116 31838
rect 3948 31500 4004 31556
rect 5292 31612 5348 31668
rect 2156 31106 2212 31108
rect 2156 31054 2158 31106
rect 2158 31054 2210 31106
rect 2210 31054 2212 31106
rect 2156 31052 2212 31054
rect 3164 30882 3220 30884
rect 3164 30830 3166 30882
rect 3166 30830 3218 30882
rect 3218 30830 3220 30882
rect 3164 30828 3220 30830
rect 2828 30716 2884 30772
rect 2044 28588 2100 28644
rect 1820 26236 1876 26292
rect 1708 24892 1764 24948
rect 2716 24780 2772 24836
rect 4396 30770 4452 30772
rect 4396 30718 4398 30770
rect 4398 30718 4450 30770
rect 4450 30718 4452 30770
rect 4396 30716 4452 30718
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5068 30380 5124 30436
rect 4060 30156 4116 30212
rect 3052 30098 3108 30100
rect 3052 30046 3054 30098
rect 3054 30046 3106 30098
rect 3106 30046 3108 30098
rect 3052 30044 3108 30046
rect 4508 30044 4564 30100
rect 3164 29708 3220 29764
rect 4172 29148 4228 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4508 28812 4564 28868
rect 3052 28530 3108 28532
rect 3052 28478 3054 28530
rect 3054 28478 3106 28530
rect 3106 28478 3108 28530
rect 3052 28476 3108 28478
rect 3948 28252 4004 28308
rect 3052 27580 3108 27636
rect 3500 27244 3556 27300
rect 7084 31666 7140 31668
rect 7084 31614 7086 31666
rect 7086 31614 7138 31666
rect 7138 31614 7140 31666
rect 7084 31612 7140 31614
rect 7084 30604 7140 30660
rect 5292 29260 5348 29316
rect 5180 28700 5236 28756
rect 6188 29538 6244 29540
rect 6188 29486 6190 29538
rect 6190 29486 6242 29538
rect 6242 29486 6244 29538
rect 6188 29484 6244 29486
rect 6076 29036 6132 29092
rect 6860 28754 6916 28756
rect 6860 28702 6862 28754
rect 6862 28702 6914 28754
rect 6914 28702 6916 28754
rect 6860 28700 6916 28702
rect 5404 28588 5460 28644
rect 6524 28642 6580 28644
rect 6524 28590 6526 28642
rect 6526 28590 6578 28642
rect 6578 28590 6580 28642
rect 6524 28588 6580 28590
rect 7196 28642 7252 28644
rect 7196 28590 7198 28642
rect 7198 28590 7250 28642
rect 7250 28590 7252 28642
rect 7196 28588 7252 28590
rect 4508 28476 4564 28532
rect 6412 28418 6468 28420
rect 6412 28366 6414 28418
rect 6414 28366 6466 28418
rect 6466 28366 6468 28418
rect 6412 28364 6468 28366
rect 7420 28364 7476 28420
rect 4732 28082 4788 28084
rect 4732 28030 4734 28082
rect 4734 28030 4786 28082
rect 4786 28030 4788 28082
rect 4732 28028 4788 28030
rect 4060 27804 4116 27860
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4060 27132 4116 27188
rect 3948 26460 4004 26516
rect 2940 26012 2996 26068
rect 3836 25228 3892 25284
rect 3052 23826 3108 23828
rect 3052 23774 3054 23826
rect 3054 23774 3106 23826
rect 3106 23774 3108 23826
rect 3052 23772 3108 23774
rect 3052 23548 3108 23604
rect 4508 26290 4564 26292
rect 4508 26238 4510 26290
rect 4510 26238 4562 26290
rect 4562 26238 4564 26290
rect 4508 26236 4564 26238
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4060 25004 4116 25060
rect 5068 25004 5124 25060
rect 4732 24946 4788 24948
rect 4732 24894 4734 24946
rect 4734 24894 4786 24946
rect 4786 24894 4788 24946
rect 4732 24892 4788 24894
rect 5964 27858 6020 27860
rect 5964 27806 5966 27858
rect 5966 27806 6018 27858
rect 6018 27806 6020 27858
rect 5964 27804 6020 27806
rect 6636 27468 6692 27524
rect 5740 26962 5796 26964
rect 5740 26910 5742 26962
rect 5742 26910 5794 26962
rect 5794 26910 5796 26962
rect 5740 26908 5796 26910
rect 5404 26236 5460 26292
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5068 24050 5124 24052
rect 5068 23998 5070 24050
rect 5070 23998 5122 24050
rect 5122 23998 5124 24050
rect 5068 23996 5124 23998
rect 4172 23100 4228 23156
rect 4060 22204 4116 22260
rect 3164 21420 3220 21476
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4844 21756 4900 21812
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5964 26236 6020 26292
rect 6524 26236 6580 26292
rect 5292 23548 5348 23604
rect 5404 23996 5460 24052
rect 5964 23154 6020 23156
rect 5964 23102 5966 23154
rect 5966 23102 6018 23154
rect 6018 23102 6020 23154
rect 5964 23100 6020 23102
rect 5852 22204 5908 22260
rect 6188 24892 6244 24948
rect 7196 26962 7252 26964
rect 7196 26910 7198 26962
rect 7198 26910 7250 26962
rect 7250 26910 7252 26962
rect 7196 26908 7252 26910
rect 8204 30716 8260 30772
rect 7868 29484 7924 29540
rect 11228 35644 11284 35700
rect 9100 32562 9156 32564
rect 9100 32510 9102 32562
rect 9102 32510 9154 32562
rect 9154 32510 9156 32562
rect 9100 32508 9156 32510
rect 9884 32562 9940 32564
rect 9884 32510 9886 32562
rect 9886 32510 9938 32562
rect 9938 32510 9940 32562
rect 9884 32508 9940 32510
rect 9212 32284 9268 32340
rect 9100 31890 9156 31892
rect 9100 31838 9102 31890
rect 9102 31838 9154 31890
rect 9154 31838 9156 31890
rect 9100 31836 9156 31838
rect 8204 29596 8260 29652
rect 8092 29372 8148 29428
rect 9436 31836 9492 31892
rect 9996 31836 10052 31892
rect 9884 31500 9940 31556
rect 9884 30828 9940 30884
rect 8988 30268 9044 30324
rect 9884 30044 9940 30100
rect 7644 28642 7700 28644
rect 7644 28590 7646 28642
rect 7646 28590 7698 28642
rect 7698 28590 7700 28642
rect 7644 28588 7700 28590
rect 8428 28028 8484 28084
rect 8316 27970 8372 27972
rect 8316 27918 8318 27970
rect 8318 27918 8370 27970
rect 8370 27918 8372 27970
rect 8316 27916 8372 27918
rect 8092 27580 8148 27636
rect 8316 26796 8372 26852
rect 7532 25676 7588 25732
rect 6748 23826 6804 23828
rect 6748 23774 6750 23826
rect 6750 23774 6802 23826
rect 6802 23774 6804 23826
rect 6748 23772 6804 23774
rect 5964 21756 6020 21812
rect 5628 21586 5684 21588
rect 5628 21534 5630 21586
rect 5630 21534 5682 21586
rect 5682 21534 5684 21586
rect 5628 21532 5684 21534
rect 5180 20188 5236 20244
rect 2268 19292 2324 19348
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 7756 25618 7812 25620
rect 7756 25566 7758 25618
rect 7758 25566 7810 25618
rect 7810 25566 7812 25618
rect 7756 25564 7812 25566
rect 7644 21868 7700 21924
rect 7868 21980 7924 22036
rect 7756 21644 7812 21700
rect 6636 19964 6692 20020
rect 7196 18396 7252 18452
rect 8764 29372 8820 29428
rect 8652 26460 8708 26516
rect 8764 28588 8820 28644
rect 10556 33516 10612 33572
rect 10668 32338 10724 32340
rect 10668 32286 10670 32338
rect 10670 32286 10722 32338
rect 10722 32286 10724 32338
rect 10668 32284 10724 32286
rect 12012 37154 12068 37156
rect 12012 37102 12014 37154
rect 12014 37102 12066 37154
rect 12066 37102 12068 37154
rect 12012 37100 12068 37102
rect 12460 36652 12516 36708
rect 12796 36764 12852 36820
rect 13020 37826 13076 37828
rect 13020 37774 13022 37826
rect 13022 37774 13074 37826
rect 13074 37774 13076 37826
rect 13020 37772 13076 37774
rect 13244 37266 13300 37268
rect 13244 37214 13246 37266
rect 13246 37214 13298 37266
rect 13298 37214 13300 37266
rect 13244 37212 13300 37214
rect 12460 36316 12516 36372
rect 12684 35980 12740 36036
rect 11452 35532 11508 35588
rect 12796 35756 12852 35812
rect 12236 34914 12292 34916
rect 12236 34862 12238 34914
rect 12238 34862 12290 34914
rect 12290 34862 12292 34914
rect 12236 34860 12292 34862
rect 11676 34690 11732 34692
rect 11676 34638 11678 34690
rect 11678 34638 11730 34690
rect 11730 34638 11732 34690
rect 11676 34636 11732 34638
rect 11340 33516 11396 33572
rect 12124 33346 12180 33348
rect 12124 33294 12126 33346
rect 12126 33294 12178 33346
rect 12178 33294 12180 33346
rect 12124 33292 12180 33294
rect 11340 31164 11396 31220
rect 12012 31836 12068 31892
rect 10220 30268 10276 30324
rect 13020 35308 13076 35364
rect 14812 43650 14868 43652
rect 14812 43598 14814 43650
rect 14814 43598 14866 43650
rect 14866 43598 14868 43650
rect 14812 43596 14868 43598
rect 15932 42642 15988 42644
rect 15932 42590 15934 42642
rect 15934 42590 15986 42642
rect 15986 42590 15988 42642
rect 15932 42588 15988 42590
rect 17836 46508 17892 46564
rect 17500 44828 17556 44884
rect 16156 42028 16212 42084
rect 15820 41916 15876 41972
rect 14700 39676 14756 39732
rect 15932 41074 15988 41076
rect 15932 41022 15934 41074
rect 15934 41022 15986 41074
rect 15986 41022 15988 41074
rect 15932 41020 15988 41022
rect 16268 40348 16324 40404
rect 15148 38668 15204 38724
rect 15820 38668 15876 38724
rect 15036 38556 15092 38612
rect 13916 36988 13972 37044
rect 13692 36370 13748 36372
rect 13692 36318 13694 36370
rect 13694 36318 13746 36370
rect 13746 36318 13748 36370
rect 13692 36316 13748 36318
rect 14028 36764 14084 36820
rect 14812 36764 14868 36820
rect 14588 35980 14644 36036
rect 14812 35756 14868 35812
rect 16604 40460 16660 40516
rect 16268 37212 16324 37268
rect 15820 36652 15876 36708
rect 16044 35756 16100 35812
rect 16828 41580 16884 41636
rect 16940 42028 16996 42084
rect 16716 39900 16772 39956
rect 16828 39676 16884 39732
rect 18844 46562 18900 46564
rect 18844 46510 18846 46562
rect 18846 46510 18898 46562
rect 18898 46510 18900 46562
rect 18844 46508 18900 46510
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19628 46396 19684 46452
rect 19516 46060 19572 46116
rect 20860 46956 20916 47012
rect 20860 45890 20916 45892
rect 20860 45838 20862 45890
rect 20862 45838 20914 45890
rect 20914 45838 20916 45890
rect 20860 45836 20916 45838
rect 18620 45612 18676 45668
rect 20300 45612 20356 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 17836 42082 17892 42084
rect 17836 42030 17838 42082
rect 17838 42030 17890 42082
rect 17890 42030 17892 42082
rect 17836 42028 17892 42030
rect 17724 41580 17780 41636
rect 17276 40572 17332 40628
rect 17164 38668 17220 38724
rect 17500 40402 17556 40404
rect 17500 40350 17502 40402
rect 17502 40350 17554 40402
rect 17554 40350 17556 40402
rect 17500 40348 17556 40350
rect 17836 40514 17892 40516
rect 17836 40462 17838 40514
rect 17838 40462 17890 40514
rect 17890 40462 17892 40514
rect 17836 40460 17892 40462
rect 17724 40348 17780 40404
rect 17724 39618 17780 39620
rect 17724 39566 17726 39618
rect 17726 39566 17778 39618
rect 17778 39566 17780 39618
rect 17724 39564 17780 39566
rect 17052 36092 17108 36148
rect 16716 35756 16772 35812
rect 15148 35420 15204 35476
rect 15260 34860 15316 34916
rect 13468 34636 13524 34692
rect 14140 34130 14196 34132
rect 14140 34078 14142 34130
rect 14142 34078 14194 34130
rect 14194 34078 14196 34130
rect 14140 34076 14196 34078
rect 13580 33964 13636 34020
rect 12460 31836 12516 31892
rect 14700 33964 14756 34020
rect 13804 33516 13860 33572
rect 13580 31836 13636 31892
rect 13692 33404 13748 33460
rect 12012 30940 12068 30996
rect 11340 30210 11396 30212
rect 11340 30158 11342 30210
rect 11342 30158 11394 30210
rect 11394 30158 11396 30210
rect 11340 30156 11396 30158
rect 13132 31218 13188 31220
rect 13132 31166 13134 31218
rect 13134 31166 13186 31218
rect 13186 31166 13188 31218
rect 13132 31164 13188 31166
rect 13244 30994 13300 30996
rect 13244 30942 13246 30994
rect 13246 30942 13298 30994
rect 13298 30942 13300 30994
rect 13244 30940 13300 30942
rect 13916 30604 13972 30660
rect 15820 34018 15876 34020
rect 15820 33966 15822 34018
rect 15822 33966 15874 34018
rect 15874 33966 15876 34018
rect 15820 33964 15876 33966
rect 14700 30940 14756 30996
rect 14700 30322 14756 30324
rect 14700 30270 14702 30322
rect 14702 30270 14754 30322
rect 14754 30270 14756 30322
rect 14700 30268 14756 30270
rect 15036 33516 15092 33572
rect 16492 35308 16548 35364
rect 17388 37212 17444 37268
rect 19516 44994 19572 44996
rect 19516 44942 19518 44994
rect 19518 44942 19570 44994
rect 19570 44942 19572 44994
rect 19516 44940 19572 44942
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 18396 42924 18452 42980
rect 18732 41804 18788 41860
rect 18732 41580 18788 41636
rect 18396 38668 18452 38724
rect 18172 36482 18228 36484
rect 18172 36430 18174 36482
rect 18174 36430 18226 36482
rect 18226 36430 18228 36482
rect 18172 36428 18228 36430
rect 18844 38220 18900 38276
rect 19404 38332 19460 38388
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 22316 48524 22372 48580
rect 21308 48076 21364 48132
rect 21644 47346 21700 47348
rect 21644 47294 21646 47346
rect 21646 47294 21698 47346
rect 21698 47294 21700 47346
rect 21644 47292 21700 47294
rect 21308 46060 21364 46116
rect 21420 45890 21476 45892
rect 21420 45838 21422 45890
rect 21422 45838 21474 45890
rect 21474 45838 21476 45890
rect 21420 45836 21476 45838
rect 21756 46956 21812 47012
rect 22428 47346 22484 47348
rect 22428 47294 22430 47346
rect 22430 47294 22482 47346
rect 22482 47294 22484 47346
rect 22428 47292 22484 47294
rect 21980 46172 22036 46228
rect 22876 47068 22932 47124
rect 22652 46060 22708 46116
rect 22540 45612 22596 45668
rect 23884 48076 23940 48132
rect 23660 46956 23716 47012
rect 23772 47068 23828 47124
rect 23772 46284 23828 46340
rect 23660 46172 23716 46228
rect 23548 45612 23604 45668
rect 21644 44828 21700 44884
rect 23660 44828 23716 44884
rect 20860 43596 20916 43652
rect 20636 41970 20692 41972
rect 20636 41918 20638 41970
rect 20638 41918 20690 41970
rect 20690 41918 20692 41970
rect 20636 41916 20692 41918
rect 19740 41298 19796 41300
rect 19740 41246 19742 41298
rect 19742 41246 19794 41298
rect 19794 41246 19796 41298
rect 19740 41244 19796 41246
rect 20748 40962 20804 40964
rect 20748 40910 20750 40962
rect 20750 40910 20802 40962
rect 20802 40910 20804 40962
rect 20748 40908 20804 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19852 40290 19908 40292
rect 19852 40238 19854 40290
rect 19854 40238 19906 40290
rect 19906 40238 19908 40290
rect 19852 40236 19908 40238
rect 20188 39452 20244 39508
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 21196 42978 21252 42980
rect 21196 42926 21198 42978
rect 21198 42926 21250 42978
rect 21250 42926 21252 42978
rect 21196 42924 21252 42926
rect 21532 41916 21588 41972
rect 21756 42028 21812 42084
rect 20972 41804 21028 41860
rect 21084 41020 21140 41076
rect 23100 42812 23156 42868
rect 22092 42252 22148 42308
rect 21980 41244 22036 41300
rect 22876 40572 22932 40628
rect 20972 39340 21028 39396
rect 21756 40124 21812 40180
rect 22316 40460 22372 40516
rect 21308 39506 21364 39508
rect 21308 39454 21310 39506
rect 21310 39454 21362 39506
rect 21362 39454 21364 39506
rect 21308 39452 21364 39454
rect 21644 39506 21700 39508
rect 21644 39454 21646 39506
rect 21646 39454 21698 39506
rect 21698 39454 21700 39506
rect 21644 39452 21700 39454
rect 20748 38892 20804 38948
rect 20300 38668 20356 38724
rect 19516 37996 19572 38052
rect 19628 37884 19684 37940
rect 18956 36428 19012 36484
rect 19180 37436 19236 37492
rect 19516 36370 19572 36372
rect 19516 36318 19518 36370
rect 19518 36318 19570 36370
rect 19570 36318 19572 36370
rect 19516 36316 19572 36318
rect 19740 37772 19796 37828
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19740 37436 19796 37492
rect 20412 37938 20468 37940
rect 20412 37886 20414 37938
rect 20414 37886 20466 37938
rect 20466 37886 20468 37938
rect 20412 37884 20468 37886
rect 20636 37772 20692 37828
rect 21308 37996 21364 38052
rect 20412 36370 20468 36372
rect 20412 36318 20414 36370
rect 20414 36318 20466 36370
rect 20466 36318 20468 36370
rect 20412 36316 20468 36318
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 17612 35756 17668 35812
rect 18172 35810 18228 35812
rect 18172 35758 18174 35810
rect 18174 35758 18226 35810
rect 18226 35758 18228 35810
rect 18172 35756 18228 35758
rect 17164 35532 17220 35588
rect 18956 35586 19012 35588
rect 18956 35534 18958 35586
rect 18958 35534 19010 35586
rect 19010 35534 19012 35586
rect 18956 35532 19012 35534
rect 18396 35308 18452 35364
rect 17164 34914 17220 34916
rect 17164 34862 17166 34914
rect 17166 34862 17218 34914
rect 17218 34862 17220 34914
rect 17164 34860 17220 34862
rect 17724 34914 17780 34916
rect 17724 34862 17726 34914
rect 17726 34862 17778 34914
rect 17778 34862 17780 34914
rect 17724 34860 17780 34862
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 17836 34300 17892 34356
rect 16268 34018 16324 34020
rect 16268 33966 16270 34018
rect 16270 33966 16322 34018
rect 16322 33966 16324 34018
rect 16268 33964 16324 33966
rect 16156 33068 16212 33124
rect 15036 32396 15092 32452
rect 9100 29426 9156 29428
rect 9100 29374 9102 29426
rect 9102 29374 9154 29426
rect 9154 29374 9156 29426
rect 9100 29372 9156 29374
rect 9660 29426 9716 29428
rect 9660 29374 9662 29426
rect 9662 29374 9714 29426
rect 9714 29374 9716 29426
rect 9660 29372 9716 29374
rect 9884 28588 9940 28644
rect 9884 27858 9940 27860
rect 9884 27806 9886 27858
rect 9886 27806 9938 27858
rect 9938 27806 9940 27858
rect 9884 27804 9940 27806
rect 9100 26012 9156 26068
rect 11564 29372 11620 29428
rect 10220 28252 10276 28308
rect 10556 27970 10612 27972
rect 10556 27918 10558 27970
rect 10558 27918 10610 27970
rect 10610 27918 10612 27970
rect 10556 27916 10612 27918
rect 10892 27858 10948 27860
rect 10892 27806 10894 27858
rect 10894 27806 10946 27858
rect 10946 27806 10948 27858
rect 10892 27804 10948 27806
rect 12348 30156 12404 30212
rect 13692 30210 13748 30212
rect 13692 30158 13694 30210
rect 13694 30158 13746 30210
rect 13746 30158 13748 30210
rect 13692 30156 13748 30158
rect 14028 30210 14084 30212
rect 14028 30158 14030 30210
rect 14030 30158 14082 30210
rect 14082 30158 14084 30210
rect 14028 30156 14084 30158
rect 12348 29932 12404 29988
rect 15036 30156 15092 30212
rect 16716 32508 16772 32564
rect 16380 30828 16436 30884
rect 16828 32450 16884 32452
rect 16828 32398 16830 32450
rect 16830 32398 16882 32450
rect 16882 32398 16884 32450
rect 16828 32396 16884 32398
rect 17052 32956 17108 33012
rect 16940 31106 16996 31108
rect 16940 31054 16942 31106
rect 16942 31054 16994 31106
rect 16994 31054 16996 31106
rect 16940 31052 16996 31054
rect 16716 30604 16772 30660
rect 14028 29932 14084 29988
rect 13244 29708 13300 29764
rect 11452 28476 11508 28532
rect 11452 27858 11508 27860
rect 11452 27806 11454 27858
rect 11454 27806 11506 27858
rect 11506 27806 11508 27858
rect 11452 27804 11508 27806
rect 11116 27244 11172 27300
rect 10108 27132 10164 27188
rect 12908 28754 12964 28756
rect 12908 28702 12910 28754
rect 12910 28702 12962 28754
rect 12962 28702 12964 28754
rect 12908 28700 12964 28702
rect 12684 27970 12740 27972
rect 12684 27918 12686 27970
rect 12686 27918 12738 27970
rect 12738 27918 12740 27970
rect 12684 27916 12740 27918
rect 11900 27634 11956 27636
rect 11900 27582 11902 27634
rect 11902 27582 11954 27634
rect 11954 27582 11956 27634
rect 11900 27580 11956 27582
rect 11564 26796 11620 26852
rect 9772 26290 9828 26292
rect 9772 26238 9774 26290
rect 9774 26238 9826 26290
rect 9826 26238 9828 26290
rect 9772 26236 9828 26238
rect 10892 26290 10948 26292
rect 10892 26238 10894 26290
rect 10894 26238 10946 26290
rect 10946 26238 10948 26290
rect 10892 26236 10948 26238
rect 9324 25676 9380 25732
rect 8316 25340 8372 25396
rect 8316 24556 8372 24612
rect 8204 21420 8260 21476
rect 7980 20802 8036 20804
rect 7980 20750 7982 20802
rect 7982 20750 8034 20802
rect 8034 20750 8036 20802
rect 7980 20748 8036 20750
rect 8988 25506 9044 25508
rect 8988 25454 8990 25506
rect 8990 25454 9042 25506
rect 9042 25454 9044 25506
rect 8988 25452 9044 25454
rect 9436 25340 9492 25396
rect 10220 25452 10276 25508
rect 9548 25228 9604 25284
rect 9772 25228 9828 25284
rect 8652 21868 8708 21924
rect 8428 20802 8484 20804
rect 8428 20750 8430 20802
rect 8430 20750 8482 20802
rect 8482 20750 8484 20802
rect 8428 20748 8484 20750
rect 7980 19906 8036 19908
rect 7980 19854 7982 19906
rect 7982 19854 8034 19906
rect 8034 19854 8036 19906
rect 7980 19852 8036 19854
rect 9324 23548 9380 23604
rect 8988 21532 9044 21588
rect 9212 22146 9268 22148
rect 9212 22094 9214 22146
rect 9214 22094 9266 22146
rect 9266 22094 9268 22146
rect 9212 22092 9268 22094
rect 9212 21756 9268 21812
rect 9436 21756 9492 21812
rect 8988 19906 9044 19908
rect 8988 19854 8990 19906
rect 8990 19854 9042 19906
rect 9042 19854 9044 19906
rect 8988 19852 9044 19854
rect 8316 19346 8372 19348
rect 8316 19294 8318 19346
rect 8318 19294 8370 19346
rect 8370 19294 8372 19346
rect 8316 19292 8372 19294
rect 6188 17724 6244 17780
rect 8652 17778 8708 17780
rect 8652 17726 8654 17778
rect 8654 17726 8706 17778
rect 8706 17726 8708 17778
rect 8652 17724 8708 17726
rect 9212 20300 9268 20356
rect 10668 24556 10724 24612
rect 11676 26460 11732 26516
rect 11452 25452 11508 25508
rect 10892 23938 10948 23940
rect 10892 23886 10894 23938
rect 10894 23886 10946 23938
rect 10946 23886 10948 23938
rect 10892 23884 10948 23886
rect 11900 23938 11956 23940
rect 11900 23886 11902 23938
rect 11902 23886 11954 23938
rect 11954 23886 11956 23938
rect 11900 23884 11956 23886
rect 10108 23324 10164 23380
rect 10220 23660 10276 23716
rect 9772 21980 9828 22036
rect 9660 21420 9716 21476
rect 9884 21084 9940 21140
rect 9660 20300 9716 20356
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 12684 25564 12740 25620
rect 12684 24780 12740 24836
rect 13916 28700 13972 28756
rect 13692 27916 13748 27972
rect 13804 27020 13860 27076
rect 15596 29260 15652 29316
rect 15708 28754 15764 28756
rect 15708 28702 15710 28754
rect 15710 28702 15762 28754
rect 15762 28702 15764 28754
rect 15708 28700 15764 28702
rect 16380 28754 16436 28756
rect 16380 28702 16382 28754
rect 16382 28702 16434 28754
rect 16434 28702 16436 28754
rect 16380 28700 16436 28702
rect 14028 28028 14084 28084
rect 15036 28364 15092 28420
rect 14812 27074 14868 27076
rect 14812 27022 14814 27074
rect 14814 27022 14866 27074
rect 14866 27022 14868 27074
rect 14812 27020 14868 27022
rect 14700 26908 14756 26964
rect 13580 26460 13636 26516
rect 16492 28418 16548 28420
rect 16492 28366 16494 28418
rect 16494 28366 16546 28418
rect 16546 28366 16548 28418
rect 16492 28364 16548 28366
rect 15372 26908 15428 26964
rect 15932 27020 15988 27076
rect 16380 27746 16436 27748
rect 16380 27694 16382 27746
rect 16382 27694 16434 27746
rect 16434 27694 16436 27746
rect 16380 27692 16436 27694
rect 16380 26908 16436 26964
rect 16828 30268 16884 30324
rect 17276 32508 17332 32564
rect 16828 29596 16884 29652
rect 15596 26796 15652 26852
rect 16380 26460 16436 26516
rect 15484 26012 15540 26068
rect 12684 23884 12740 23940
rect 12572 23660 12628 23716
rect 12124 23548 12180 23604
rect 10892 23324 10948 23380
rect 10892 22876 10948 22932
rect 10780 22092 10836 22148
rect 10556 21756 10612 21812
rect 11004 21644 11060 21700
rect 11900 21868 11956 21924
rect 12572 21980 12628 22036
rect 12460 21756 12516 21812
rect 11788 20636 11844 20692
rect 11340 18396 11396 18452
rect 12684 20860 12740 20916
rect 12684 20300 12740 20356
rect 12908 23938 12964 23940
rect 12908 23886 12910 23938
rect 12910 23886 12962 23938
rect 12962 23886 12964 23938
rect 12908 23884 12964 23886
rect 12908 23548 12964 23604
rect 13356 24722 13412 24724
rect 13356 24670 13358 24722
rect 13358 24670 13410 24722
rect 13410 24670 13412 24722
rect 13356 24668 13412 24670
rect 13356 23548 13412 23604
rect 13244 22930 13300 22932
rect 13244 22878 13246 22930
rect 13246 22878 13298 22930
rect 13298 22878 13300 22930
rect 13244 22876 13300 22878
rect 13020 21084 13076 21140
rect 13580 22370 13636 22372
rect 13580 22318 13582 22370
rect 13582 22318 13634 22370
rect 13634 22318 13636 22370
rect 13580 22316 13636 22318
rect 13468 20914 13524 20916
rect 13468 20862 13470 20914
rect 13470 20862 13522 20914
rect 13522 20862 13524 20914
rect 13468 20860 13524 20862
rect 13916 21868 13972 21924
rect 13804 21756 13860 21812
rect 13692 20636 13748 20692
rect 15260 20914 15316 20916
rect 15260 20862 15262 20914
rect 15262 20862 15314 20914
rect 15314 20862 15316 20914
rect 15260 20860 15316 20862
rect 16380 25788 16436 25844
rect 15820 25228 15876 25284
rect 15708 24444 15764 24500
rect 16380 23996 16436 24052
rect 15820 22316 15876 22372
rect 15596 21196 15652 21252
rect 15708 20748 15764 20804
rect 15484 19906 15540 19908
rect 15484 19854 15486 19906
rect 15486 19854 15538 19906
rect 15538 19854 15540 19906
rect 15484 19852 15540 19854
rect 14924 19628 14980 19684
rect 16268 21644 16324 21700
rect 16380 22092 16436 22148
rect 16156 21196 16212 21252
rect 9884 15932 9940 15988
rect 10892 15986 10948 15988
rect 10892 15934 10894 15986
rect 10894 15934 10946 15986
rect 10946 15934 10948 15986
rect 10892 15932 10948 15934
rect 16380 20802 16436 20804
rect 16380 20750 16382 20802
rect 16382 20750 16434 20802
rect 16434 20750 16436 20802
rect 16380 20748 16436 20750
rect 16380 20524 16436 20580
rect 16492 18284 16548 18340
rect 17612 32396 17668 32452
rect 22428 39452 22484 39508
rect 24220 48524 24276 48580
rect 24332 47516 24388 47572
rect 25228 48524 25284 48580
rect 25452 49644 25508 49700
rect 24668 47346 24724 47348
rect 24668 47294 24670 47346
rect 24670 47294 24722 47346
rect 24722 47294 24724 47346
rect 24668 47292 24724 47294
rect 24444 46450 24500 46452
rect 24444 46398 24446 46450
rect 24446 46398 24498 46450
rect 24498 46398 24500 46450
rect 24444 46396 24500 46398
rect 24332 45612 24388 45668
rect 24108 44828 24164 44884
rect 24220 43820 24276 43876
rect 23772 42588 23828 42644
rect 25676 49756 25732 49812
rect 26124 49698 26180 49700
rect 26124 49646 26126 49698
rect 26126 49646 26178 49698
rect 26178 49646 26180 49698
rect 26124 49644 26180 49646
rect 25340 47964 25396 48020
rect 25116 47516 25172 47572
rect 25340 47404 25396 47460
rect 26572 48860 26628 48916
rect 25676 48130 25732 48132
rect 25676 48078 25678 48130
rect 25678 48078 25730 48130
rect 25730 48078 25732 48130
rect 25676 48076 25732 48078
rect 25900 47964 25956 48020
rect 25116 46620 25172 46676
rect 25116 45890 25172 45892
rect 25116 45838 25118 45890
rect 25118 45838 25170 45890
rect 25170 45838 25172 45890
rect 25116 45836 25172 45838
rect 24892 44940 24948 44996
rect 25564 46956 25620 47012
rect 27916 51436 27972 51492
rect 27244 49756 27300 49812
rect 27356 48802 27412 48804
rect 27356 48750 27358 48802
rect 27358 48750 27410 48802
rect 27410 48750 27412 48802
rect 27356 48748 27412 48750
rect 27132 47292 27188 47348
rect 26460 46620 26516 46676
rect 25676 45164 25732 45220
rect 24780 43820 24836 43876
rect 25788 44044 25844 44100
rect 25004 42252 25060 42308
rect 23996 41970 24052 41972
rect 23996 41918 23998 41970
rect 23998 41918 24050 41970
rect 24050 41918 24052 41970
rect 23996 41916 24052 41918
rect 23660 41804 23716 41860
rect 23548 40908 23604 40964
rect 24108 40402 24164 40404
rect 24108 40350 24110 40402
rect 24110 40350 24162 40402
rect 24162 40350 24164 40402
rect 24108 40348 24164 40350
rect 22876 39506 22932 39508
rect 22876 39454 22878 39506
rect 22878 39454 22930 39506
rect 22930 39454 22932 39506
rect 22876 39452 22932 39454
rect 22204 39004 22260 39060
rect 21644 37772 21700 37828
rect 21644 37266 21700 37268
rect 21644 37214 21646 37266
rect 21646 37214 21698 37266
rect 21698 37214 21700 37266
rect 21644 37212 21700 37214
rect 21532 35196 21588 35252
rect 20972 34636 21028 34692
rect 20860 34188 20916 34244
rect 20748 34076 20804 34132
rect 20412 33404 20468 33460
rect 20076 33292 20132 33348
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 18396 32562 18452 32564
rect 18396 32510 18398 32562
rect 18398 32510 18450 32562
rect 18450 32510 18452 32562
rect 18396 32508 18452 32510
rect 17724 32172 17780 32228
rect 19516 32450 19572 32452
rect 19516 32398 19518 32450
rect 19518 32398 19570 32450
rect 19570 32398 19572 32450
rect 19516 32396 19572 32398
rect 17724 31778 17780 31780
rect 17724 31726 17726 31778
rect 17726 31726 17778 31778
rect 17778 31726 17780 31778
rect 17724 31724 17780 31726
rect 18844 31500 18900 31556
rect 17836 30828 17892 30884
rect 18508 30604 18564 30660
rect 18620 30210 18676 30212
rect 18620 30158 18622 30210
rect 18622 30158 18674 30210
rect 18674 30158 18676 30210
rect 18620 30156 18676 30158
rect 17500 29650 17556 29652
rect 17500 29598 17502 29650
rect 17502 29598 17554 29650
rect 17554 29598 17556 29650
rect 17500 29596 17556 29598
rect 17948 29650 18004 29652
rect 17948 29598 17950 29650
rect 17950 29598 18002 29650
rect 18002 29598 18004 29650
rect 17948 29596 18004 29598
rect 20076 31948 20132 32004
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20860 32620 20916 32676
rect 22092 36316 22148 36372
rect 21756 33852 21812 33908
rect 21980 34076 22036 34132
rect 21644 33740 21700 33796
rect 21420 33458 21476 33460
rect 21420 33406 21422 33458
rect 21422 33406 21474 33458
rect 21474 33406 21476 33458
rect 21420 33404 21476 33406
rect 21084 32396 21140 32452
rect 21196 32732 21252 32788
rect 21644 32396 21700 32452
rect 20972 31724 21028 31780
rect 20860 31666 20916 31668
rect 20860 31614 20862 31666
rect 20862 31614 20914 31666
rect 20914 31614 20916 31666
rect 20860 31612 20916 31614
rect 20300 30940 20356 30996
rect 20188 30492 20244 30548
rect 20300 30268 20356 30324
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19068 29596 19124 29652
rect 17724 28924 17780 28980
rect 17948 28082 18004 28084
rect 17948 28030 17950 28082
rect 17950 28030 18002 28082
rect 18002 28030 18004 28082
rect 17948 28028 18004 28030
rect 20748 30268 20804 30324
rect 20300 29650 20356 29652
rect 20300 29598 20302 29650
rect 20302 29598 20354 29650
rect 20354 29598 20356 29650
rect 20300 29596 20356 29598
rect 22764 38668 22820 38724
rect 22652 38162 22708 38164
rect 22652 38110 22654 38162
rect 22654 38110 22706 38162
rect 22706 38110 22708 38162
rect 22652 38108 22708 38110
rect 22652 36594 22708 36596
rect 22652 36542 22654 36594
rect 22654 36542 22706 36594
rect 22706 36542 22708 36594
rect 22652 36540 22708 36542
rect 24332 41858 24388 41860
rect 24332 41806 24334 41858
rect 24334 41806 24386 41858
rect 24386 41806 24388 41858
rect 24332 41804 24388 41806
rect 24780 41804 24836 41860
rect 24444 41298 24500 41300
rect 24444 41246 24446 41298
rect 24446 41246 24498 41298
rect 24498 41246 24500 41298
rect 24444 41244 24500 41246
rect 25452 41858 25508 41860
rect 25452 41806 25454 41858
rect 25454 41806 25506 41858
rect 25506 41806 25508 41858
rect 25452 41804 25508 41806
rect 24668 40402 24724 40404
rect 24668 40350 24670 40402
rect 24670 40350 24722 40402
rect 24722 40350 24724 40402
rect 24668 40348 24724 40350
rect 24332 39618 24388 39620
rect 24332 39566 24334 39618
rect 24334 39566 24386 39618
rect 24386 39566 24388 39618
rect 24332 39564 24388 39566
rect 25340 40236 25396 40292
rect 24780 40124 24836 40180
rect 23996 38050 24052 38052
rect 23996 37998 23998 38050
rect 23998 37998 24050 38050
rect 24050 37998 24052 38050
rect 23996 37996 24052 37998
rect 24668 37996 24724 38052
rect 24780 39900 24836 39956
rect 24556 37884 24612 37940
rect 24220 37324 24276 37380
rect 24556 36482 24612 36484
rect 24556 36430 24558 36482
rect 24558 36430 24610 36482
rect 24610 36430 24612 36482
rect 24556 36428 24612 36430
rect 23212 35868 23268 35924
rect 22876 35698 22932 35700
rect 22876 35646 22878 35698
rect 22878 35646 22930 35698
rect 22930 35646 22932 35698
rect 22876 35644 22932 35646
rect 24220 35644 24276 35700
rect 24444 35644 24500 35700
rect 24220 34972 24276 35028
rect 22540 33346 22596 33348
rect 22540 33294 22542 33346
rect 22542 33294 22594 33346
rect 22594 33294 22596 33346
rect 22540 33292 22596 33294
rect 22764 33516 22820 33572
rect 23548 33516 23604 33572
rect 25228 37378 25284 37380
rect 25228 37326 25230 37378
rect 25230 37326 25282 37378
rect 25282 37326 25284 37378
rect 25228 37324 25284 37326
rect 25900 42252 25956 42308
rect 25676 41804 25732 41860
rect 25788 41692 25844 41748
rect 25564 40514 25620 40516
rect 25564 40462 25566 40514
rect 25566 40462 25618 40514
rect 25618 40462 25620 40514
rect 25564 40460 25620 40462
rect 26684 45106 26740 45108
rect 26684 45054 26686 45106
rect 26686 45054 26738 45106
rect 26738 45054 26740 45106
rect 26684 45052 26740 45054
rect 26572 42028 26628 42084
rect 26460 41692 26516 41748
rect 27132 41970 27188 41972
rect 27132 41918 27134 41970
rect 27134 41918 27186 41970
rect 27186 41918 27188 41970
rect 27132 41916 27188 41918
rect 26684 41244 26740 41300
rect 25788 40572 25844 40628
rect 25340 36876 25396 36932
rect 25340 35644 25396 35700
rect 27356 45164 27412 45220
rect 27916 49698 27972 49700
rect 27916 49646 27918 49698
rect 27918 49646 27970 49698
rect 27970 49646 27972 49698
rect 27916 49644 27972 49646
rect 28140 49644 28196 49700
rect 28028 48860 28084 48916
rect 27916 47180 27972 47236
rect 28252 48802 28308 48804
rect 28252 48750 28254 48802
rect 28254 48750 28306 48802
rect 28306 48750 28308 48802
rect 28252 48748 28308 48750
rect 28140 46844 28196 46900
rect 28140 46674 28196 46676
rect 28140 46622 28142 46674
rect 28142 46622 28194 46674
rect 28194 46622 28196 46674
rect 28140 46620 28196 46622
rect 28476 48748 28532 48804
rect 30380 53842 30436 53844
rect 30380 53790 30382 53842
rect 30382 53790 30434 53842
rect 30434 53790 30436 53842
rect 30380 53788 30436 53790
rect 29036 51490 29092 51492
rect 29036 51438 29038 51490
rect 29038 51438 29090 51490
rect 29090 51438 29092 51490
rect 29036 51436 29092 51438
rect 28700 48860 28756 48916
rect 28812 48748 28868 48804
rect 28364 46284 28420 46340
rect 29036 46620 29092 46676
rect 29036 46114 29092 46116
rect 29036 46062 29038 46114
rect 29038 46062 29090 46114
rect 29090 46062 29092 46114
rect 29036 46060 29092 46062
rect 28364 44098 28420 44100
rect 28364 44046 28366 44098
rect 28366 44046 28418 44098
rect 28418 44046 28420 44098
rect 28364 44044 28420 44046
rect 27916 42476 27972 42532
rect 28140 41916 28196 41972
rect 27132 40908 27188 40964
rect 26460 36428 26516 36484
rect 26012 35698 26068 35700
rect 26012 35646 26014 35698
rect 26014 35646 26066 35698
rect 26066 35646 26068 35698
rect 26012 35644 26068 35646
rect 26348 35026 26404 35028
rect 26348 34974 26350 35026
rect 26350 34974 26402 35026
rect 26402 34974 26404 35026
rect 26348 34972 26404 34974
rect 28028 41692 28084 41748
rect 27916 41580 27972 41636
rect 28252 42812 28308 42868
rect 29148 45052 29204 45108
rect 28700 43650 28756 43652
rect 28700 43598 28702 43650
rect 28702 43598 28754 43650
rect 28754 43598 28756 43650
rect 28700 43596 28756 43598
rect 28476 42476 28532 42532
rect 28476 40684 28532 40740
rect 27916 39730 27972 39732
rect 27916 39678 27918 39730
rect 27918 39678 27970 39730
rect 27970 39678 27972 39730
rect 27916 39676 27972 39678
rect 28588 40348 28644 40404
rect 28700 40460 28756 40516
rect 28924 40402 28980 40404
rect 28924 40350 28926 40402
rect 28926 40350 28978 40402
rect 28978 40350 28980 40402
rect 28924 40348 28980 40350
rect 28812 38946 28868 38948
rect 28812 38894 28814 38946
rect 28814 38894 28866 38946
rect 28866 38894 28868 38946
rect 28812 38892 28868 38894
rect 28028 38668 28084 38724
rect 27692 38332 27748 38388
rect 27804 37212 27860 37268
rect 28364 38220 28420 38276
rect 25788 33292 25844 33348
rect 24556 32956 24612 33012
rect 23548 32508 23604 32564
rect 22204 31836 22260 31892
rect 22316 32396 22372 32452
rect 21308 30940 21364 30996
rect 21308 30268 21364 30324
rect 21644 30210 21700 30212
rect 21644 30158 21646 30210
rect 21646 30158 21698 30210
rect 21698 30158 21700 30210
rect 21644 30156 21700 30158
rect 23324 32450 23380 32452
rect 23324 32398 23326 32450
rect 23326 32398 23378 32450
rect 23378 32398 23380 32450
rect 23324 32396 23380 32398
rect 22988 31948 23044 32004
rect 23772 32396 23828 32452
rect 23548 30882 23604 30884
rect 23548 30830 23550 30882
rect 23550 30830 23602 30882
rect 23602 30830 23604 30882
rect 23548 30828 23604 30830
rect 23212 30380 23268 30436
rect 22316 30210 22372 30212
rect 22316 30158 22318 30210
rect 22318 30158 22370 30210
rect 22370 30158 22372 30210
rect 22316 30156 22372 30158
rect 21644 29426 21700 29428
rect 21644 29374 21646 29426
rect 21646 29374 21698 29426
rect 21698 29374 21700 29426
rect 21644 29372 21700 29374
rect 19852 29314 19908 29316
rect 19852 29262 19854 29314
rect 19854 29262 19906 29314
rect 19906 29262 19908 29314
rect 19852 29260 19908 29262
rect 22540 29148 22596 29204
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17612 27746 17668 27748
rect 17612 27694 17614 27746
rect 17614 27694 17666 27746
rect 17666 27694 17668 27746
rect 17612 27692 17668 27694
rect 18172 27692 18228 27748
rect 19740 27746 19796 27748
rect 19740 27694 19742 27746
rect 19742 27694 19794 27746
rect 19794 27694 19796 27746
rect 19740 27692 19796 27694
rect 17276 26066 17332 26068
rect 17276 26014 17278 26066
rect 17278 26014 17330 26066
rect 17330 26014 17332 26066
rect 17276 26012 17332 26014
rect 17276 25788 17332 25844
rect 16828 24444 16884 24500
rect 17388 25228 17444 25284
rect 17612 24722 17668 24724
rect 17612 24670 17614 24722
rect 17614 24670 17666 24722
rect 17666 24670 17668 24722
rect 17612 24668 17668 24670
rect 17164 22370 17220 22372
rect 17164 22318 17166 22370
rect 17166 22318 17218 22370
rect 17218 22318 17220 22370
rect 17164 22316 17220 22318
rect 17052 22146 17108 22148
rect 17052 22094 17054 22146
rect 17054 22094 17106 22146
rect 17106 22094 17108 22146
rect 17052 22092 17108 22094
rect 17276 21756 17332 21812
rect 16716 20860 16772 20916
rect 16828 20524 16884 20580
rect 16828 19964 16884 20020
rect 16828 19346 16884 19348
rect 16828 19294 16830 19346
rect 16830 19294 16882 19346
rect 16882 19294 16884 19346
rect 16828 19292 16884 19294
rect 17500 22316 17556 22372
rect 17500 20130 17556 20132
rect 17500 20078 17502 20130
rect 17502 20078 17554 20130
rect 17554 20078 17556 20130
rect 17500 20076 17556 20078
rect 17612 21980 17668 22036
rect 17388 19852 17444 19908
rect 17500 18956 17556 19012
rect 19740 27020 19796 27076
rect 20300 27244 20356 27300
rect 20076 26962 20132 26964
rect 20076 26910 20078 26962
rect 20078 26910 20130 26962
rect 20130 26910 20132 26962
rect 20076 26908 20132 26910
rect 19964 26796 20020 26852
rect 20748 27692 20804 27748
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18284 26460 18340 26516
rect 18060 25676 18116 25732
rect 17948 25004 18004 25060
rect 17948 24722 18004 24724
rect 17948 24670 17950 24722
rect 17950 24670 18002 24722
rect 18002 24670 18004 24722
rect 17948 24668 18004 24670
rect 17836 20300 17892 20356
rect 18060 20188 18116 20244
rect 18172 20524 18228 20580
rect 17836 20018 17892 20020
rect 17836 19966 17838 20018
rect 17838 19966 17890 20018
rect 17890 19966 17892 20018
rect 17836 19964 17892 19966
rect 17724 19292 17780 19348
rect 19516 26236 19572 26292
rect 19404 25730 19460 25732
rect 19404 25678 19406 25730
rect 19406 25678 19458 25730
rect 19458 25678 19460 25730
rect 19404 25676 19460 25678
rect 18844 24444 18900 24500
rect 18732 20578 18788 20580
rect 18732 20526 18734 20578
rect 18734 20526 18786 20578
rect 18786 20526 18788 20578
rect 18732 20524 18788 20526
rect 18620 20300 18676 20356
rect 18508 20188 18564 20244
rect 18508 19516 18564 19572
rect 18844 20018 18900 20020
rect 18844 19966 18846 20018
rect 18846 19966 18898 20018
rect 18898 19966 18900 20018
rect 18844 19964 18900 19966
rect 19292 25340 19348 25396
rect 19180 25116 19236 25172
rect 19180 24780 19236 24836
rect 19068 24050 19124 24052
rect 19068 23998 19070 24050
rect 19070 23998 19122 24050
rect 19122 23998 19124 24050
rect 19068 23996 19124 23998
rect 19068 21756 19124 21812
rect 19068 20076 19124 20132
rect 19068 18508 19124 18564
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 19628 25116 19684 25172
rect 20188 25452 20244 25508
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 25228 20356 25284
rect 19628 24834 19684 24836
rect 19628 24782 19630 24834
rect 19630 24782 19682 24834
rect 19682 24782 19684 24834
rect 19628 24780 19684 24782
rect 19852 24498 19908 24500
rect 19852 24446 19854 24498
rect 19854 24446 19906 24498
rect 19906 24446 19908 24498
rect 19852 24444 19908 24446
rect 20300 23884 20356 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 20860 19348 20916
rect 19292 19964 19348 20020
rect 19516 23100 19572 23156
rect 20300 23154 20356 23156
rect 20300 23102 20302 23154
rect 20302 23102 20354 23154
rect 20354 23102 20356 23154
rect 20300 23100 20356 23102
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19740 20914 19796 20916
rect 19740 20862 19742 20914
rect 19742 20862 19794 20914
rect 19794 20862 19796 20914
rect 19740 20860 19796 20862
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19516 19516 19572 19572
rect 19516 19180 19572 19236
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20412 20914 20468 20916
rect 20412 20862 20414 20914
rect 20414 20862 20466 20914
rect 20466 20862 20468 20914
rect 20412 20860 20468 20862
rect 20300 19010 20356 19012
rect 20300 18958 20302 19010
rect 20302 18958 20354 19010
rect 20354 18958 20356 19010
rect 20300 18956 20356 18958
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21308 27298 21364 27300
rect 21308 27246 21310 27298
rect 21310 27246 21362 27298
rect 21362 27246 21364 27298
rect 21308 27244 21364 27246
rect 22316 27804 22372 27860
rect 21532 27074 21588 27076
rect 21532 27022 21534 27074
rect 21534 27022 21586 27074
rect 21586 27022 21588 27074
rect 21532 27020 21588 27022
rect 22428 27074 22484 27076
rect 22428 27022 22430 27074
rect 22430 27022 22482 27074
rect 22482 27022 22484 27074
rect 22428 27020 22484 27022
rect 20860 26460 20916 26516
rect 20636 25506 20692 25508
rect 20636 25454 20638 25506
rect 20638 25454 20690 25506
rect 20690 25454 20692 25506
rect 20636 25452 20692 25454
rect 20748 25228 20804 25284
rect 20748 24892 20804 24948
rect 21532 26684 21588 26740
rect 21756 26348 21812 26404
rect 21644 26290 21700 26292
rect 21644 26238 21646 26290
rect 21646 26238 21698 26290
rect 21698 26238 21700 26290
rect 21644 26236 21700 26238
rect 21420 25394 21476 25396
rect 21420 25342 21422 25394
rect 21422 25342 21474 25394
rect 21474 25342 21476 25394
rect 21420 25340 21476 25342
rect 21308 24892 21364 24948
rect 21196 23938 21252 23940
rect 21196 23886 21198 23938
rect 21198 23886 21250 23938
rect 21250 23886 21252 23938
rect 21196 23884 21252 23886
rect 20748 22316 20804 22372
rect 20636 20076 20692 20132
rect 20636 19346 20692 19348
rect 20636 19294 20638 19346
rect 20638 19294 20690 19346
rect 20690 19294 20692 19346
rect 20636 19292 20692 19294
rect 20412 16716 20468 16772
rect 19740 16604 19796 16660
rect 20300 16604 20356 16660
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21420 19346 21476 19348
rect 21420 19294 21422 19346
rect 21422 19294 21474 19346
rect 21474 19294 21476 19346
rect 21420 19292 21476 19294
rect 23996 31724 24052 31780
rect 24220 31612 24276 31668
rect 23996 30268 24052 30324
rect 24332 30380 24388 30436
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 24668 31778 24724 31780
rect 24668 31726 24670 31778
rect 24670 31726 24722 31778
rect 24722 31726 24724 31778
rect 24668 31724 24724 31726
rect 25900 32562 25956 32564
rect 25900 32510 25902 32562
rect 25902 32510 25954 32562
rect 25954 32510 25956 32562
rect 25900 32508 25956 32510
rect 25004 31554 25060 31556
rect 25004 31502 25006 31554
rect 25006 31502 25058 31554
rect 25058 31502 25060 31554
rect 25004 31500 25060 31502
rect 25452 31218 25508 31220
rect 25452 31166 25454 31218
rect 25454 31166 25506 31218
rect 25506 31166 25508 31218
rect 25452 31164 25508 31166
rect 27132 32508 27188 32564
rect 27692 33292 27748 33348
rect 26684 32396 26740 32452
rect 26572 31612 26628 31668
rect 26012 30882 26068 30884
rect 26012 30830 26014 30882
rect 26014 30830 26066 30882
rect 26066 30830 26068 30882
rect 26012 30828 26068 30830
rect 25900 30604 25956 30660
rect 24556 29260 24612 29316
rect 25116 29932 25172 29988
rect 23548 29036 23604 29092
rect 24444 29036 24500 29092
rect 22092 22540 22148 22596
rect 21756 20860 21812 20916
rect 22092 19180 22148 19236
rect 21532 18396 21588 18452
rect 21868 18338 21924 18340
rect 21868 18286 21870 18338
rect 21870 18286 21922 18338
rect 21922 18286 21924 18338
rect 21868 18284 21924 18286
rect 24220 28140 24276 28196
rect 23772 27916 23828 27972
rect 23212 27804 23268 27860
rect 22764 22540 22820 22596
rect 23100 27580 23156 27636
rect 22764 22370 22820 22372
rect 22764 22318 22766 22370
rect 22766 22318 22818 22370
rect 22818 22318 22820 22370
rect 22764 22316 22820 22318
rect 23660 27858 23716 27860
rect 23660 27806 23662 27858
rect 23662 27806 23714 27858
rect 23714 27806 23716 27858
rect 23660 27804 23716 27806
rect 23660 27074 23716 27076
rect 23660 27022 23662 27074
rect 23662 27022 23714 27074
rect 23714 27022 23716 27074
rect 23660 27020 23716 27022
rect 24108 27804 24164 27860
rect 23884 26908 23940 26964
rect 23996 26402 24052 26404
rect 23996 26350 23998 26402
rect 23998 26350 24050 26402
rect 24050 26350 24052 26402
rect 23996 26348 24052 26350
rect 24220 27692 24276 27748
rect 24668 27746 24724 27748
rect 24668 27694 24670 27746
rect 24670 27694 24722 27746
rect 24722 27694 24724 27746
rect 24668 27692 24724 27694
rect 24668 27132 24724 27188
rect 25340 29426 25396 29428
rect 25340 29374 25342 29426
rect 25342 29374 25394 29426
rect 25394 29374 25396 29426
rect 25340 29372 25396 29374
rect 25788 29036 25844 29092
rect 25788 28866 25844 28868
rect 25788 28814 25790 28866
rect 25790 28814 25842 28866
rect 25842 28814 25844 28866
rect 25788 28812 25844 28814
rect 26012 28028 26068 28084
rect 25228 27692 25284 27748
rect 24332 24892 24388 24948
rect 23324 24722 23380 24724
rect 23324 24670 23326 24722
rect 23326 24670 23378 24722
rect 23378 24670 23380 24722
rect 23324 24668 23380 24670
rect 23324 23884 23380 23940
rect 24332 23660 24388 23716
rect 22540 19292 22596 19348
rect 23996 22092 24052 22148
rect 23212 20188 23268 20244
rect 23212 19292 23268 19348
rect 23884 21586 23940 21588
rect 23884 21534 23886 21586
rect 23886 21534 23938 21586
rect 23938 21534 23940 21586
rect 23884 21532 23940 21534
rect 23548 20018 23604 20020
rect 23548 19966 23550 20018
rect 23550 19966 23602 20018
rect 23602 19966 23604 20018
rect 23548 19964 23604 19966
rect 23772 19068 23828 19124
rect 23884 19292 23940 19348
rect 23996 18508 24052 18564
rect 23660 18396 23716 18452
rect 24220 20242 24276 20244
rect 24220 20190 24222 20242
rect 24222 20190 24274 20242
rect 24274 20190 24276 20242
rect 24220 20188 24276 20190
rect 24108 17724 24164 17780
rect 25116 25228 25172 25284
rect 24556 24668 24612 24724
rect 24668 24780 24724 24836
rect 25228 26236 25284 26292
rect 24892 23714 24948 23716
rect 24892 23662 24894 23714
rect 24894 23662 24946 23714
rect 24946 23662 24948 23714
rect 24892 23660 24948 23662
rect 24780 23154 24836 23156
rect 24780 23102 24782 23154
rect 24782 23102 24834 23154
rect 24834 23102 24836 23154
rect 24780 23100 24836 23102
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 24332 16716 24388 16772
rect 24668 21644 24724 21700
rect 24780 21420 24836 21476
rect 24668 19964 24724 20020
rect 25116 23154 25172 23156
rect 25116 23102 25118 23154
rect 25118 23102 25170 23154
rect 25170 23102 25172 23154
rect 25116 23100 25172 23102
rect 25340 22428 25396 22484
rect 25228 22316 25284 22372
rect 25116 22092 25172 22148
rect 25340 21868 25396 21924
rect 25676 26290 25732 26292
rect 25676 26238 25678 26290
rect 25678 26238 25730 26290
rect 25730 26238 25732 26290
rect 25676 26236 25732 26238
rect 26348 30380 26404 30436
rect 26236 30156 26292 30212
rect 26236 29372 26292 29428
rect 27132 30828 27188 30884
rect 26572 28140 26628 28196
rect 26236 27804 26292 27860
rect 27244 30210 27300 30212
rect 27244 30158 27246 30210
rect 27246 30158 27298 30210
rect 27298 30158 27300 30210
rect 27244 30156 27300 30158
rect 29708 49868 29764 49924
rect 29596 48748 29652 48804
rect 29932 49196 29988 49252
rect 29372 44828 29428 44884
rect 29484 46844 29540 46900
rect 29820 45778 29876 45780
rect 29820 45726 29822 45778
rect 29822 45726 29874 45778
rect 29874 45726 29876 45778
rect 29820 45724 29876 45726
rect 29820 44434 29876 44436
rect 29820 44382 29822 44434
rect 29822 44382 29874 44434
rect 29874 44382 29876 44434
rect 29820 44380 29876 44382
rect 29260 42754 29316 42756
rect 29260 42702 29262 42754
rect 29262 42702 29314 42754
rect 29314 42702 29316 42754
rect 29260 42700 29316 42702
rect 31052 49868 31108 49924
rect 30716 48860 30772 48916
rect 30268 48748 30324 48804
rect 30268 48188 30324 48244
rect 30828 48242 30884 48244
rect 30828 48190 30830 48242
rect 30830 48190 30882 48242
rect 30882 48190 30884 48242
rect 30828 48188 30884 48190
rect 30156 47180 30212 47236
rect 30940 45106 30996 45108
rect 30940 45054 30942 45106
rect 30942 45054 30994 45106
rect 30994 45054 30996 45106
rect 30940 45052 30996 45054
rect 30268 42252 30324 42308
rect 29148 39676 29204 39732
rect 29372 42028 29428 42084
rect 29148 37884 29204 37940
rect 28028 34972 28084 35028
rect 28476 34748 28532 34804
rect 28700 32956 28756 33012
rect 28476 32562 28532 32564
rect 28476 32510 28478 32562
rect 28478 32510 28530 32562
rect 28530 32510 28532 32562
rect 28476 32508 28532 32510
rect 28140 31836 28196 31892
rect 27804 31612 27860 31668
rect 28588 31164 28644 31220
rect 28252 30210 28308 30212
rect 28252 30158 28254 30210
rect 28254 30158 28306 30210
rect 28306 30158 28308 30210
rect 28252 30156 28308 30158
rect 27580 29986 27636 29988
rect 27580 29934 27582 29986
rect 27582 29934 27634 29986
rect 27634 29934 27636 29986
rect 27580 29932 27636 29934
rect 27244 28082 27300 28084
rect 27244 28030 27246 28082
rect 27246 28030 27298 28082
rect 27298 28030 27300 28082
rect 27244 28028 27300 28030
rect 26684 26850 26740 26852
rect 26684 26798 26686 26850
rect 26686 26798 26738 26850
rect 26738 26798 26740 26850
rect 26684 26796 26740 26798
rect 26124 24668 26180 24724
rect 25788 21980 25844 22036
rect 26460 22428 26516 22484
rect 25788 21644 25844 21700
rect 25900 21474 25956 21476
rect 25900 21422 25902 21474
rect 25902 21422 25954 21474
rect 25954 21422 25956 21474
rect 25900 21420 25956 21422
rect 25340 19964 25396 20020
rect 25452 19122 25508 19124
rect 25452 19070 25454 19122
rect 25454 19070 25506 19122
rect 25506 19070 25508 19122
rect 25452 19068 25508 19070
rect 26124 18172 26180 18228
rect 24556 15932 24612 15988
rect 26908 22316 26964 22372
rect 26572 19346 26628 19348
rect 26572 19294 26574 19346
rect 26574 19294 26626 19346
rect 26626 19294 26628 19346
rect 26572 19292 26628 19294
rect 27244 24892 27300 24948
rect 27468 27634 27524 27636
rect 27468 27582 27470 27634
rect 27470 27582 27522 27634
rect 27522 27582 27524 27634
rect 27468 27580 27524 27582
rect 28252 28588 28308 28644
rect 28588 28476 28644 28532
rect 28028 27020 28084 27076
rect 27468 25228 27524 25284
rect 27916 23996 27972 24052
rect 27356 22594 27412 22596
rect 27356 22542 27358 22594
rect 27358 22542 27410 22594
rect 27410 22542 27412 22594
rect 27356 22540 27412 22542
rect 27916 23100 27972 23156
rect 27356 21980 27412 22036
rect 27468 21868 27524 21924
rect 27580 21586 27636 21588
rect 27580 21534 27582 21586
rect 27582 21534 27634 21586
rect 27634 21534 27636 21586
rect 27580 21532 27636 21534
rect 28364 26796 28420 26852
rect 28252 26514 28308 26516
rect 28252 26462 28254 26514
rect 28254 26462 28306 26514
rect 28306 26462 28308 26514
rect 28252 26460 28308 26462
rect 28140 25340 28196 25396
rect 28252 17724 28308 17780
rect 27244 15986 27300 15988
rect 27244 15934 27246 15986
rect 27246 15934 27298 15986
rect 27298 15934 27300 15986
rect 27244 15932 27300 15934
rect 28588 26684 28644 26740
rect 29484 41020 29540 41076
rect 31388 49196 31444 49252
rect 31164 48300 31220 48356
rect 31724 47404 31780 47460
rect 31724 45724 31780 45780
rect 31500 44322 31556 44324
rect 31500 44270 31502 44322
rect 31502 44270 31554 44322
rect 31554 44270 31556 44322
rect 31500 44268 31556 44270
rect 31388 42700 31444 42756
rect 32060 49026 32116 49028
rect 32060 48974 32062 49026
rect 32062 48974 32114 49026
rect 32114 48974 32116 49026
rect 32060 48972 32116 48974
rect 31948 48242 32004 48244
rect 31948 48190 31950 48242
rect 31950 48190 32002 48242
rect 32002 48190 32004 48242
rect 31948 48188 32004 48190
rect 33404 52220 33460 52276
rect 32956 51996 33012 52052
rect 32620 48300 32676 48356
rect 32732 48860 32788 48916
rect 32284 48188 32340 48244
rect 32060 45612 32116 45668
rect 32620 48130 32676 48132
rect 32620 48078 32622 48130
rect 32622 48078 32674 48130
rect 32674 48078 32676 48130
rect 32620 48076 32676 48078
rect 32844 47458 32900 47460
rect 32844 47406 32846 47458
rect 32846 47406 32898 47458
rect 32898 47406 32900 47458
rect 32844 47404 32900 47406
rect 32508 45276 32564 45332
rect 32284 44380 32340 44436
rect 32396 43372 32452 43428
rect 31164 41692 31220 41748
rect 30604 40684 30660 40740
rect 30604 40460 30660 40516
rect 32620 44828 32676 44884
rect 33180 49868 33236 49924
rect 33068 48076 33124 48132
rect 32844 44268 32900 44324
rect 33068 43650 33124 43652
rect 33068 43598 33070 43650
rect 33070 43598 33122 43650
rect 33122 43598 33124 43650
rect 33068 43596 33124 43598
rect 34412 52274 34468 52276
rect 34412 52222 34414 52274
rect 34414 52222 34466 52274
rect 34466 52222 34468 52274
rect 34412 52220 34468 52222
rect 33404 48972 33460 49028
rect 33516 48748 33572 48804
rect 33740 45330 33796 45332
rect 33740 45278 33742 45330
rect 33742 45278 33794 45330
rect 33794 45278 33796 45330
rect 33740 45276 33796 45278
rect 33740 44380 33796 44436
rect 33628 44044 33684 44100
rect 33292 43372 33348 43428
rect 37324 53564 37380 53620
rect 34636 48860 34692 48916
rect 33964 45612 34020 45668
rect 32396 41692 32452 41748
rect 31724 40460 31780 40516
rect 30940 39900 30996 39956
rect 31164 40348 31220 40404
rect 29932 39788 29988 39844
rect 31948 40348 32004 40404
rect 32172 40236 32228 40292
rect 32620 41804 32676 41860
rect 32732 41186 32788 41188
rect 32732 41134 32734 41186
rect 32734 41134 32786 41186
rect 32786 41134 32788 41186
rect 32732 41132 32788 41134
rect 32284 40460 32340 40516
rect 32060 39900 32116 39956
rect 31164 38834 31220 38836
rect 31164 38782 31166 38834
rect 31166 38782 31218 38834
rect 31218 38782 31220 38834
rect 31164 38780 31220 38782
rect 31948 38946 32004 38948
rect 31948 38894 31950 38946
rect 31950 38894 32002 38946
rect 32002 38894 32004 38946
rect 31948 38892 32004 38894
rect 30940 38108 30996 38164
rect 30828 37938 30884 37940
rect 30828 37886 30830 37938
rect 30830 37886 30882 37938
rect 30882 37886 30884 37938
rect 30828 37884 30884 37886
rect 29484 37266 29540 37268
rect 29484 37214 29486 37266
rect 29486 37214 29538 37266
rect 29538 37214 29540 37266
rect 29484 37212 29540 37214
rect 29596 36876 29652 36932
rect 29932 36204 29988 36260
rect 30604 33346 30660 33348
rect 30604 33294 30606 33346
rect 30606 33294 30658 33346
rect 30658 33294 30660 33346
rect 30604 33292 30660 33294
rect 32620 39788 32676 39844
rect 31164 37938 31220 37940
rect 31164 37886 31166 37938
rect 31166 37886 31218 37938
rect 31218 37886 31220 37938
rect 31164 37884 31220 37886
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35756 52220 35812 52276
rect 35420 52050 35476 52052
rect 35420 51998 35422 52050
rect 35422 51998 35474 52050
rect 35474 51998 35476 52050
rect 35420 51996 35476 51998
rect 34860 48748 34916 48804
rect 34972 51436 35028 51492
rect 34076 41746 34132 41748
rect 34076 41694 34078 41746
rect 34078 41694 34130 41746
rect 34130 41694 34132 41746
rect 34076 41692 34132 41694
rect 33964 40572 34020 40628
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 50764 35252 50820
rect 35308 49922 35364 49924
rect 35308 49870 35310 49922
rect 35310 49870 35362 49922
rect 35362 49870 35364 49922
rect 35308 49868 35364 49870
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35420 48188 35476 48244
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 33516 40236 33572 40292
rect 33292 38892 33348 38948
rect 34524 40236 34580 40292
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34972 41692 35028 41748
rect 36652 53004 36708 53060
rect 35868 50764 35924 50820
rect 36428 52780 36484 52836
rect 36316 49868 36372 49924
rect 36092 48242 36148 48244
rect 36092 48190 36094 48242
rect 36094 48190 36146 48242
rect 36146 48190 36148 48242
rect 36092 48188 36148 48190
rect 35980 47404 36036 47460
rect 36540 49532 36596 49588
rect 36764 48242 36820 48244
rect 36764 48190 36766 48242
rect 36766 48190 36818 48242
rect 36818 48190 36820 48242
rect 36764 48188 36820 48190
rect 36764 47404 36820 47460
rect 36988 49922 37044 49924
rect 36988 49870 36990 49922
rect 36990 49870 37042 49922
rect 37042 49870 37044 49922
rect 36988 49868 37044 49870
rect 39564 53618 39620 53620
rect 39564 53566 39566 53618
rect 39566 53566 39618 53618
rect 39618 53566 39620 53618
rect 39564 53564 39620 53566
rect 38668 53058 38724 53060
rect 38668 53006 38670 53058
rect 38670 53006 38722 53058
rect 38722 53006 38724 53058
rect 38668 53004 38724 53006
rect 37660 52834 37716 52836
rect 37660 52782 37662 52834
rect 37662 52782 37714 52834
rect 37714 52782 37716 52834
rect 37660 52780 37716 52782
rect 37996 52274 38052 52276
rect 37996 52222 37998 52274
rect 37998 52222 38050 52274
rect 38050 52222 38052 52274
rect 37996 52220 38052 52222
rect 39452 52220 39508 52276
rect 37772 51490 37828 51492
rect 37772 51438 37774 51490
rect 37774 51438 37826 51490
rect 37826 51438 37828 51490
rect 37772 51436 37828 51438
rect 39004 50652 39060 50708
rect 38220 50540 38276 50596
rect 35980 44044 36036 44100
rect 37436 45106 37492 45108
rect 37436 45054 37438 45106
rect 37438 45054 37490 45106
rect 37490 45054 37492 45106
rect 37436 45052 37492 45054
rect 37996 48188 38052 48244
rect 36428 44268 36484 44324
rect 36988 44322 37044 44324
rect 36988 44270 36990 44322
rect 36990 44270 37042 44322
rect 37042 44270 37044 44322
rect 36988 44268 37044 44270
rect 36540 43538 36596 43540
rect 36540 43486 36542 43538
rect 36542 43486 36594 43538
rect 36594 43486 36596 43538
rect 36540 43484 36596 43486
rect 36876 42754 36932 42756
rect 36876 42702 36878 42754
rect 36878 42702 36930 42754
rect 36930 42702 36932 42754
rect 36876 42700 36932 42702
rect 38220 47180 38276 47236
rect 39116 49532 39172 49588
rect 39116 48972 39172 49028
rect 38892 48076 38948 48132
rect 37660 43932 37716 43988
rect 36092 41692 36148 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 36316 42028 36372 42084
rect 35196 40962 35252 40964
rect 35196 40910 35198 40962
rect 35198 40910 35250 40962
rect 35250 40910 35252 40962
rect 35196 40908 35252 40910
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 33292 38668 33348 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 38274 35140 38276
rect 35084 38222 35086 38274
rect 35086 38222 35138 38274
rect 35138 38222 35140 38274
rect 35084 38220 35140 38222
rect 33404 37884 33460 37940
rect 31164 36540 31220 36596
rect 30156 33234 30212 33236
rect 30156 33182 30158 33234
rect 30158 33182 30210 33234
rect 30210 33182 30212 33234
rect 30156 33180 30212 33182
rect 29372 31836 29428 31892
rect 33404 37378 33460 37380
rect 33404 37326 33406 37378
rect 33406 37326 33458 37378
rect 33458 37326 33460 37378
rect 33404 37324 33460 37326
rect 34188 37378 34244 37380
rect 34188 37326 34190 37378
rect 34190 37326 34242 37378
rect 34242 37326 34244 37378
rect 34188 37324 34244 37326
rect 32732 36482 32788 36484
rect 32732 36430 32734 36482
rect 32734 36430 32786 36482
rect 32786 36430 32788 36482
rect 32732 36428 32788 36430
rect 33516 36540 33572 36596
rect 33068 36482 33124 36484
rect 33068 36430 33070 36482
rect 33070 36430 33122 36482
rect 33122 36430 33124 36482
rect 33068 36428 33124 36430
rect 31836 35868 31892 35924
rect 33068 35810 33124 35812
rect 33068 35758 33070 35810
rect 33070 35758 33122 35810
rect 33122 35758 33124 35810
rect 33068 35756 33124 35758
rect 33404 35810 33460 35812
rect 33404 35758 33406 35810
rect 33406 35758 33458 35810
rect 33458 35758 33460 35810
rect 33404 35756 33460 35758
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34076 35810 34132 35812
rect 34076 35758 34078 35810
rect 34078 35758 34130 35810
rect 34130 35758 34132 35810
rect 34076 35756 34132 35758
rect 34860 36428 34916 36484
rect 31276 34354 31332 34356
rect 31276 34302 31278 34354
rect 31278 34302 31330 34354
rect 31330 34302 31332 34354
rect 31276 34300 31332 34302
rect 31164 31836 31220 31892
rect 29036 30828 29092 30884
rect 29260 31778 29316 31780
rect 29260 31726 29262 31778
rect 29262 31726 29314 31778
rect 29314 31726 29316 31778
rect 29260 31724 29316 31726
rect 29260 30210 29316 30212
rect 29260 30158 29262 30210
rect 29262 30158 29314 30210
rect 29314 30158 29316 30210
rect 29260 30156 29316 30158
rect 28924 29202 28980 29204
rect 28924 29150 28926 29202
rect 28926 29150 28978 29202
rect 28978 29150 28980 29202
rect 28924 29148 28980 29150
rect 29708 29538 29764 29540
rect 29708 29486 29710 29538
rect 29710 29486 29762 29538
rect 29762 29486 29764 29538
rect 29708 29484 29764 29486
rect 29708 28642 29764 28644
rect 29708 28590 29710 28642
rect 29710 28590 29762 28642
rect 29762 28590 29764 28642
rect 29708 28588 29764 28590
rect 29932 28476 29988 28532
rect 29596 27916 29652 27972
rect 30156 28364 30212 28420
rect 28700 24220 28756 24276
rect 29372 26684 29428 26740
rect 29260 25452 29316 25508
rect 29372 26460 29428 26516
rect 29148 25228 29204 25284
rect 29484 25676 29540 25732
rect 28924 24556 28980 24612
rect 29148 24050 29204 24052
rect 29148 23998 29150 24050
rect 29150 23998 29202 24050
rect 29202 23998 29204 24050
rect 29148 23996 29204 23998
rect 29148 23154 29204 23156
rect 29148 23102 29150 23154
rect 29150 23102 29202 23154
rect 29202 23102 29204 23154
rect 29148 23100 29204 23102
rect 28588 22258 28644 22260
rect 28588 22206 28590 22258
rect 28590 22206 28642 22258
rect 28642 22206 28644 22258
rect 28588 22204 28644 22206
rect 28476 18508 28532 18564
rect 28812 20300 28868 20356
rect 29148 22764 29204 22820
rect 29148 22540 29204 22596
rect 29708 25564 29764 25620
rect 30044 25228 30100 25284
rect 30044 24556 30100 24612
rect 29596 23548 29652 23604
rect 29708 24220 29764 24276
rect 29484 21532 29540 21588
rect 29596 20188 29652 20244
rect 29932 23100 29988 23156
rect 30156 22764 30212 22820
rect 30156 22204 30212 22260
rect 30492 29484 30548 29540
rect 31164 29372 31220 29428
rect 30716 28754 30772 28756
rect 30716 28702 30718 28754
rect 30718 28702 30770 28754
rect 30770 28702 30772 28754
rect 30716 28700 30772 28702
rect 30940 28418 30996 28420
rect 30940 28366 30942 28418
rect 30942 28366 30994 28418
rect 30994 28366 30996 28418
rect 30940 28364 30996 28366
rect 30380 25676 30436 25732
rect 30828 25564 30884 25620
rect 30380 25340 30436 25396
rect 30492 22988 30548 23044
rect 30492 22204 30548 22260
rect 30604 23548 30660 23604
rect 30156 18508 30212 18564
rect 30940 25282 30996 25284
rect 30940 25230 30942 25282
rect 30942 25230 30994 25282
rect 30994 25230 30996 25282
rect 30940 25228 30996 25230
rect 30940 24722 30996 24724
rect 30940 24670 30942 24722
rect 30942 24670 30994 24722
rect 30994 24670 30996 24722
rect 30940 24668 30996 24670
rect 31836 35196 31892 35252
rect 32396 35644 32452 35700
rect 32060 34242 32116 34244
rect 32060 34190 32062 34242
rect 32062 34190 32114 34242
rect 32114 34190 32116 34242
rect 32060 34188 32116 34190
rect 36652 41244 36708 41300
rect 36988 41692 37044 41748
rect 37100 40962 37156 40964
rect 37100 40910 37102 40962
rect 37102 40910 37154 40962
rect 37154 40910 37156 40962
rect 37100 40908 37156 40910
rect 37212 40626 37268 40628
rect 37212 40574 37214 40626
rect 37214 40574 37266 40626
rect 37266 40574 37268 40626
rect 37212 40572 37268 40574
rect 40460 50428 40516 50484
rect 40460 47570 40516 47572
rect 40460 47518 40462 47570
rect 40462 47518 40514 47570
rect 40514 47518 40516 47570
rect 40460 47516 40516 47518
rect 40348 46786 40404 46788
rect 40348 46734 40350 46786
rect 40350 46734 40402 46786
rect 40402 46734 40404 46786
rect 40348 46732 40404 46734
rect 40684 51996 40740 52052
rect 40796 50540 40852 50596
rect 41356 50092 41412 50148
rect 41132 48802 41188 48804
rect 41132 48750 41134 48802
rect 41134 48750 41186 48802
rect 41186 48750 41188 48802
rect 41132 48748 41188 48750
rect 41356 48860 41412 48916
rect 40908 48130 40964 48132
rect 40908 48078 40910 48130
rect 40910 48078 40962 48130
rect 40962 48078 40964 48130
rect 40908 48076 40964 48078
rect 40796 47516 40852 47572
rect 41020 45948 41076 46004
rect 39900 45164 39956 45220
rect 39004 42700 39060 42756
rect 39004 41916 39060 41972
rect 38220 41298 38276 41300
rect 38220 41246 38222 41298
rect 38222 41246 38274 41298
rect 38274 41246 38276 41298
rect 38220 41244 38276 41246
rect 39564 41970 39620 41972
rect 39564 41918 39566 41970
rect 39566 41918 39618 41970
rect 39618 41918 39620 41970
rect 39564 41916 39620 41918
rect 41244 46732 41300 46788
rect 42700 54402 42756 54404
rect 42700 54350 42702 54402
rect 42702 54350 42754 54402
rect 42754 54350 42756 54402
rect 42700 54348 42756 54350
rect 43036 53788 43092 53844
rect 42364 52220 42420 52276
rect 41692 52108 41748 52164
rect 41580 49196 41636 49252
rect 41804 52050 41860 52052
rect 41804 51998 41806 52050
rect 41806 51998 41858 52050
rect 41858 51998 41860 52050
rect 41804 51996 41860 51998
rect 42476 50316 42532 50372
rect 41916 48972 41972 49028
rect 42252 48914 42308 48916
rect 42252 48862 42254 48914
rect 42254 48862 42306 48914
rect 42306 48862 42308 48914
rect 42252 48860 42308 48862
rect 41916 47516 41972 47572
rect 42476 47964 42532 48020
rect 42028 47180 42084 47236
rect 42252 47180 42308 47236
rect 40908 43820 40964 43876
rect 41020 43484 41076 43540
rect 40796 41970 40852 41972
rect 40796 41918 40798 41970
rect 40798 41918 40850 41970
rect 40850 41918 40852 41970
rect 40796 41916 40852 41918
rect 40012 41244 40068 41300
rect 38556 41074 38612 41076
rect 38556 41022 38558 41074
rect 38558 41022 38610 41074
rect 38610 41022 38612 41074
rect 38556 41020 38612 41022
rect 40124 41020 40180 41076
rect 38556 40348 38612 40404
rect 38444 40290 38500 40292
rect 38444 40238 38446 40290
rect 38446 40238 38498 40290
rect 38498 40238 38500 40290
rect 38444 40236 38500 40238
rect 37436 38892 37492 38948
rect 37436 38162 37492 38164
rect 37436 38110 37438 38162
rect 37438 38110 37490 38162
rect 37490 38110 37492 38162
rect 37436 38108 37492 38110
rect 37436 37324 37492 37380
rect 36540 36706 36596 36708
rect 36540 36654 36542 36706
rect 36542 36654 36594 36706
rect 36594 36654 36596 36706
rect 36540 36652 36596 36654
rect 35644 36428 35700 36484
rect 35980 36316 36036 36372
rect 36988 36370 37044 36372
rect 36988 36318 36990 36370
rect 36990 36318 37042 36370
rect 37042 36318 37044 36370
rect 36988 36316 37044 36318
rect 35532 35980 35588 36036
rect 31836 33292 31892 33348
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 37996 38108 38052 38164
rect 38556 37212 38612 37268
rect 40908 39618 40964 39620
rect 40908 39566 40910 39618
rect 40910 39566 40962 39618
rect 40962 39566 40964 39618
rect 40908 39564 40964 39566
rect 40908 39116 40964 39172
rect 40236 38892 40292 38948
rect 41804 45948 41860 46004
rect 41468 45218 41524 45220
rect 41468 45166 41470 45218
rect 41470 45166 41522 45218
rect 41522 45166 41524 45218
rect 41468 45164 41524 45166
rect 41468 44940 41524 44996
rect 41692 44156 41748 44212
rect 41468 42812 41524 42868
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 45836 53842 45892 53844
rect 45836 53790 45838 53842
rect 45838 53790 45890 53842
rect 45890 53790 45892 53842
rect 45836 53788 45892 53790
rect 43708 52108 43764 52164
rect 44492 53564 44548 53620
rect 42924 48914 42980 48916
rect 42924 48862 42926 48914
rect 42926 48862 42978 48914
rect 42978 48862 42980 48914
rect 42924 48860 42980 48862
rect 42812 48802 42868 48804
rect 42812 48750 42814 48802
rect 42814 48750 42866 48802
rect 42866 48750 42868 48802
rect 42812 48748 42868 48750
rect 43148 47964 43204 48020
rect 43484 48860 43540 48916
rect 42924 47234 42980 47236
rect 42924 47182 42926 47234
rect 42926 47182 42978 47234
rect 42978 47182 42980 47234
rect 42924 47180 42980 47182
rect 42924 45612 42980 45668
rect 43148 45218 43204 45220
rect 43148 45166 43150 45218
rect 43150 45166 43202 45218
rect 43202 45166 43204 45218
rect 43148 45164 43204 45166
rect 42700 44940 42756 44996
rect 43596 44940 43652 44996
rect 43596 44210 43652 44212
rect 43596 44158 43598 44210
rect 43598 44158 43650 44210
rect 43650 44158 43652 44210
rect 43596 44156 43652 44158
rect 42812 43932 42868 43988
rect 44268 48188 44324 48244
rect 44380 47180 44436 47236
rect 47068 53618 47124 53620
rect 47068 53566 47070 53618
rect 47070 53566 47122 53618
rect 47122 53566 47124 53618
rect 47068 53564 47124 53566
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 44604 53004 44660 53060
rect 45948 53058 46004 53060
rect 45948 53006 45950 53058
rect 45950 53006 46002 53058
rect 46002 53006 46004 53058
rect 45948 53004 46004 53006
rect 44940 50316 44996 50372
rect 45948 51436 46004 51492
rect 45836 50706 45892 50708
rect 45836 50654 45838 50706
rect 45838 50654 45890 50706
rect 45890 50654 45892 50706
rect 45836 50652 45892 50654
rect 45724 50092 45780 50148
rect 46060 50652 46116 50708
rect 45388 49868 45444 49924
rect 45612 49756 45668 49812
rect 44716 49196 44772 49252
rect 44828 49644 44884 49700
rect 45388 49532 45444 49588
rect 44828 48188 44884 48244
rect 44716 46732 44772 46788
rect 45612 49084 45668 49140
rect 45612 48242 45668 48244
rect 45612 48190 45614 48242
rect 45614 48190 45666 48242
rect 45666 48190 45668 48242
rect 45612 48188 45668 48190
rect 44940 47068 44996 47124
rect 44828 45948 44884 46004
rect 42588 42812 42644 42868
rect 41804 42028 41860 42084
rect 43372 41298 43428 41300
rect 43372 41246 43374 41298
rect 43374 41246 43426 41298
rect 43426 41246 43428 41298
rect 43372 41244 43428 41246
rect 42476 41186 42532 41188
rect 42476 41134 42478 41186
rect 42478 41134 42530 41186
rect 42530 41134 42532 41186
rect 42476 41132 42532 41134
rect 43148 40908 43204 40964
rect 42700 40348 42756 40404
rect 42812 40460 42868 40516
rect 41692 39564 41748 39620
rect 41244 39116 41300 39172
rect 41804 39116 41860 39172
rect 41580 39004 41636 39060
rect 39676 38444 39732 38500
rect 39452 37436 39508 37492
rect 37772 36482 37828 36484
rect 37772 36430 37774 36482
rect 37774 36430 37826 36482
rect 37826 36430 37828 36482
rect 37772 36428 37828 36430
rect 38556 34972 38612 35028
rect 35196 34860 35252 34916
rect 37884 34914 37940 34916
rect 37884 34862 37886 34914
rect 37886 34862 37938 34914
rect 37938 34862 37940 34914
rect 37884 34860 37940 34862
rect 36092 34412 36148 34468
rect 32956 33906 33012 33908
rect 32956 33854 32958 33906
rect 32958 33854 33010 33906
rect 33010 33854 33012 33906
rect 32956 33852 33012 33854
rect 32508 33404 32564 33460
rect 31500 28476 31556 28532
rect 31724 28418 31780 28420
rect 31724 28366 31726 28418
rect 31726 28366 31778 28418
rect 31778 28366 31780 28418
rect 31724 28364 31780 28366
rect 36540 34412 36596 34468
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 33458 35140 33460
rect 35084 33406 35086 33458
rect 35086 33406 35138 33458
rect 35138 33406 35140 33458
rect 35084 33404 35140 33406
rect 35644 33458 35700 33460
rect 35644 33406 35646 33458
rect 35646 33406 35698 33458
rect 35698 33406 35700 33458
rect 35644 33404 35700 33406
rect 36428 33404 36484 33460
rect 34524 33180 34580 33236
rect 32172 31724 32228 31780
rect 32172 30882 32228 30884
rect 32172 30830 32174 30882
rect 32174 30830 32226 30882
rect 32226 30830 32228 30882
rect 32172 30828 32228 30830
rect 32172 29986 32228 29988
rect 32172 29934 32174 29986
rect 32174 29934 32226 29986
rect 32226 29934 32228 29986
rect 32172 29932 32228 29934
rect 32060 29596 32116 29652
rect 32060 29426 32116 29428
rect 32060 29374 32062 29426
rect 32062 29374 32114 29426
rect 32114 29374 32116 29426
rect 32060 29372 32116 29374
rect 31836 28028 31892 28084
rect 31388 27132 31444 27188
rect 31388 25506 31444 25508
rect 31388 25454 31390 25506
rect 31390 25454 31442 25506
rect 31442 25454 31444 25506
rect 31388 25452 31444 25454
rect 31388 24780 31444 24836
rect 32060 23660 32116 23716
rect 32060 23212 32116 23268
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 33740 31836 33796 31892
rect 33404 31778 33460 31780
rect 33404 31726 33406 31778
rect 33406 31726 33458 31778
rect 33458 31726 33460 31778
rect 33404 31724 33460 31726
rect 33068 30268 33124 30324
rect 33180 30828 33236 30884
rect 32620 29260 32676 29316
rect 32396 28476 32452 28532
rect 32396 27858 32452 27860
rect 32396 27806 32398 27858
rect 32398 27806 32450 27858
rect 32450 27806 32452 27858
rect 32396 27804 32452 27806
rect 32508 28028 32564 28084
rect 32396 23324 32452 23380
rect 31612 21532 31668 21588
rect 32284 22092 32340 22148
rect 31276 20300 31332 20356
rect 31164 20188 31220 20244
rect 32396 21756 32452 21812
rect 32396 21532 32452 21588
rect 31836 18172 31892 18228
rect 32732 26850 32788 26852
rect 32732 26798 32734 26850
rect 32734 26798 32786 26850
rect 32786 26798 32788 26850
rect 32732 26796 32788 26798
rect 32508 21420 32564 21476
rect 32620 20412 32676 20468
rect 33068 29932 33124 29988
rect 33068 29260 33124 29316
rect 33516 30210 33572 30212
rect 33516 30158 33518 30210
rect 33518 30158 33570 30210
rect 33570 30158 33572 30210
rect 33516 30156 33572 30158
rect 33292 29372 33348 29428
rect 33404 28700 33460 28756
rect 33740 29596 33796 29652
rect 33964 28700 34020 28756
rect 34636 29260 34692 29316
rect 33628 28364 33684 28420
rect 32956 23548 33012 23604
rect 33068 23266 33124 23268
rect 33068 23214 33070 23266
rect 33070 23214 33122 23266
rect 33122 23214 33124 23266
rect 33068 23212 33124 23214
rect 33292 22988 33348 23044
rect 33068 22370 33124 22372
rect 33068 22318 33070 22370
rect 33070 22318 33122 22370
rect 33122 22318 33124 22370
rect 33068 22316 33124 22318
rect 33404 21532 33460 21588
rect 33404 21308 33460 21364
rect 32732 16940 32788 16996
rect 33852 27858 33908 27860
rect 33852 27806 33854 27858
rect 33854 27806 33906 27858
rect 33906 27806 33908 27858
rect 33852 27804 33908 27806
rect 33628 26796 33684 26852
rect 33740 26514 33796 26516
rect 33740 26462 33742 26514
rect 33742 26462 33794 26514
rect 33794 26462 33796 26514
rect 33740 26460 33796 26462
rect 33964 27186 34020 27188
rect 33964 27134 33966 27186
rect 33966 27134 34018 27186
rect 34018 27134 34020 27186
rect 33964 27132 34020 27134
rect 34524 26908 34580 26964
rect 34076 24834 34132 24836
rect 34076 24782 34078 24834
rect 34078 24782 34130 24834
rect 34130 24782 34132 24834
rect 34076 24780 34132 24782
rect 34748 26684 34804 26740
rect 36092 33180 36148 33236
rect 37436 34130 37492 34132
rect 37436 34078 37438 34130
rect 37438 34078 37490 34130
rect 37490 34078 37492 34130
rect 37436 34076 37492 34078
rect 36540 33292 36596 33348
rect 36092 32562 36148 32564
rect 36092 32510 36094 32562
rect 36094 32510 36146 32562
rect 36146 32510 36148 32562
rect 36092 32508 36148 32510
rect 37324 33180 37380 33236
rect 36988 31890 37044 31892
rect 36988 31838 36990 31890
rect 36990 31838 37042 31890
rect 37042 31838 37044 31890
rect 36988 31836 37044 31838
rect 36540 31778 36596 31780
rect 36540 31726 36542 31778
rect 36542 31726 36594 31778
rect 36594 31726 36596 31778
rect 36540 31724 36596 31726
rect 37436 32562 37492 32564
rect 37436 32510 37438 32562
rect 37438 32510 37490 32562
rect 37490 32510 37492 32562
rect 37436 32508 37492 32510
rect 38892 36428 38948 36484
rect 39676 36540 39732 36596
rect 40348 37154 40404 37156
rect 40348 37102 40350 37154
rect 40350 37102 40402 37154
rect 40402 37102 40404 37154
rect 40348 37100 40404 37102
rect 41804 37996 41860 38052
rect 41692 36706 41748 36708
rect 41692 36654 41694 36706
rect 41694 36654 41746 36706
rect 41746 36654 41748 36706
rect 41692 36652 41748 36654
rect 41020 36540 41076 36596
rect 40124 36316 40180 36372
rect 40908 36370 40964 36372
rect 40908 36318 40910 36370
rect 40910 36318 40962 36370
rect 40962 36318 40964 36370
rect 40908 36316 40964 36318
rect 41468 35698 41524 35700
rect 41468 35646 41470 35698
rect 41470 35646 41522 35698
rect 41522 35646 41524 35698
rect 41468 35644 41524 35646
rect 41132 35084 41188 35140
rect 42700 38780 42756 38836
rect 42924 38220 42980 38276
rect 43036 38668 43092 38724
rect 42140 37884 42196 37940
rect 42924 37938 42980 37940
rect 42924 37886 42926 37938
rect 42926 37886 42978 37938
rect 42978 37886 42980 37938
rect 42924 37884 42980 37886
rect 41916 36876 41972 36932
rect 43036 36876 43092 36932
rect 43708 41074 43764 41076
rect 43708 41022 43710 41074
rect 43710 41022 43762 41074
rect 43762 41022 43764 41074
rect 43708 41020 43764 41022
rect 43708 40796 43764 40852
rect 46172 49698 46228 49700
rect 46172 49646 46174 49698
rect 46174 49646 46226 49698
rect 46226 49646 46228 49698
rect 46172 49644 46228 49646
rect 47068 50482 47124 50484
rect 47068 50430 47070 50482
rect 47070 50430 47122 50482
rect 47122 50430 47124 50482
rect 47068 50428 47124 50430
rect 46844 49922 46900 49924
rect 46844 49870 46846 49922
rect 46846 49870 46898 49922
rect 46898 49870 46900 49922
rect 46844 49868 46900 49870
rect 46396 49644 46452 49700
rect 47068 49644 47124 49700
rect 46396 48860 46452 48916
rect 45388 45276 45444 45332
rect 46508 48748 46564 48804
rect 45164 45164 45220 45220
rect 45724 45666 45780 45668
rect 45724 45614 45726 45666
rect 45726 45614 45778 45666
rect 45778 45614 45780 45666
rect 45724 45612 45780 45614
rect 46172 45388 46228 45444
rect 46284 47068 46340 47124
rect 46844 46844 46900 46900
rect 47292 45330 47348 45332
rect 47292 45278 47294 45330
rect 47294 45278 47346 45330
rect 47346 45278 47348 45330
rect 47292 45276 47348 45278
rect 45388 44156 45444 44212
rect 45388 43932 45444 43988
rect 44940 42754 44996 42756
rect 44940 42702 44942 42754
rect 44942 42702 44994 42754
rect 44994 42702 44996 42754
rect 44940 42700 44996 42702
rect 43932 41244 43988 41300
rect 43708 39564 43764 39620
rect 44044 40796 44100 40852
rect 44940 40402 44996 40404
rect 44940 40350 44942 40402
rect 44942 40350 44994 40402
rect 44994 40350 44996 40402
rect 44940 40348 44996 40350
rect 44492 39676 44548 39732
rect 44380 38780 44436 38836
rect 43148 37884 43204 37940
rect 43820 37884 43876 37940
rect 43148 37100 43204 37156
rect 42028 36594 42084 36596
rect 42028 36542 42030 36594
rect 42030 36542 42082 36594
rect 42082 36542 42084 36594
rect 42028 36540 42084 36542
rect 42812 36594 42868 36596
rect 42812 36542 42814 36594
rect 42814 36542 42866 36594
rect 42866 36542 42868 36594
rect 42812 36540 42868 36542
rect 45164 43372 45220 43428
rect 46508 44994 46564 44996
rect 46508 44942 46510 44994
rect 46510 44942 46562 44994
rect 46562 44942 46564 44994
rect 46508 44940 46564 44942
rect 47180 44994 47236 44996
rect 47180 44942 47182 44994
rect 47182 44942 47234 44994
rect 47234 44942 47236 44994
rect 47180 44940 47236 44942
rect 46620 44322 46676 44324
rect 46620 44270 46622 44322
rect 46622 44270 46674 44322
rect 46674 44270 46676 44322
rect 46620 44268 46676 44270
rect 46396 43932 46452 43988
rect 45948 43820 46004 43876
rect 48412 49756 48468 49812
rect 48636 51996 48692 52052
rect 47516 49698 47572 49700
rect 47516 49646 47518 49698
rect 47518 49646 47570 49698
rect 47570 49646 47572 49698
rect 47516 49644 47572 49646
rect 47964 49644 48020 49700
rect 47740 48636 47796 48692
rect 47628 46844 47684 46900
rect 48412 48860 48468 48916
rect 48076 47068 48132 47124
rect 48636 50706 48692 50708
rect 48636 50654 48638 50706
rect 48638 50654 48690 50706
rect 48690 50654 48692 50706
rect 48636 50652 48692 50654
rect 48636 50428 48692 50484
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 51100 52108 51156 52164
rect 49420 49698 49476 49700
rect 49420 49646 49422 49698
rect 49422 49646 49474 49698
rect 49474 49646 49476 49698
rect 49420 49644 49476 49646
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50764 51490 50820 51492
rect 50764 51438 50766 51490
rect 50766 51438 50818 51490
rect 50818 51438 50820 51490
rect 50764 51436 50820 51438
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49980 49698 50036 49700
rect 49980 49646 49982 49698
rect 49982 49646 50034 49698
rect 50034 49646 50036 49698
rect 49980 49644 50036 49646
rect 49868 49532 49924 49588
rect 49868 48748 49924 48804
rect 49756 48636 49812 48692
rect 49532 48076 49588 48132
rect 49308 47180 49364 47236
rect 49420 47404 49476 47460
rect 48524 47068 48580 47124
rect 49308 45948 49364 46004
rect 48188 45330 48244 45332
rect 48188 45278 48190 45330
rect 48190 45278 48242 45330
rect 48242 45278 48244 45330
rect 48188 45276 48244 45278
rect 49644 46172 49700 46228
rect 49084 43820 49140 43876
rect 48972 43708 49028 43764
rect 47404 43484 47460 43540
rect 47740 43650 47796 43652
rect 47740 43598 47742 43650
rect 47742 43598 47794 43650
rect 47794 43598 47796 43650
rect 47740 43596 47796 43598
rect 45276 41970 45332 41972
rect 45276 41918 45278 41970
rect 45278 41918 45330 41970
rect 45330 41918 45332 41970
rect 45276 41916 45332 41918
rect 45500 41298 45556 41300
rect 45500 41246 45502 41298
rect 45502 41246 45554 41298
rect 45554 41246 45556 41298
rect 45500 41244 45556 41246
rect 48188 43650 48244 43652
rect 48188 43598 48190 43650
rect 48190 43598 48242 43650
rect 48242 43598 48244 43650
rect 48188 43596 48244 43598
rect 48860 43426 48916 43428
rect 48860 43374 48862 43426
rect 48862 43374 48914 43426
rect 48914 43374 48916 43426
rect 48860 43372 48916 43374
rect 47740 42700 47796 42756
rect 46508 42476 46564 42532
rect 46172 41298 46228 41300
rect 46172 41246 46174 41298
rect 46174 41246 46226 41298
rect 46226 41246 46228 41298
rect 46172 41244 46228 41246
rect 47628 42530 47684 42532
rect 47628 42478 47630 42530
rect 47630 42478 47682 42530
rect 47682 42478 47684 42530
rect 47628 42476 47684 42478
rect 46844 41298 46900 41300
rect 46844 41246 46846 41298
rect 46846 41246 46898 41298
rect 46898 41246 46900 41298
rect 46844 41244 46900 41246
rect 45164 41074 45220 41076
rect 45164 41022 45166 41074
rect 45166 41022 45218 41074
rect 45218 41022 45220 41074
rect 45164 41020 45220 41022
rect 48300 43148 48356 43204
rect 48412 42642 48468 42644
rect 48412 42590 48414 42642
rect 48414 42590 48466 42642
rect 48466 42590 48468 42642
rect 48412 42588 48468 42590
rect 49196 43372 49252 43428
rect 48076 41186 48132 41188
rect 48076 41134 48078 41186
rect 48078 41134 48130 41186
rect 48130 41134 48132 41186
rect 48076 41132 48132 41134
rect 45724 40796 45780 40852
rect 45388 39618 45444 39620
rect 45388 39566 45390 39618
rect 45390 39566 45442 39618
rect 45442 39566 45444 39618
rect 45388 39564 45444 39566
rect 45388 39058 45444 39060
rect 45388 39006 45390 39058
rect 45390 39006 45442 39058
rect 45442 39006 45444 39058
rect 45388 39004 45444 39006
rect 47068 38946 47124 38948
rect 47068 38894 47070 38946
rect 47070 38894 47122 38946
rect 47122 38894 47124 38946
rect 47068 38892 47124 38894
rect 45052 38780 45108 38836
rect 44380 36428 44436 36484
rect 45388 38220 45444 38276
rect 44828 37100 44884 37156
rect 45500 37884 45556 37940
rect 45500 37324 45556 37380
rect 44828 36540 44884 36596
rect 44492 35922 44548 35924
rect 44492 35870 44494 35922
rect 44494 35870 44546 35922
rect 44546 35870 44548 35922
rect 44492 35868 44548 35870
rect 45276 36764 45332 36820
rect 47964 40626 48020 40628
rect 47964 40574 47966 40626
rect 47966 40574 48018 40626
rect 48018 40574 48020 40626
rect 47964 40572 48020 40574
rect 49868 45276 49924 45332
rect 49868 44434 49924 44436
rect 49868 44382 49870 44434
rect 49870 44382 49922 44434
rect 49922 44382 49924 44434
rect 49868 44380 49924 44382
rect 50204 45164 50260 45220
rect 49756 44268 49812 44324
rect 49756 43820 49812 43876
rect 50876 49420 50932 49476
rect 51772 49644 51828 49700
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 53788 50540 53844 50596
rect 53900 50428 53956 50484
rect 53340 49868 53396 49924
rect 52556 49644 52612 49700
rect 51884 49532 51940 49588
rect 53676 49138 53732 49140
rect 53676 49086 53678 49138
rect 53678 49086 53730 49138
rect 53730 49086 53732 49138
rect 53676 49084 53732 49086
rect 51884 49026 51940 49028
rect 51884 48974 51886 49026
rect 51886 48974 51938 49026
rect 51938 48974 51940 49026
rect 51884 48972 51940 48974
rect 52780 49026 52836 49028
rect 52780 48974 52782 49026
rect 52782 48974 52834 49026
rect 52834 48974 52836 49026
rect 52780 48972 52836 48974
rect 53004 48972 53060 49028
rect 52220 48748 52276 48804
rect 52444 47852 52500 47908
rect 50876 46732 50932 46788
rect 50428 45612 50484 45668
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 52220 46508 52276 46564
rect 51548 45218 51604 45220
rect 51548 45166 51550 45218
rect 51550 45166 51602 45218
rect 51602 45166 51604 45218
rect 51548 45164 51604 45166
rect 51100 44434 51156 44436
rect 51100 44382 51102 44434
rect 51102 44382 51154 44434
rect 51154 44382 51156 44434
rect 51100 44380 51156 44382
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50316 43708 50372 43764
rect 49532 43650 49588 43652
rect 49532 43598 49534 43650
rect 49534 43598 49586 43650
rect 49586 43598 49588 43650
rect 49532 43596 49588 43598
rect 49980 43596 50036 43652
rect 50876 43596 50932 43652
rect 50988 43538 51044 43540
rect 50988 43486 50990 43538
rect 50990 43486 51042 43538
rect 51042 43486 51044 43538
rect 50988 43484 51044 43486
rect 51548 43596 51604 43652
rect 51436 43484 51492 43540
rect 50204 43426 50260 43428
rect 50204 43374 50206 43426
rect 50206 43374 50258 43426
rect 50258 43374 50260 43426
rect 50204 43372 50260 43374
rect 51548 43372 51604 43428
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 51772 43650 51828 43652
rect 51772 43598 51774 43650
rect 51774 43598 51826 43650
rect 51826 43598 51828 43650
rect 51772 43596 51828 43598
rect 52332 46450 52388 46452
rect 52332 46398 52334 46450
rect 52334 46398 52386 46450
rect 52386 46398 52388 46450
rect 52332 46396 52388 46398
rect 52892 47516 52948 47572
rect 52332 45724 52388 45780
rect 52668 45612 52724 45668
rect 52668 44940 52724 44996
rect 52332 44828 52388 44884
rect 51436 41244 51492 41300
rect 52108 41298 52164 41300
rect 52108 41246 52110 41298
rect 52110 41246 52162 41298
rect 52162 41246 52164 41298
rect 52108 41244 52164 41246
rect 51100 40962 51156 40964
rect 51100 40910 51102 40962
rect 51102 40910 51154 40962
rect 51154 40910 51156 40962
rect 51100 40908 51156 40910
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50316 40124 50372 40180
rect 51436 40124 51492 40180
rect 50204 40012 50260 40068
rect 48412 39900 48468 39956
rect 49196 39730 49252 39732
rect 49196 39678 49198 39730
rect 49198 39678 49250 39730
rect 49250 39678 49252 39730
rect 49196 39676 49252 39678
rect 47404 38668 47460 38724
rect 47292 37378 47348 37380
rect 47292 37326 47294 37378
rect 47294 37326 47346 37378
rect 47346 37326 47348 37378
rect 47292 37324 47348 37326
rect 46732 37154 46788 37156
rect 46732 37102 46734 37154
rect 46734 37102 46786 37154
rect 46786 37102 46788 37154
rect 46732 37100 46788 37102
rect 45836 35980 45892 36036
rect 46396 36540 46452 36596
rect 41804 34748 41860 34804
rect 42924 34802 42980 34804
rect 42924 34750 42926 34802
rect 42926 34750 42978 34802
rect 42978 34750 42980 34802
rect 42924 34748 42980 34750
rect 43596 34748 43652 34804
rect 41132 34076 41188 34132
rect 40460 33906 40516 33908
rect 40460 33854 40462 33906
rect 40462 33854 40514 33906
rect 40514 33854 40516 33906
rect 40460 33852 40516 33854
rect 39900 33404 39956 33460
rect 40348 33292 40404 33348
rect 39340 32956 39396 33012
rect 39900 33068 39956 33124
rect 41468 34130 41524 34132
rect 41468 34078 41470 34130
rect 41470 34078 41522 34130
rect 41522 34078 41524 34130
rect 41468 34076 41524 34078
rect 41916 33516 41972 33572
rect 41244 33292 41300 33348
rect 38668 32284 38724 32340
rect 40460 31948 40516 32004
rect 37324 31666 37380 31668
rect 37324 31614 37326 31666
rect 37326 31614 37378 31666
rect 37378 31614 37380 31666
rect 37324 31612 37380 31614
rect 37324 31276 37380 31332
rect 36092 31218 36148 31220
rect 36092 31166 36094 31218
rect 36094 31166 36146 31218
rect 36146 31166 36148 31218
rect 36092 31164 36148 31166
rect 37772 31276 37828 31332
rect 36652 30770 36708 30772
rect 36652 30718 36654 30770
rect 36654 30718 36706 30770
rect 36706 30718 36708 30770
rect 36652 30716 36708 30718
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35644 30268 35700 30324
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 27804 35140 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 36204 29426 36260 29428
rect 36204 29374 36206 29426
rect 36206 29374 36258 29426
rect 36258 29374 36260 29426
rect 36204 29372 36260 29374
rect 36316 28700 36372 28756
rect 35756 27804 35812 27860
rect 37100 29260 37156 29316
rect 38220 30156 38276 30212
rect 38332 31612 38388 31668
rect 38332 30940 38388 30996
rect 41132 31612 41188 31668
rect 39900 31218 39956 31220
rect 39900 31166 39902 31218
rect 39902 31166 39954 31218
rect 39954 31166 39956 31218
rect 39900 31164 39956 31166
rect 39788 30994 39844 30996
rect 39788 30942 39790 30994
rect 39790 30942 39842 30994
rect 39842 30942 39844 30994
rect 39788 30940 39844 30942
rect 42924 33458 42980 33460
rect 42924 33406 42926 33458
rect 42926 33406 42978 33458
rect 42978 33406 42980 33458
rect 42924 33404 42980 33406
rect 43260 33458 43316 33460
rect 43260 33406 43262 33458
rect 43262 33406 43314 33458
rect 43314 33406 43316 33458
rect 43260 33404 43316 33406
rect 42924 32844 42980 32900
rect 41916 31666 41972 31668
rect 41916 31614 41918 31666
rect 41918 31614 41970 31666
rect 41970 31614 41972 31666
rect 41916 31612 41972 31614
rect 41692 31500 41748 31556
rect 43372 31554 43428 31556
rect 43372 31502 43374 31554
rect 43374 31502 43426 31554
rect 43426 31502 43428 31554
rect 43372 31500 43428 31502
rect 41468 30994 41524 30996
rect 41468 30942 41470 30994
rect 41470 30942 41522 30994
rect 41522 30942 41524 30994
rect 41468 30940 41524 30942
rect 38668 30828 38724 30884
rect 40684 30210 40740 30212
rect 40684 30158 40686 30210
rect 40686 30158 40738 30210
rect 40738 30158 40740 30210
rect 40684 30156 40740 30158
rect 40012 29986 40068 29988
rect 40012 29934 40014 29986
rect 40014 29934 40066 29986
rect 40066 29934 40068 29986
rect 40012 29932 40068 29934
rect 38444 29372 38500 29428
rect 38892 29372 38948 29428
rect 38332 28700 38388 28756
rect 37660 28418 37716 28420
rect 37660 28366 37662 28418
rect 37662 28366 37714 28418
rect 37714 28366 37716 28418
rect 37660 28364 37716 28366
rect 37548 28140 37604 28196
rect 38556 29314 38612 29316
rect 38556 29262 38558 29314
rect 38558 29262 38610 29314
rect 38610 29262 38612 29314
rect 38556 29260 38612 29262
rect 37100 27074 37156 27076
rect 37100 27022 37102 27074
rect 37102 27022 37154 27074
rect 37154 27022 37156 27074
rect 37100 27020 37156 27022
rect 36092 26962 36148 26964
rect 36092 26910 36094 26962
rect 36094 26910 36146 26962
rect 36146 26910 36148 26962
rect 36092 26908 36148 26910
rect 34748 26460 34804 26516
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34076 23660 34132 23716
rect 33740 23324 33796 23380
rect 33964 22988 34020 23044
rect 34300 23884 34356 23940
rect 34300 22316 34356 22372
rect 34412 23548 34468 23604
rect 34076 21474 34132 21476
rect 34076 21422 34078 21474
rect 34078 21422 34130 21474
rect 34130 21422 34132 21474
rect 34076 21420 34132 21422
rect 33740 20412 33796 20468
rect 34636 21868 34692 21924
rect 34524 21756 34580 21812
rect 34636 18508 34692 18564
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35084 23938 35140 23940
rect 35084 23886 35086 23938
rect 35086 23886 35138 23938
rect 35138 23886 35140 23938
rect 35084 23884 35140 23886
rect 34860 21756 34916 21812
rect 34972 22316 35028 22372
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35756 22988 35812 23044
rect 35532 22092 35588 22148
rect 35756 21868 35812 21924
rect 35196 21698 35252 21700
rect 35196 21646 35198 21698
rect 35198 21646 35250 21698
rect 35250 21646 35252 21698
rect 35196 21644 35252 21646
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36876 26684 36932 26740
rect 36428 25452 36484 25508
rect 36428 23884 36484 23940
rect 36092 23548 36148 23604
rect 37100 23938 37156 23940
rect 37100 23886 37102 23938
rect 37102 23886 37154 23938
rect 37154 23886 37156 23938
rect 37100 23884 37156 23886
rect 37100 23548 37156 23604
rect 35868 21644 35924 21700
rect 35308 16994 35364 16996
rect 35308 16942 35310 16994
rect 35310 16942 35362 16994
rect 35362 16942 35364 16994
rect 35308 16940 35364 16942
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35756 21362 35812 21364
rect 35756 21310 35758 21362
rect 35758 21310 35810 21362
rect 35810 21310 35812 21362
rect 35756 21308 35812 21310
rect 36540 21868 36596 21924
rect 35980 20860 36036 20916
rect 36652 20188 36708 20244
rect 35756 18508 35812 18564
rect 36988 20914 37044 20916
rect 36988 20862 36990 20914
rect 36990 20862 37042 20914
rect 37042 20862 37044 20914
rect 36988 20860 37044 20862
rect 37324 25228 37380 25284
rect 37436 24220 37492 24276
rect 37324 22876 37380 22932
rect 38108 23100 38164 23156
rect 37660 22988 37716 23044
rect 38220 21868 38276 21924
rect 37996 20636 38052 20692
rect 37996 20188 38052 20244
rect 38556 27020 38612 27076
rect 38780 28140 38836 28196
rect 38444 25788 38500 25844
rect 38444 25506 38500 25508
rect 38444 25454 38446 25506
rect 38446 25454 38498 25506
rect 38498 25454 38500 25506
rect 38444 25452 38500 25454
rect 38444 23154 38500 23156
rect 38444 23102 38446 23154
rect 38446 23102 38498 23154
rect 38498 23102 38500 23154
rect 38444 23100 38500 23102
rect 38444 21756 38500 21812
rect 40572 28812 40628 28868
rect 40908 29932 40964 29988
rect 40684 29372 40740 29428
rect 39900 28364 39956 28420
rect 39676 27804 39732 27860
rect 40236 27970 40292 27972
rect 40236 27918 40238 27970
rect 40238 27918 40290 27970
rect 40290 27918 40292 27970
rect 40236 27916 40292 27918
rect 40012 27692 40068 27748
rect 40684 27074 40740 27076
rect 40684 27022 40686 27074
rect 40686 27022 40738 27074
rect 40738 27022 40740 27074
rect 40684 27020 40740 27022
rect 39004 25228 39060 25284
rect 39564 25564 39620 25620
rect 39900 25788 39956 25844
rect 39116 24556 39172 24612
rect 39004 23660 39060 23716
rect 38892 23154 38948 23156
rect 38892 23102 38894 23154
rect 38894 23102 38946 23154
rect 38946 23102 38948 23154
rect 38892 23100 38948 23102
rect 38892 20636 38948 20692
rect 39564 23154 39620 23156
rect 39564 23102 39566 23154
rect 39566 23102 39618 23154
rect 39618 23102 39620 23154
rect 39564 23100 39620 23102
rect 39788 23042 39844 23044
rect 39788 22990 39790 23042
rect 39790 22990 39842 23042
rect 39842 22990 39844 23042
rect 39788 22988 39844 22990
rect 39452 21586 39508 21588
rect 39452 21534 39454 21586
rect 39454 21534 39506 21586
rect 39506 21534 39508 21586
rect 39452 21532 39508 21534
rect 39788 21586 39844 21588
rect 39788 21534 39790 21586
rect 39790 21534 39842 21586
rect 39842 21534 39844 21586
rect 39788 21532 39844 21534
rect 40348 24610 40404 24612
rect 40348 24558 40350 24610
rect 40350 24558 40402 24610
rect 40402 24558 40404 24610
rect 40348 24556 40404 24558
rect 40124 24220 40180 24276
rect 40012 20300 40068 20356
rect 40348 23772 40404 23828
rect 40684 24332 40740 24388
rect 40908 25004 40964 25060
rect 44492 34018 44548 34020
rect 44492 33966 44494 34018
rect 44494 33966 44546 34018
rect 44546 33966 44548 34018
rect 44492 33964 44548 33966
rect 43932 33740 43988 33796
rect 43932 33458 43988 33460
rect 43932 33406 43934 33458
rect 43934 33406 43986 33458
rect 43986 33406 43988 33458
rect 43932 33404 43988 33406
rect 45052 33740 45108 33796
rect 43820 33122 43876 33124
rect 43820 33070 43822 33122
rect 43822 33070 43874 33122
rect 43874 33070 43876 33122
rect 43820 33068 43876 33070
rect 43708 32844 43764 32900
rect 44940 32786 44996 32788
rect 44940 32734 44942 32786
rect 44942 32734 44994 32786
rect 44994 32734 44996 32786
rect 44940 32732 44996 32734
rect 44716 32396 44772 32452
rect 43708 31500 43764 31556
rect 43596 30156 43652 30212
rect 41692 29708 41748 29764
rect 41580 29596 41636 29652
rect 41916 29596 41972 29652
rect 42252 29426 42308 29428
rect 42252 29374 42254 29426
rect 42254 29374 42306 29426
rect 42306 29374 42308 29426
rect 42252 29372 42308 29374
rect 41916 27916 41972 27972
rect 41468 27692 41524 27748
rect 41356 27074 41412 27076
rect 41356 27022 41358 27074
rect 41358 27022 41410 27074
rect 41410 27022 41412 27074
rect 41356 27020 41412 27022
rect 41132 24892 41188 24948
rect 40796 23772 40852 23828
rect 40460 23548 40516 23604
rect 40572 22540 40628 22596
rect 41020 23772 41076 23828
rect 41020 21532 41076 21588
rect 41020 20188 41076 20244
rect 41132 24332 41188 24388
rect 40796 19068 40852 19124
rect 41356 22764 41412 22820
rect 41244 18956 41300 19012
rect 41916 25564 41972 25620
rect 41580 25340 41636 25396
rect 42364 25394 42420 25396
rect 42364 25342 42366 25394
rect 42366 25342 42418 25394
rect 42418 25342 42420 25394
rect 42364 25340 42420 25342
rect 42140 24892 42196 24948
rect 41692 24556 41748 24612
rect 41580 23660 41636 23716
rect 41356 18396 41412 18452
rect 41804 20300 41860 20356
rect 42364 24556 42420 24612
rect 42252 21532 42308 21588
rect 42700 25618 42756 25620
rect 42700 25566 42702 25618
rect 42702 25566 42754 25618
rect 42754 25566 42756 25618
rect 42700 25564 42756 25566
rect 43932 29708 43988 29764
rect 45388 33346 45444 33348
rect 45388 33294 45390 33346
rect 45390 33294 45442 33346
rect 45442 33294 45444 33346
rect 45388 33292 45444 33294
rect 45388 32562 45444 32564
rect 45388 32510 45390 32562
rect 45390 32510 45442 32562
rect 45442 32510 45444 32562
rect 45388 32508 45444 32510
rect 45388 32172 45444 32228
rect 46060 33740 46116 33796
rect 46284 33180 46340 33236
rect 47068 36482 47124 36484
rect 47068 36430 47070 36482
rect 47070 36430 47122 36482
rect 47122 36430 47124 36482
rect 47068 36428 47124 36430
rect 47852 37436 47908 37492
rect 48972 38722 49028 38724
rect 48972 38670 48974 38722
rect 48974 38670 49026 38722
rect 49026 38670 49028 38722
rect 48972 38668 49028 38670
rect 47964 37324 48020 37380
rect 48412 37826 48468 37828
rect 48412 37774 48414 37826
rect 48414 37774 48466 37826
rect 48466 37774 48468 37826
rect 48412 37772 48468 37774
rect 48524 37324 48580 37380
rect 49196 38332 49252 38388
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 49644 38444 49700 38500
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 48860 37324 48916 37380
rect 48188 37100 48244 37156
rect 48412 36988 48468 37044
rect 48076 36482 48132 36484
rect 48076 36430 48078 36482
rect 48078 36430 48130 36482
rect 48130 36430 48132 36482
rect 48076 36428 48132 36430
rect 48972 37436 49028 37492
rect 49532 37378 49588 37380
rect 49532 37326 49534 37378
rect 49534 37326 49586 37378
rect 49586 37326 49588 37378
rect 49532 37324 49588 37326
rect 50652 37100 50708 37156
rect 47628 35532 47684 35588
rect 52444 39676 52500 39732
rect 53452 48188 53508 48244
rect 53564 48130 53620 48132
rect 53564 48078 53566 48130
rect 53566 48078 53618 48130
rect 53618 48078 53620 48130
rect 53564 48076 53620 48078
rect 53228 47964 53284 48020
rect 54124 49922 54180 49924
rect 54124 49870 54126 49922
rect 54126 49870 54178 49922
rect 54178 49870 54180 49922
rect 54124 49868 54180 49870
rect 54348 49532 54404 49588
rect 55020 49532 55076 49588
rect 54684 48914 54740 48916
rect 54684 48862 54686 48914
rect 54686 48862 54738 48914
rect 54738 48862 54740 48914
rect 54684 48860 54740 48862
rect 54012 47964 54068 48020
rect 53228 46786 53284 46788
rect 53228 46734 53230 46786
rect 53230 46734 53282 46786
rect 53282 46734 53284 46786
rect 53228 46732 53284 46734
rect 56252 49868 56308 49924
rect 55356 49532 55412 49588
rect 55468 48188 55524 48244
rect 55692 48300 55748 48356
rect 55132 47852 55188 47908
rect 56476 49420 56532 49476
rect 57820 50482 57876 50484
rect 57820 50430 57822 50482
rect 57822 50430 57874 50482
rect 57874 50430 57876 50482
rect 57820 50428 57876 50430
rect 58828 49922 58884 49924
rect 58828 49870 58830 49922
rect 58830 49870 58882 49922
rect 58882 49870 58884 49922
rect 58828 49868 58884 49870
rect 56812 48972 56868 49028
rect 57484 48914 57540 48916
rect 57484 48862 57486 48914
rect 57486 48862 57538 48914
rect 57538 48862 57540 48914
rect 57484 48860 57540 48862
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 57596 48300 57652 48356
rect 57596 47740 57652 47796
rect 57484 47570 57540 47572
rect 57484 47518 57486 47570
rect 57486 47518 57538 47570
rect 57538 47518 57540 47570
rect 57484 47516 57540 47518
rect 56140 47292 56196 47348
rect 54572 46172 54628 46228
rect 55692 45836 55748 45892
rect 53116 45276 53172 45332
rect 58492 47346 58548 47348
rect 58492 47294 58494 47346
rect 58494 47294 58546 47346
rect 58546 47294 58548 47346
rect 58492 47292 58548 47294
rect 56252 47068 56308 47124
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 58828 47068 58884 47124
rect 58828 46786 58884 46788
rect 58828 46734 58830 46786
rect 58830 46734 58882 46786
rect 58882 46734 58884 46786
rect 58828 46732 58884 46734
rect 59388 46786 59444 46788
rect 59388 46734 59390 46786
rect 59390 46734 59442 46786
rect 59442 46734 59444 46786
rect 59388 46732 59444 46734
rect 57484 46002 57540 46004
rect 57484 45950 57486 46002
rect 57486 45950 57538 46002
rect 57538 45950 57540 46002
rect 57484 45948 57540 45950
rect 52780 43708 52836 43764
rect 52780 43484 52836 43540
rect 53004 44380 53060 44436
rect 55356 45218 55412 45220
rect 55356 45166 55358 45218
rect 55358 45166 55410 45218
rect 55410 45166 55412 45218
rect 55356 45164 55412 45166
rect 56700 44994 56756 44996
rect 56700 44942 56702 44994
rect 56702 44942 56754 44994
rect 56754 44942 56756 44994
rect 56700 44940 56756 44942
rect 59276 45890 59332 45892
rect 59276 45838 59278 45890
rect 59278 45838 59330 45890
rect 59330 45838 59332 45890
rect 59276 45836 59332 45838
rect 58492 45778 58548 45780
rect 58492 45726 58494 45778
rect 58494 45726 58546 45778
rect 58546 45726 58548 45778
rect 58492 45724 58548 45726
rect 57596 45276 57652 45332
rect 61404 46396 61460 46452
rect 59500 45612 59556 45668
rect 54124 44716 54180 44772
rect 55468 44156 55524 44212
rect 54908 43650 54964 43652
rect 54908 43598 54910 43650
rect 54910 43598 54962 43650
rect 54962 43598 54964 43650
rect 54908 43596 54964 43598
rect 54684 43538 54740 43540
rect 54684 43486 54686 43538
rect 54686 43486 54738 43538
rect 54738 43486 54740 43538
rect 54684 43484 54740 43486
rect 55132 43372 55188 43428
rect 53228 43260 53284 43316
rect 56028 43708 56084 43764
rect 56140 43596 56196 43652
rect 55356 42194 55412 42196
rect 55356 42142 55358 42194
rect 55358 42142 55410 42194
rect 55410 42142 55412 42194
rect 55356 42140 55412 42142
rect 55580 41244 55636 41300
rect 53116 40402 53172 40404
rect 53116 40350 53118 40402
rect 53118 40350 53170 40402
rect 53170 40350 53172 40402
rect 53116 40348 53172 40350
rect 53676 40124 53732 40180
rect 53004 39676 53060 39732
rect 53788 39676 53844 39732
rect 53228 38946 53284 38948
rect 53228 38894 53230 38946
rect 53230 38894 53282 38946
rect 53282 38894 53284 38946
rect 53228 38892 53284 38894
rect 53788 38780 53844 38836
rect 52780 38050 52836 38052
rect 52780 37998 52782 38050
rect 52782 37998 52834 38050
rect 52834 37998 52836 38050
rect 52780 37996 52836 37998
rect 53340 38108 53396 38164
rect 50876 36652 50932 36708
rect 52220 37826 52276 37828
rect 52220 37774 52222 37826
rect 52222 37774 52274 37826
rect 52274 37774 52276 37826
rect 52220 37772 52276 37774
rect 53116 37324 53172 37380
rect 53228 36540 53284 36596
rect 50428 36428 50484 36484
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50428 35196 50484 35252
rect 50988 35196 51044 35252
rect 50652 34690 50708 34692
rect 50652 34638 50654 34690
rect 50654 34638 50706 34690
rect 50706 34638 50708 34690
rect 50652 34636 50708 34638
rect 50556 34522 50612 34524
rect 48748 34412 48804 34468
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 47068 33852 47124 33908
rect 47964 33740 48020 33796
rect 47068 33516 47124 33572
rect 47628 33234 47684 33236
rect 47628 33182 47630 33234
rect 47630 33182 47682 33234
rect 47682 33182 47684 33234
rect 47628 33180 47684 33182
rect 46396 32732 46452 32788
rect 47180 32956 47236 33012
rect 48412 32732 48468 32788
rect 45612 32508 45668 32564
rect 44492 30770 44548 30772
rect 44492 30718 44494 30770
rect 44494 30718 44546 30770
rect 44546 30718 44548 30770
rect 44492 30716 44548 30718
rect 44156 29596 44212 29652
rect 44156 29372 44212 29428
rect 43148 25564 43204 25620
rect 42924 23996 42980 24052
rect 43148 25004 43204 25060
rect 42700 23548 42756 23604
rect 42588 21420 42644 21476
rect 42364 20188 42420 20244
rect 42924 22540 42980 22596
rect 42364 19292 42420 19348
rect 42588 19122 42644 19124
rect 42588 19070 42590 19122
rect 42590 19070 42642 19122
rect 42642 19070 42644 19122
rect 42588 19068 42644 19070
rect 42588 18396 42644 18452
rect 42812 18060 42868 18116
rect 44380 28364 44436 28420
rect 45164 30604 45220 30660
rect 44716 29596 44772 29652
rect 48076 32562 48132 32564
rect 48076 32510 48078 32562
rect 48078 32510 48130 32562
rect 48130 32510 48132 32562
rect 48076 32508 48132 32510
rect 45724 32450 45780 32452
rect 45724 32398 45726 32450
rect 45726 32398 45778 32450
rect 45778 32398 45780 32450
rect 45724 32396 45780 32398
rect 46172 32284 46228 32340
rect 47068 32284 47124 32340
rect 47068 31724 47124 31780
rect 47852 31554 47908 31556
rect 47852 31502 47854 31554
rect 47854 31502 47906 31554
rect 47906 31502 47908 31554
rect 47852 31500 47908 31502
rect 45612 31276 45668 31332
rect 45388 29484 45444 29540
rect 46060 30716 46116 30772
rect 45948 29202 46004 29204
rect 45948 29150 45950 29202
rect 45950 29150 46002 29202
rect 46002 29150 46004 29202
rect 45948 29148 46004 29150
rect 45612 28812 45668 28868
rect 45500 28642 45556 28644
rect 45500 28590 45502 28642
rect 45502 28590 45554 28642
rect 45554 28590 45556 28642
rect 45500 28588 45556 28590
rect 43932 27244 43988 27300
rect 44156 27020 44212 27076
rect 44044 26012 44100 26068
rect 44044 25618 44100 25620
rect 44044 25566 44046 25618
rect 44046 25566 44098 25618
rect 44098 25566 44100 25618
rect 44044 25564 44100 25566
rect 43708 24108 43764 24164
rect 43932 22204 43988 22260
rect 43708 19628 43764 19684
rect 44828 27858 44884 27860
rect 44828 27806 44830 27858
rect 44830 27806 44882 27858
rect 44882 27806 44884 27858
rect 44828 27804 44884 27806
rect 45388 27074 45444 27076
rect 45388 27022 45390 27074
rect 45390 27022 45442 27074
rect 45442 27022 45444 27074
rect 45388 27020 45444 27022
rect 44492 26514 44548 26516
rect 44492 26462 44494 26514
rect 44494 26462 44546 26514
rect 44546 26462 44548 26514
rect 44492 26460 44548 26462
rect 45052 26796 45108 26852
rect 45500 26124 45556 26180
rect 45388 25676 45444 25732
rect 45612 25228 45668 25284
rect 44380 23436 44436 23492
rect 44828 22652 44884 22708
rect 45276 24220 45332 24276
rect 44268 19628 44324 19684
rect 44380 19346 44436 19348
rect 44380 19294 44382 19346
rect 44382 19294 44434 19346
rect 44434 19294 44436 19346
rect 44380 19292 44436 19294
rect 44492 19068 44548 19124
rect 44940 22092 44996 22148
rect 45836 22652 45892 22708
rect 45388 21980 45444 22036
rect 45612 21868 45668 21924
rect 45052 20130 45108 20132
rect 45052 20078 45054 20130
rect 45054 20078 45106 20130
rect 45106 20078 45108 20130
rect 45052 20076 45108 20078
rect 44716 19964 44772 20020
rect 45388 19852 45444 19908
rect 45052 19346 45108 19348
rect 45052 19294 45054 19346
rect 45054 19294 45106 19346
rect 45106 19294 45108 19346
rect 45052 19292 45108 19294
rect 45724 21532 45780 21588
rect 44604 18620 44660 18676
rect 46284 30210 46340 30212
rect 46284 30158 46286 30210
rect 46286 30158 46338 30210
rect 46338 30158 46340 30210
rect 46284 30156 46340 30158
rect 46732 30156 46788 30212
rect 46284 29650 46340 29652
rect 46284 29598 46286 29650
rect 46286 29598 46338 29650
rect 46338 29598 46340 29650
rect 46284 29596 46340 29598
rect 49308 34300 49364 34356
rect 48860 34130 48916 34132
rect 48860 34078 48862 34130
rect 48862 34078 48914 34130
rect 48914 34078 48916 34130
rect 48860 34076 48916 34078
rect 49196 33346 49252 33348
rect 49196 33294 49198 33346
rect 49198 33294 49250 33346
rect 49250 33294 49252 33346
rect 49196 33292 49252 33294
rect 48748 33180 48804 33236
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 52556 36482 52612 36484
rect 52556 36430 52558 36482
rect 52558 36430 52610 36482
rect 52610 36430 52612 36482
rect 52556 36428 52612 36430
rect 51324 35196 51380 35252
rect 52108 35196 52164 35252
rect 53900 37378 53956 37380
rect 53900 37326 53902 37378
rect 53902 37326 53954 37378
rect 53954 37326 53956 37378
rect 53900 37324 53956 37326
rect 54236 37266 54292 37268
rect 54236 37214 54238 37266
rect 54238 37214 54290 37266
rect 54290 37214 54292 37266
rect 54236 37212 54292 37214
rect 53676 36316 53732 36372
rect 53676 35922 53732 35924
rect 53676 35870 53678 35922
rect 53678 35870 53730 35922
rect 53730 35870 53732 35922
rect 53676 35868 53732 35870
rect 54684 37324 54740 37380
rect 55468 40460 55524 40516
rect 58828 44828 58884 44884
rect 58940 45164 58996 45220
rect 60620 45666 60676 45668
rect 60620 45614 60622 45666
rect 60622 45614 60674 45666
rect 60674 45614 60676 45666
rect 60620 45612 60676 45614
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 57596 44268 57652 44324
rect 58268 44210 58324 44212
rect 58268 44158 58270 44210
rect 58270 44158 58322 44210
rect 58322 44158 58324 44210
rect 58268 44156 58324 44158
rect 57596 44044 57652 44100
rect 56700 43484 56756 43540
rect 56252 42642 56308 42644
rect 56252 42590 56254 42642
rect 56254 42590 56306 42642
rect 56306 42590 56308 42642
rect 56252 42588 56308 42590
rect 56252 42028 56308 42084
rect 56700 41970 56756 41972
rect 56700 41918 56702 41970
rect 56702 41918 56754 41970
rect 56754 41918 56756 41970
rect 56700 41916 56756 41918
rect 56812 43708 56868 43764
rect 57148 43426 57204 43428
rect 57148 43374 57150 43426
rect 57150 43374 57202 43426
rect 57202 43374 57204 43426
rect 57148 43372 57204 43374
rect 58492 43708 58548 43764
rect 60396 44994 60452 44996
rect 60396 44942 60398 44994
rect 60398 44942 60450 44994
rect 60450 44942 60452 44994
rect 60396 44940 60452 44942
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 61516 44434 61572 44436
rect 61516 44382 61518 44434
rect 61518 44382 61570 44434
rect 61570 44382 61572 44434
rect 61516 44380 61572 44382
rect 60060 44156 60116 44212
rect 59500 43762 59556 43764
rect 59500 43710 59502 43762
rect 59502 43710 59554 43762
rect 59554 43710 59556 43762
rect 59500 43708 59556 43710
rect 59276 43372 59332 43428
rect 58828 43148 58884 43204
rect 57036 42812 57092 42868
rect 58828 42364 58884 42420
rect 59276 42140 59332 42196
rect 56812 41244 56868 41300
rect 56140 40684 56196 40740
rect 57596 41858 57652 41860
rect 57596 41806 57598 41858
rect 57598 41806 57650 41858
rect 57650 41806 57652 41858
rect 57596 41804 57652 41806
rect 55580 37324 55636 37380
rect 56700 39394 56756 39396
rect 56700 39342 56702 39394
rect 56702 39342 56754 39394
rect 56754 39342 56756 39394
rect 56700 39340 56756 39342
rect 59500 41970 59556 41972
rect 59500 41918 59502 41970
rect 59502 41918 59554 41970
rect 59554 41918 59556 41970
rect 59500 41916 59556 41918
rect 59388 41804 59444 41860
rect 62524 44210 62580 44212
rect 62524 44158 62526 44210
rect 62526 44158 62578 44210
rect 62578 44158 62580 44210
rect 62524 44156 62580 44158
rect 61404 43650 61460 43652
rect 61404 43598 61406 43650
rect 61406 43598 61458 43650
rect 61458 43598 61460 43650
rect 61404 43596 61460 43598
rect 60396 43426 60452 43428
rect 60396 43374 60398 43426
rect 60398 43374 60450 43426
rect 60450 43374 60452 43426
rect 60396 43372 60452 43374
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 61516 42866 61572 42868
rect 61516 42814 61518 42866
rect 61518 42814 61570 42866
rect 61570 42814 61572 42866
rect 61516 42812 61572 42814
rect 62524 42642 62580 42644
rect 62524 42590 62526 42642
rect 62526 42590 62578 42642
rect 62578 42590 62580 42642
rect 62524 42588 62580 42590
rect 61404 42082 61460 42084
rect 61404 42030 61406 42082
rect 61406 42030 61458 42082
rect 61458 42030 61460 42082
rect 61404 42028 61460 42030
rect 59612 41692 59668 41748
rect 58492 41074 58548 41076
rect 58492 41022 58494 41074
rect 58494 41022 58546 41074
rect 58546 41022 58548 41074
rect 58492 41020 58548 41022
rect 62188 41858 62244 41860
rect 62188 41806 62190 41858
rect 62190 41806 62242 41858
rect 62242 41806 62244 41858
rect 62188 41804 62244 41806
rect 62412 41692 62468 41748
rect 62972 41692 63028 41748
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 60396 41132 60452 41188
rect 61404 40908 61460 40964
rect 58828 40514 58884 40516
rect 58828 40462 58830 40514
rect 58830 40462 58882 40514
rect 58882 40462 58884 40514
rect 58828 40460 58884 40462
rect 61516 40348 61572 40404
rect 60396 40012 60452 40068
rect 57596 39788 57652 39844
rect 58940 39900 58996 39956
rect 57932 39730 57988 39732
rect 57932 39678 57934 39730
rect 57934 39678 57986 39730
rect 57986 39678 57988 39730
rect 57932 39676 57988 39678
rect 57484 39004 57540 39060
rect 57596 39564 57652 39620
rect 56700 38780 56756 38836
rect 62524 40684 62580 40740
rect 61740 40124 61796 40180
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 61404 39340 61460 39396
rect 57596 38220 57652 38276
rect 56700 37378 56756 37380
rect 56700 37326 56702 37378
rect 56702 37326 56754 37378
rect 56754 37326 56756 37378
rect 56700 37324 56756 37326
rect 55468 37212 55524 37268
rect 54348 35644 54404 35700
rect 54460 35868 54516 35924
rect 51436 33740 51492 33796
rect 51212 32732 51268 32788
rect 48524 32396 48580 32452
rect 48300 31836 48356 31892
rect 48076 30268 48132 30324
rect 47740 30044 47796 30100
rect 46844 29596 46900 29652
rect 47740 28700 47796 28756
rect 47852 27692 47908 27748
rect 48188 28924 48244 28980
rect 49756 32450 49812 32452
rect 49756 32398 49758 32450
rect 49758 32398 49810 32450
rect 49810 32398 49812 32450
rect 49756 32396 49812 32398
rect 50764 32284 50820 32340
rect 53676 34412 53732 34468
rect 52332 34354 52388 34356
rect 52332 34302 52334 34354
rect 52334 34302 52386 34354
rect 52386 34302 52388 34354
rect 52332 34300 52388 34302
rect 52444 34130 52500 34132
rect 52444 34078 52446 34130
rect 52446 34078 52498 34130
rect 52498 34078 52500 34130
rect 52444 34076 52500 34078
rect 53116 33628 53172 33684
rect 52220 33122 52276 33124
rect 52220 33070 52222 33122
rect 52222 33070 52274 33122
rect 52274 33070 52276 33122
rect 52220 33068 52276 33070
rect 49308 30994 49364 30996
rect 49308 30942 49310 30994
rect 49310 30942 49362 30994
rect 49362 30942 49364 30994
rect 49308 30940 49364 30942
rect 48748 30268 48804 30324
rect 48524 28866 48580 28868
rect 48524 28814 48526 28866
rect 48526 28814 48578 28866
rect 48578 28814 48580 28866
rect 48524 28812 48580 28814
rect 48412 27916 48468 27972
rect 46956 26012 47012 26068
rect 47628 25228 47684 25284
rect 47740 24946 47796 24948
rect 47740 24894 47742 24946
rect 47742 24894 47794 24946
rect 47794 24894 47796 24946
rect 47740 24892 47796 24894
rect 46060 23772 46116 23828
rect 46508 24108 46564 24164
rect 46060 23436 46116 23492
rect 46060 23100 46116 23156
rect 46060 21868 46116 21924
rect 45948 21532 46004 21588
rect 46060 21420 46116 21476
rect 45836 18956 45892 19012
rect 44716 18060 44772 18116
rect 45948 17500 46004 17556
rect 46284 22204 46340 22260
rect 46956 23100 47012 23156
rect 46732 20130 46788 20132
rect 46732 20078 46734 20130
rect 46734 20078 46786 20130
rect 46786 20078 46788 20130
rect 46732 20076 46788 20078
rect 47068 20130 47124 20132
rect 47068 20078 47070 20130
rect 47070 20078 47122 20130
rect 47122 20078 47124 20130
rect 47068 20076 47124 20078
rect 46396 19628 46452 19684
rect 47068 19122 47124 19124
rect 47068 19070 47070 19122
rect 47070 19070 47122 19122
rect 47122 19070 47124 19122
rect 47068 19068 47124 19070
rect 46844 18562 46900 18564
rect 46844 18510 46846 18562
rect 46846 18510 46898 18562
rect 46898 18510 46900 18562
rect 46844 18508 46900 18510
rect 47068 18396 47124 18452
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50876 30492 50932 30548
rect 51548 31554 51604 31556
rect 51548 31502 51550 31554
rect 51550 31502 51602 31554
rect 51602 31502 51604 31554
rect 51548 31500 51604 31502
rect 50428 30098 50484 30100
rect 50428 30046 50430 30098
rect 50430 30046 50482 30098
rect 50482 30046 50484 30098
rect 50428 30044 50484 30046
rect 49644 29932 49700 29988
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 49308 29426 49364 29428
rect 49308 29374 49310 29426
rect 49310 29374 49362 29426
rect 49362 29374 49364 29426
rect 49308 29372 49364 29374
rect 49756 28924 49812 28980
rect 49644 28028 49700 28084
rect 48748 27804 48804 27860
rect 49196 27746 49252 27748
rect 49196 27694 49198 27746
rect 49198 27694 49250 27746
rect 49250 27694 49252 27746
rect 49196 27692 49252 27694
rect 49532 27746 49588 27748
rect 49532 27694 49534 27746
rect 49534 27694 49586 27746
rect 49586 27694 49588 27746
rect 49532 27692 49588 27694
rect 49084 27020 49140 27076
rect 49084 26460 49140 26516
rect 48412 25564 48468 25620
rect 48748 26012 48804 26068
rect 48972 25506 49028 25508
rect 48972 25454 48974 25506
rect 48974 25454 49026 25506
rect 49026 25454 49028 25506
rect 48972 25452 49028 25454
rect 49196 25676 49252 25732
rect 49308 25340 49364 25396
rect 49196 24780 49252 24836
rect 47964 23548 48020 23604
rect 47516 20076 47572 20132
rect 47852 18562 47908 18564
rect 47852 18510 47854 18562
rect 47854 18510 47906 18562
rect 47906 18510 47908 18562
rect 47852 18508 47908 18510
rect 48300 22540 48356 22596
rect 48412 22258 48468 22260
rect 48412 22206 48414 22258
rect 48414 22206 48466 22258
rect 48466 22206 48468 22258
rect 48412 22204 48468 22206
rect 48860 24668 48916 24724
rect 49420 24610 49476 24612
rect 49420 24558 49422 24610
rect 49422 24558 49474 24610
rect 49474 24558 49476 24610
rect 49420 24556 49476 24558
rect 51100 28924 51156 28980
rect 49980 28588 50036 28644
rect 49980 27858 50036 27860
rect 49980 27806 49982 27858
rect 49982 27806 50034 27858
rect 50034 27806 50036 27858
rect 49980 27804 50036 27806
rect 50316 28364 50372 28420
rect 49756 27692 49812 27748
rect 48860 23324 48916 23380
rect 48860 23154 48916 23156
rect 48860 23102 48862 23154
rect 48862 23102 48914 23154
rect 48914 23102 48916 23154
rect 48860 23100 48916 23102
rect 48524 21756 48580 21812
rect 48412 21026 48468 21028
rect 48412 20974 48414 21026
rect 48414 20974 48466 21026
rect 48466 20974 48468 21026
rect 48412 20972 48468 20974
rect 48188 20130 48244 20132
rect 48188 20078 48190 20130
rect 48190 20078 48242 20130
rect 48242 20078 48244 20130
rect 48188 20076 48244 20078
rect 48860 22092 48916 22148
rect 48636 20188 48692 20244
rect 49308 23154 49364 23156
rect 49308 23102 49310 23154
rect 49310 23102 49362 23154
rect 49362 23102 49364 23154
rect 49308 23100 49364 23102
rect 51100 28364 51156 28420
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 51212 28028 51268 28084
rect 50652 27356 50708 27412
rect 53900 32844 53956 32900
rect 54236 32844 54292 32900
rect 53900 32508 53956 32564
rect 54908 35420 54964 35476
rect 62524 38892 62580 38948
rect 60396 38332 60452 38388
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 61516 38162 61572 38164
rect 61516 38110 61518 38162
rect 61518 38110 61570 38162
rect 61570 38110 61572 38162
rect 61516 38108 61572 38110
rect 58828 37996 58884 38052
rect 61404 37772 61460 37828
rect 60396 37154 60452 37156
rect 60396 37102 60398 37154
rect 60398 37102 60450 37154
rect 60450 37102 60452 37154
rect 60396 37100 60452 37102
rect 58828 36988 58884 37044
rect 57596 36876 57652 36932
rect 56252 36764 56308 36820
rect 56588 36482 56644 36484
rect 56588 36430 56590 36482
rect 56590 36430 56642 36482
rect 56642 36430 56644 36482
rect 56588 36428 56644 36430
rect 55580 35420 55636 35476
rect 54572 35196 54628 35252
rect 55356 34636 55412 34692
rect 56364 35138 56420 35140
rect 56364 35086 56366 35138
rect 56366 35086 56418 35138
rect 56418 35086 56420 35138
rect 56364 35084 56420 35086
rect 58492 36652 58548 36708
rect 57596 35026 57652 35028
rect 57596 34974 57598 35026
rect 57598 34974 57650 35026
rect 57650 34974 57652 35026
rect 57596 34972 57652 34974
rect 56140 34748 56196 34804
rect 54684 33404 54740 33460
rect 56476 32956 56532 33012
rect 53788 31948 53844 32004
rect 52556 30828 52612 30884
rect 53228 31836 53284 31892
rect 52332 30770 52388 30772
rect 52332 30718 52334 30770
rect 52334 30718 52386 30770
rect 52386 30718 52388 30770
rect 52332 30716 52388 30718
rect 52220 30156 52276 30212
rect 52668 30268 52724 30324
rect 51996 30098 52052 30100
rect 51996 30046 51998 30098
rect 51998 30046 52050 30098
rect 52050 30046 52052 30098
rect 51996 30044 52052 30046
rect 51660 28754 51716 28756
rect 51660 28702 51662 28754
rect 51662 28702 51714 28754
rect 51714 28702 51716 28754
rect 51660 28700 51716 28702
rect 52332 29202 52388 29204
rect 52332 29150 52334 29202
rect 52334 29150 52386 29202
rect 52386 29150 52388 29202
rect 52332 29148 52388 29150
rect 51996 28754 52052 28756
rect 51996 28702 51998 28754
rect 51998 28702 52050 28754
rect 52050 28702 52052 28754
rect 51996 28700 52052 28702
rect 51996 28364 52052 28420
rect 52444 28364 52500 28420
rect 52780 30098 52836 30100
rect 52780 30046 52782 30098
rect 52782 30046 52834 30098
rect 52834 30046 52836 30098
rect 52780 30044 52836 30046
rect 53228 29820 53284 29876
rect 53900 30210 53956 30212
rect 53900 30158 53902 30210
rect 53902 30158 53954 30210
rect 53954 30158 53956 30210
rect 53900 30156 53956 30158
rect 52668 28642 52724 28644
rect 52668 28590 52670 28642
rect 52670 28590 52722 28642
rect 52722 28590 52724 28642
rect 52668 28588 52724 28590
rect 50764 27074 50820 27076
rect 50764 27022 50766 27074
rect 50766 27022 50818 27074
rect 50818 27022 50820 27074
rect 50764 27020 50820 27022
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50316 26348 50372 26404
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50204 24946 50260 24948
rect 50204 24894 50206 24946
rect 50206 24894 50258 24946
rect 50258 24894 50260 24946
rect 50204 24892 50260 24894
rect 50876 24834 50932 24836
rect 50876 24782 50878 24834
rect 50878 24782 50930 24834
rect 50930 24782 50932 24834
rect 50876 24780 50932 24782
rect 51212 24722 51268 24724
rect 51212 24670 51214 24722
rect 51214 24670 51266 24722
rect 51266 24670 51268 24722
rect 51212 24668 51268 24670
rect 50092 24050 50148 24052
rect 50092 23998 50094 24050
rect 50094 23998 50146 24050
rect 50146 23998 50148 24050
rect 50092 23996 50148 23998
rect 51100 23826 51156 23828
rect 51100 23774 51102 23826
rect 51102 23774 51154 23826
rect 51154 23774 51156 23826
rect 51100 23772 51156 23774
rect 49756 23548 49812 23604
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 49644 23324 49700 23380
rect 49084 22370 49140 22372
rect 49084 22318 49086 22370
rect 49086 22318 49138 22370
rect 49138 22318 49140 22370
rect 49084 22316 49140 22318
rect 49644 22092 49700 22148
rect 50204 23100 50260 23156
rect 49644 21644 49700 21700
rect 49532 21196 49588 21252
rect 49756 21532 49812 21588
rect 48860 20130 48916 20132
rect 48860 20078 48862 20130
rect 48862 20078 48914 20130
rect 48914 20078 48916 20130
rect 48860 20076 48916 20078
rect 48636 19964 48692 20020
rect 49644 19740 49700 19796
rect 50428 22540 50484 22596
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50764 20130 50820 20132
rect 50764 20078 50766 20130
rect 50766 20078 50818 20130
rect 50818 20078 50820 20130
rect 50764 20076 50820 20078
rect 53004 28028 53060 28084
rect 52332 26066 52388 26068
rect 52332 26014 52334 26066
rect 52334 26014 52386 26066
rect 52386 26014 52388 26066
rect 52332 26012 52388 26014
rect 51772 25116 51828 25172
rect 53116 27916 53172 27972
rect 53228 27692 53284 27748
rect 53564 27244 53620 27300
rect 53228 27074 53284 27076
rect 53228 27022 53230 27074
rect 53230 27022 53282 27074
rect 53282 27022 53284 27074
rect 53228 27020 53284 27022
rect 53676 26460 53732 26516
rect 51996 24780 52052 24836
rect 51772 23772 51828 23828
rect 52444 24668 52500 24724
rect 53452 24892 53508 24948
rect 52892 24668 52948 24724
rect 53116 23884 53172 23940
rect 51884 22988 51940 23044
rect 52332 22930 52388 22932
rect 52332 22878 52334 22930
rect 52334 22878 52386 22930
rect 52386 22878 52388 22930
rect 52332 22876 52388 22878
rect 51884 22092 51940 22148
rect 51436 19964 51492 20020
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 54348 28700 54404 28756
rect 54348 28028 54404 28084
rect 55468 30322 55524 30324
rect 55468 30270 55470 30322
rect 55470 30270 55522 30322
rect 55522 30270 55524 30322
rect 55468 30268 55524 30270
rect 55580 30044 55636 30100
rect 54908 27970 54964 27972
rect 54908 27918 54910 27970
rect 54910 27918 54962 27970
rect 54962 27918 54964 27970
rect 54908 27916 54964 27918
rect 55244 27970 55300 27972
rect 55244 27918 55246 27970
rect 55246 27918 55298 27970
rect 55298 27918 55300 27970
rect 55244 27916 55300 27918
rect 56252 31554 56308 31556
rect 56252 31502 56254 31554
rect 56254 31502 56306 31554
rect 56306 31502 56308 31554
rect 56252 31500 56308 31502
rect 57596 34018 57652 34020
rect 57596 33966 57598 34018
rect 57598 33966 57650 34018
rect 57650 33966 57652 34018
rect 57596 33964 57652 33966
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 62524 36652 62580 36708
rect 61516 36594 61572 36596
rect 61516 36542 61518 36594
rect 61518 36542 61570 36594
rect 61570 36542 61572 36594
rect 61516 36540 61572 36542
rect 62524 36370 62580 36372
rect 62524 36318 62526 36370
rect 62526 36318 62578 36370
rect 62578 36318 62580 36370
rect 62524 36316 62580 36318
rect 58828 35810 58884 35812
rect 58828 35758 58830 35810
rect 58830 35758 58882 35810
rect 58882 35758 58884 35810
rect 58828 35756 58884 35758
rect 60396 35586 60452 35588
rect 60396 35534 60398 35586
rect 60398 35534 60450 35586
rect 60450 35534 60452 35586
rect 60396 35532 60452 35534
rect 59388 35420 59444 35476
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 61404 35084 61460 35140
rect 58828 34802 58884 34804
rect 58828 34750 58830 34802
rect 58830 34750 58882 34802
rect 58882 34750 58884 34802
rect 58828 34748 58884 34750
rect 59500 34690 59556 34692
rect 59500 34638 59502 34690
rect 59502 34638 59554 34690
rect 59554 34638 59556 34690
rect 59500 34636 59556 34638
rect 62524 34802 62580 34804
rect 62524 34750 62526 34802
rect 62526 34750 62578 34802
rect 62578 34750 62580 34802
rect 62524 34748 62580 34750
rect 61516 34412 61572 34468
rect 61404 34300 61460 34356
rect 58828 34242 58884 34244
rect 58828 34190 58830 34242
rect 58830 34190 58882 34242
rect 58882 34190 58884 34242
rect 58828 34188 58884 34190
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 61516 33516 61572 33572
rect 60396 33292 60452 33348
rect 62524 33234 62580 33236
rect 62524 33182 62526 33234
rect 62526 33182 62578 33234
rect 62578 33182 62580 33234
rect 62524 33180 62580 33182
rect 61404 33068 61460 33124
rect 60396 32732 60452 32788
rect 58828 32674 58884 32676
rect 58828 32622 58830 32674
rect 58830 32622 58882 32674
rect 58882 32622 58884 32674
rect 58828 32620 58884 32622
rect 57708 32508 57764 32564
rect 57596 32450 57652 32452
rect 57596 32398 57598 32450
rect 57598 32398 57650 32450
rect 57650 32398 57652 32450
rect 57596 32396 57652 32398
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 57036 31724 57092 31780
rect 56140 31276 56196 31332
rect 57036 31164 57092 31220
rect 57148 31388 57204 31444
rect 61516 31890 61572 31892
rect 61516 31838 61518 31890
rect 61518 31838 61570 31890
rect 61570 31838 61572 31890
rect 61516 31836 61572 31838
rect 58492 31666 58548 31668
rect 58492 31614 58494 31666
rect 58494 31614 58546 31666
rect 58546 31614 58548 31666
rect 58492 31612 58548 31614
rect 65548 31500 65604 31556
rect 64316 31388 64372 31444
rect 62524 31276 62580 31332
rect 57484 31052 57540 31108
rect 55916 30268 55972 30324
rect 57484 30604 57540 30660
rect 56476 30268 56532 30324
rect 56028 28588 56084 28644
rect 56028 27970 56084 27972
rect 56028 27918 56030 27970
rect 56030 27918 56082 27970
rect 56082 27918 56084 27970
rect 56028 27916 56084 27918
rect 56252 27916 56308 27972
rect 55580 27580 55636 27636
rect 57596 29484 57652 29540
rect 58828 29036 58884 29092
rect 60508 31218 60564 31220
rect 60508 31166 60510 31218
rect 60510 31166 60562 31218
rect 60562 31166 60564 31218
rect 60508 31164 60564 31166
rect 60172 30994 60228 30996
rect 60172 30942 60174 30994
rect 60174 30942 60226 30994
rect 60226 30942 60228 30994
rect 60172 30940 60228 30942
rect 61516 30828 61572 30884
rect 64988 30994 65044 30996
rect 64988 30942 64990 30994
rect 64990 30942 65042 30994
rect 65042 30942 65044 30994
rect 64988 30940 65044 30942
rect 66108 30994 66164 30996
rect 66108 30942 66110 30994
rect 66110 30942 66162 30994
rect 66162 30942 66164 30994
rect 66108 30940 66164 30942
rect 62412 30716 62468 30772
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 61404 30044 61460 30100
rect 61516 29820 61572 29876
rect 60396 29314 60452 29316
rect 60396 29262 60398 29314
rect 60398 29262 60450 29314
rect 60450 29262 60452 29314
rect 60396 29260 60452 29262
rect 61404 28812 61460 28868
rect 62524 28924 62580 28980
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 59276 28642 59332 28644
rect 59276 28590 59278 28642
rect 59278 28590 59330 28642
rect 59330 28590 59332 28642
rect 59276 28588 59332 28590
rect 57596 28476 57652 28532
rect 62524 28530 62580 28532
rect 62524 28478 62526 28530
rect 62526 28478 62578 28530
rect 62578 28478 62580 28530
rect 62524 28476 62580 28478
rect 58492 27804 58548 27860
rect 57484 27186 57540 27188
rect 57484 27134 57486 27186
rect 57486 27134 57538 27186
rect 57538 27134 57540 27186
rect 57484 27132 57540 27134
rect 58492 26796 58548 26852
rect 56364 26684 56420 26740
rect 54572 26402 54628 26404
rect 54572 26350 54574 26402
rect 54574 26350 54626 26402
rect 54626 26350 54628 26402
rect 54572 26348 54628 26350
rect 58828 26402 58884 26404
rect 58828 26350 58830 26402
rect 58830 26350 58882 26402
rect 58882 26350 58884 26402
rect 58828 26348 58884 26350
rect 55132 25116 55188 25172
rect 53900 23884 53956 23940
rect 53676 22652 53732 22708
rect 52892 21644 52948 21700
rect 53228 21420 53284 21476
rect 57596 26178 57652 26180
rect 57596 26126 57598 26178
rect 57598 26126 57650 26178
rect 57650 26126 57652 26178
rect 57596 26124 57652 26126
rect 57596 25340 57652 25396
rect 55916 25282 55972 25284
rect 55916 25230 55918 25282
rect 55918 25230 55970 25282
rect 55970 25230 55972 25282
rect 55916 25228 55972 25230
rect 56476 24780 56532 24836
rect 54908 24498 54964 24500
rect 54908 24446 54910 24498
rect 54910 24446 54962 24498
rect 54962 24446 54964 24498
rect 54908 24444 54964 24446
rect 58716 25564 58772 25620
rect 61404 27970 61460 27972
rect 61404 27918 61406 27970
rect 61406 27918 61458 27970
rect 61458 27918 61460 27970
rect 61404 27916 61460 27918
rect 60396 27746 60452 27748
rect 60396 27694 60398 27746
rect 60398 27694 60450 27746
rect 60450 27694 60452 27746
rect 60396 27692 60452 27694
rect 59276 27580 59332 27636
rect 65916 27466 65972 27468
rect 60284 27356 60340 27412
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 58940 25452 58996 25508
rect 61516 27020 61572 27076
rect 61404 26684 61460 26740
rect 62524 26012 62580 26068
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 58828 24834 58884 24836
rect 58828 24782 58830 24834
rect 58830 24782 58882 24834
rect 58882 24782 58884 24834
rect 58828 24780 58884 24782
rect 57708 24220 57764 24276
rect 55468 23996 55524 24052
rect 55916 23996 55972 24052
rect 54348 22540 54404 22596
rect 53900 22204 53956 22260
rect 52220 20636 52276 20692
rect 53676 21196 53732 21252
rect 52556 19906 52612 19908
rect 52556 19854 52558 19906
rect 52558 19854 52610 19906
rect 52610 19854 52612 19906
rect 52556 19852 52612 19854
rect 54012 21644 54068 21700
rect 54796 20972 54852 21028
rect 54684 20690 54740 20692
rect 54684 20638 54686 20690
rect 54686 20638 54738 20690
rect 54738 20638 54740 20690
rect 54684 20636 54740 20638
rect 55580 22540 55636 22596
rect 55692 22204 55748 22260
rect 58604 24050 58660 24052
rect 58604 23998 58606 24050
rect 58606 23998 58658 24050
rect 58658 23998 58660 24050
rect 58604 23996 58660 23998
rect 59612 25282 59668 25284
rect 59612 25230 59614 25282
rect 59614 25230 59666 25282
rect 59666 25230 59668 25282
rect 59612 25228 59668 25230
rect 60396 24892 60452 24948
rect 61404 24444 61460 24500
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 59500 23996 59556 24052
rect 56476 23938 56532 23940
rect 56476 23886 56478 23938
rect 56478 23886 56530 23938
rect 56530 23886 56532 23938
rect 56476 23884 56532 23886
rect 58268 23826 58324 23828
rect 58268 23774 58270 23826
rect 58270 23774 58322 23826
rect 58322 23774 58324 23826
rect 58268 23772 58324 23774
rect 56252 23212 56308 23268
rect 58828 23266 58884 23268
rect 58828 23214 58830 23266
rect 58830 23214 58882 23266
rect 58882 23214 58884 23266
rect 58828 23212 58884 23214
rect 57596 23042 57652 23044
rect 57596 22990 57598 23042
rect 57598 22990 57650 23042
rect 57650 22990 57652 23042
rect 57596 22988 57652 22990
rect 58492 22876 58548 22932
rect 57484 22482 57540 22484
rect 57484 22430 57486 22482
rect 57486 22430 57538 22482
rect 57538 22430 57540 22482
rect 57484 22428 57540 22430
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 59612 22204 59668 22260
rect 56140 21644 56196 21700
rect 58828 21698 58884 21700
rect 58828 21646 58830 21698
rect 58830 21646 58882 21698
rect 58882 21646 58884 21698
rect 58828 21644 58884 21646
rect 57596 21474 57652 21476
rect 57596 21422 57598 21474
rect 57598 21422 57650 21474
rect 57650 21422 57652 21474
rect 57596 21420 57652 21422
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 55916 20076 55972 20132
rect 54460 20018 54516 20020
rect 54460 19966 54462 20018
rect 54462 19966 54514 20018
rect 54514 19966 54516 20018
rect 54460 19964 54516 19966
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 52668 19068 52724 19124
rect 55020 19122 55076 19124
rect 55020 19070 55022 19122
rect 55022 19070 55074 19122
rect 55074 19070 55076 19122
rect 55020 19068 55076 19070
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 49644 17554 49700 17556
rect 49644 17502 49646 17554
rect 49646 17502 49698 17554
rect 49698 17502 49700 17554
rect 49644 17500 49700 17502
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 41692 15932 41748 15988
rect 43708 15986 43764 15988
rect 43708 15934 43710 15986
rect 43710 15934 43762 15986
rect 43762 15934 43764 15986
rect 43708 15932 43764 15934
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 67200 62580 68000 62608
rect 66210 62524 66220 62580
rect 66276 62524 68000 62580
rect 67200 62496 68000 62524
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 41458 54348 41468 54404
rect 41524 54348 42700 54404
rect 42756 54348 42766 54404
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 28578 53788 28588 53844
rect 28644 53788 30380 53844
rect 30436 53788 30446 53844
rect 43026 53788 43036 53844
rect 43092 53788 45836 53844
rect 45892 53788 45902 53844
rect 37314 53564 37324 53620
rect 37380 53564 39564 53620
rect 39620 53564 39630 53620
rect 44482 53564 44492 53620
rect 44548 53564 47068 53620
rect 47124 53564 47134 53620
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 36642 53004 36652 53060
rect 36708 53004 38668 53060
rect 38724 53004 38734 53060
rect 44594 53004 44604 53060
rect 44660 53004 45948 53060
rect 46004 53004 46014 53060
rect 36418 52780 36428 52836
rect 36484 52780 37660 52836
rect 37716 52780 37726 52836
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 33394 52220 33404 52276
rect 33460 52220 34412 52276
rect 34468 52220 34478 52276
rect 35746 52220 35756 52276
rect 35812 52220 37996 52276
rect 38052 52220 38062 52276
rect 39442 52220 39452 52276
rect 39508 52220 42364 52276
rect 42420 52220 42430 52276
rect 41682 52108 41692 52164
rect 41748 52108 43708 52164
rect 43764 52108 43774 52164
rect 48636 52108 51100 52164
rect 51156 52108 51166 52164
rect 48636 52052 48692 52108
rect 32946 51996 32956 52052
rect 33012 51996 35420 52052
rect 35476 51996 35486 52052
rect 40674 51996 40684 52052
rect 40740 51996 41804 52052
rect 41860 51996 41870 52052
rect 48626 51996 48636 52052
rect 48692 51996 48702 52052
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 27906 51436 27916 51492
rect 27972 51436 29036 51492
rect 29092 51436 29102 51492
rect 34962 51436 34972 51492
rect 35028 51436 37772 51492
rect 37828 51436 37838 51492
rect 45938 51436 45948 51492
rect 46004 51436 50764 51492
rect 50820 51436 50830 51492
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 35186 50764 35196 50820
rect 35252 50764 35868 50820
rect 35924 50764 35934 50820
rect 38994 50652 39004 50708
rect 39060 50652 45836 50708
rect 45892 50652 45902 50708
rect 46050 50652 46060 50708
rect 46116 50652 48636 50708
rect 48692 50652 48702 50708
rect 38210 50540 38220 50596
rect 38276 50540 40796 50596
rect 40852 50540 40862 50596
rect 48636 50540 53788 50596
rect 53844 50540 53854 50596
rect 48636 50484 48692 50540
rect 40450 50428 40460 50484
rect 40516 50428 47068 50484
rect 47124 50428 47134 50484
rect 48626 50428 48636 50484
rect 48692 50428 48702 50484
rect 53890 50428 53900 50484
rect 53956 50428 57820 50484
rect 57876 50428 57886 50484
rect 42466 50316 42476 50372
rect 42532 50316 44940 50372
rect 44996 50316 45006 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 41346 50092 41356 50148
rect 41412 50092 45724 50148
rect 45780 50092 45790 50148
rect 29698 49868 29708 49924
rect 29764 49868 31052 49924
rect 31108 49868 31118 49924
rect 33170 49868 33180 49924
rect 33236 49868 35308 49924
rect 35364 49868 35374 49924
rect 36306 49868 36316 49924
rect 36372 49868 36988 49924
rect 37044 49868 37054 49924
rect 45378 49868 45388 49924
rect 45444 49868 46844 49924
rect 46900 49868 46910 49924
rect 53330 49868 53340 49924
rect 53396 49868 54124 49924
rect 54180 49868 54190 49924
rect 56242 49868 56252 49924
rect 56308 49868 58828 49924
rect 58884 49868 58894 49924
rect 25666 49756 25676 49812
rect 25732 49756 27244 49812
rect 27300 49756 27310 49812
rect 45602 49756 45612 49812
rect 45668 49756 48412 49812
rect 48468 49756 48478 49812
rect 25442 49644 25452 49700
rect 25508 49644 26124 49700
rect 26180 49644 27916 49700
rect 27972 49644 28140 49700
rect 28196 49644 28206 49700
rect 44818 49644 44828 49700
rect 44884 49644 46172 49700
rect 46228 49644 46238 49700
rect 46386 49644 46396 49700
rect 46452 49644 47068 49700
rect 47124 49644 47516 49700
rect 47572 49644 47582 49700
rect 47954 49644 47964 49700
rect 48020 49644 49420 49700
rect 49476 49644 49980 49700
rect 50036 49644 51604 49700
rect 51762 49644 51772 49700
rect 51828 49644 52556 49700
rect 52612 49644 52622 49700
rect 51548 49588 51604 49644
rect 36530 49532 36540 49588
rect 36596 49532 39116 49588
rect 39172 49532 39182 49588
rect 45378 49532 45388 49588
rect 45444 49532 49868 49588
rect 49924 49532 49934 49588
rect 51548 49532 51884 49588
rect 51940 49532 54348 49588
rect 54404 49532 55020 49588
rect 55076 49532 55356 49588
rect 55412 49532 55422 49588
rect 50866 49420 50876 49476
rect 50932 49420 56476 49476
rect 56532 49420 56542 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 29922 49196 29932 49252
rect 29988 49196 31388 49252
rect 31444 49196 31454 49252
rect 41570 49196 41580 49252
rect 41636 49196 44716 49252
rect 44772 49196 44782 49252
rect 45602 49084 45612 49140
rect 45668 49084 53676 49140
rect 53732 49084 53742 49140
rect 32050 48972 32060 49028
rect 32116 48972 33404 49028
rect 33460 48972 33470 49028
rect 39106 48972 39116 49028
rect 39172 48972 41916 49028
rect 41972 48972 41982 49028
rect 51874 48972 51884 49028
rect 51940 48972 52780 49028
rect 52836 48972 52846 49028
rect 52994 48972 53004 49028
rect 53060 48972 56812 49028
rect 56868 48972 56878 49028
rect 26562 48860 26572 48916
rect 26628 48860 28028 48916
rect 28084 48860 28094 48916
rect 28690 48860 28700 48916
rect 28756 48860 30716 48916
rect 30772 48860 30782 48916
rect 32722 48860 32732 48916
rect 32788 48860 34636 48916
rect 34692 48860 34702 48916
rect 41346 48860 41356 48916
rect 41412 48860 42252 48916
rect 42308 48860 42924 48916
rect 42980 48860 43484 48916
rect 43540 48860 46396 48916
rect 46452 48860 46462 48916
rect 48402 48860 48412 48916
rect 48468 48860 54684 48916
rect 54740 48860 54750 48916
rect 55412 48860 57484 48916
rect 57540 48860 57550 48916
rect 55412 48804 55468 48860
rect 27346 48748 27356 48804
rect 27412 48748 28252 48804
rect 28308 48748 28318 48804
rect 28466 48748 28476 48804
rect 28532 48748 28812 48804
rect 28868 48748 28878 48804
rect 29586 48748 29596 48804
rect 29652 48748 30268 48804
rect 30324 48748 30334 48804
rect 33506 48748 33516 48804
rect 33572 48748 34860 48804
rect 34916 48748 34926 48804
rect 41122 48748 41132 48804
rect 41188 48748 42812 48804
rect 42868 48748 42878 48804
rect 46498 48748 46508 48804
rect 46564 48748 49868 48804
rect 49924 48748 49934 48804
rect 52210 48748 52220 48804
rect 52276 48748 55468 48804
rect 47730 48636 47740 48692
rect 47796 48636 49756 48692
rect 49812 48636 49822 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 20290 48524 20300 48580
rect 20356 48524 22316 48580
rect 22372 48524 22382 48580
rect 24210 48524 24220 48580
rect 24276 48524 25228 48580
rect 25284 48524 25294 48580
rect 31154 48300 31164 48356
rect 31220 48300 32620 48356
rect 32676 48300 32686 48356
rect 55682 48300 55692 48356
rect 55748 48300 57596 48356
rect 57652 48300 57662 48356
rect 30258 48188 30268 48244
rect 30324 48188 30828 48244
rect 30884 48188 31948 48244
rect 32004 48188 32284 48244
rect 32340 48188 35420 48244
rect 35476 48188 36092 48244
rect 36148 48188 36158 48244
rect 36754 48188 36764 48244
rect 36820 48188 37996 48244
rect 38052 48188 38062 48244
rect 44258 48188 44268 48244
rect 44324 48188 44828 48244
rect 44884 48188 45612 48244
rect 45668 48188 45678 48244
rect 53442 48188 53452 48244
rect 53508 48188 55468 48244
rect 55524 48188 55534 48244
rect 19730 48076 19740 48132
rect 19796 48076 21308 48132
rect 21364 48076 21374 48132
rect 23874 48076 23884 48132
rect 23940 48076 25676 48132
rect 25732 48076 25742 48132
rect 32610 48076 32620 48132
rect 32676 48076 33068 48132
rect 33124 48076 33134 48132
rect 38882 48076 38892 48132
rect 38948 48076 40908 48132
rect 40964 48076 40974 48132
rect 49522 48076 49532 48132
rect 49588 48076 53564 48132
rect 53620 48076 53630 48132
rect 25330 47964 25340 48020
rect 25396 47964 25900 48020
rect 25956 47964 25966 48020
rect 42466 47964 42476 48020
rect 42532 47964 43148 48020
rect 43204 47964 43214 48020
rect 53218 47964 53228 48020
rect 53284 47964 54012 48020
rect 54068 47964 54078 48020
rect 52434 47852 52444 47908
rect 52500 47852 55132 47908
rect 55188 47852 55198 47908
rect 0 47796 800 47824
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 0 47740 4228 47796
rect 0 47712 800 47740
rect 4172 47684 4228 47740
rect 55412 47740 57596 47796
rect 57652 47740 57662 47796
rect 4172 47628 10892 47684
rect 10948 47628 10958 47684
rect 55412 47572 55468 47740
rect 24322 47516 24332 47572
rect 24388 47516 25116 47572
rect 25172 47516 25182 47572
rect 38612 47516 40460 47572
rect 40516 47516 40796 47572
rect 40852 47516 41916 47572
rect 41972 47516 41982 47572
rect 52882 47516 52892 47572
rect 52948 47516 55468 47572
rect 57474 47516 57484 47572
rect 57540 47516 57550 47572
rect 38612 47460 38668 47516
rect 57484 47460 57540 47516
rect 22428 47404 25340 47460
rect 25396 47404 25406 47460
rect 31714 47404 31724 47460
rect 31780 47404 32844 47460
rect 32900 47404 35980 47460
rect 36036 47404 36764 47460
rect 36820 47404 38668 47460
rect 49410 47404 49420 47460
rect 49476 47404 57540 47460
rect 22428 47348 22484 47404
rect 21634 47292 21644 47348
rect 21700 47292 22428 47348
rect 22484 47292 22494 47348
rect 24658 47292 24668 47348
rect 24724 47292 27132 47348
rect 27188 47292 27198 47348
rect 56130 47292 56140 47348
rect 56196 47292 58492 47348
rect 58548 47292 58558 47348
rect 17154 47180 17164 47236
rect 17220 47180 18508 47236
rect 18564 47180 18574 47236
rect 27906 47180 27916 47236
rect 27972 47180 30156 47236
rect 30212 47180 30222 47236
rect 38210 47180 38220 47236
rect 38276 47180 42028 47236
rect 42084 47180 42094 47236
rect 42242 47180 42252 47236
rect 42308 47180 42924 47236
rect 42980 47180 42990 47236
rect 44370 47180 44380 47236
rect 44436 47180 49308 47236
rect 49364 47180 49374 47236
rect 22866 47068 22876 47124
rect 22932 47068 23772 47124
rect 23828 47068 23838 47124
rect 44930 47068 44940 47124
rect 44996 47068 46284 47124
rect 46340 47068 48076 47124
rect 48132 47068 48524 47124
rect 48580 47068 48590 47124
rect 56242 47068 56252 47124
rect 56308 47068 58828 47124
rect 58884 47068 58894 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 20850 46956 20860 47012
rect 20916 46956 21756 47012
rect 21812 46956 21822 47012
rect 23650 46956 23660 47012
rect 23716 46956 25564 47012
rect 25620 46956 25630 47012
rect 28130 46844 28140 46900
rect 28196 46844 29484 46900
rect 29540 46844 29550 46900
rect 46834 46844 46844 46900
rect 46900 46844 47628 46900
rect 47684 46844 47694 46900
rect 55412 46844 59444 46900
rect 55412 46788 55468 46844
rect 59388 46788 59444 46844
rect 40338 46732 40348 46788
rect 40404 46732 41244 46788
rect 41300 46732 41310 46788
rect 44706 46732 44716 46788
rect 44772 46732 50876 46788
rect 50932 46732 50942 46788
rect 53218 46732 53228 46788
rect 53284 46732 55468 46788
rect 58818 46732 58828 46788
rect 58884 46732 58894 46788
rect 59378 46732 59388 46788
rect 59444 46732 59454 46788
rect 25106 46620 25116 46676
rect 25172 46620 26460 46676
rect 26516 46620 28140 46676
rect 28196 46620 29036 46676
rect 29092 46620 29102 46676
rect 58828 46564 58884 46732
rect 17826 46508 17836 46564
rect 17892 46508 18844 46564
rect 18900 46508 18910 46564
rect 52210 46508 52220 46564
rect 52276 46508 58884 46564
rect 19618 46396 19628 46452
rect 19684 46396 24444 46452
rect 24500 46396 24510 46452
rect 52322 46396 52332 46452
rect 52388 46396 61404 46452
rect 61460 46396 61470 46452
rect 23762 46284 23772 46340
rect 23828 46284 28364 46340
rect 28420 46284 28430 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 21970 46172 21980 46228
rect 22036 46172 23660 46228
rect 23716 46172 23726 46228
rect 49634 46172 49644 46228
rect 49700 46172 54572 46228
rect 54628 46172 54638 46228
rect 19506 46060 19516 46116
rect 19572 46060 21308 46116
rect 21364 46060 21374 46116
rect 22642 46060 22652 46116
rect 22708 46060 29036 46116
rect 29092 46060 29102 46116
rect 41010 45948 41020 46004
rect 41076 45948 41804 46004
rect 41860 45948 44828 46004
rect 44884 45948 44894 46004
rect 49298 45948 49308 46004
rect 49364 45948 57484 46004
rect 57540 45948 57550 46004
rect 20850 45836 20860 45892
rect 20916 45836 21420 45892
rect 21476 45836 25116 45892
rect 25172 45836 25182 45892
rect 55682 45836 55692 45892
rect 55748 45836 59276 45892
rect 59332 45836 59342 45892
rect 29810 45724 29820 45780
rect 29876 45724 31724 45780
rect 31780 45724 31790 45780
rect 52322 45724 52332 45780
rect 52388 45724 58492 45780
rect 58548 45724 58558 45780
rect 17154 45612 17164 45668
rect 17220 45612 18620 45668
rect 18676 45612 18686 45668
rect 20290 45612 20300 45668
rect 20356 45612 22540 45668
rect 22596 45612 22606 45668
rect 23538 45612 23548 45668
rect 23604 45612 24332 45668
rect 24388 45612 24398 45668
rect 32050 45612 32060 45668
rect 32116 45612 33964 45668
rect 34020 45612 34030 45668
rect 42914 45612 42924 45668
rect 42980 45612 45724 45668
rect 45780 45612 50428 45668
rect 50484 45612 52668 45668
rect 52724 45612 52734 45668
rect 59490 45612 59500 45668
rect 59556 45612 60620 45668
rect 60676 45612 60686 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 40236 45388 46172 45444
rect 46228 45388 46238 45444
rect 40236 45332 40292 45388
rect 32498 45276 32508 45332
rect 32564 45276 33740 45332
rect 33796 45276 33806 45332
rect 38612 45276 40292 45332
rect 45378 45276 45388 45332
rect 45444 45276 47292 45332
rect 47348 45276 47358 45332
rect 48178 45276 48188 45332
rect 48244 45276 49868 45332
rect 49924 45276 49934 45332
rect 53106 45276 53116 45332
rect 53172 45276 57596 45332
rect 57652 45276 57662 45332
rect 25666 45164 25676 45220
rect 25732 45164 27356 45220
rect 27412 45164 27422 45220
rect 38612 45108 38668 45276
rect 39890 45164 39900 45220
rect 39956 45164 41468 45220
rect 41524 45164 41534 45220
rect 43138 45164 43148 45220
rect 43204 45164 45164 45220
rect 45220 45164 45230 45220
rect 50194 45164 50204 45220
rect 50260 45164 51548 45220
rect 51604 45164 51614 45220
rect 55346 45164 55356 45220
rect 55412 45164 58940 45220
rect 58996 45164 59006 45220
rect 26674 45052 26684 45108
rect 26740 45052 29148 45108
rect 29204 45052 30940 45108
rect 30996 45052 31006 45108
rect 37426 45052 37436 45108
rect 37492 45052 38668 45108
rect 19506 44940 19516 44996
rect 19572 44940 24892 44996
rect 24948 44940 24958 44996
rect 41458 44940 41468 44996
rect 41524 44940 42700 44996
rect 42756 44940 42766 44996
rect 43586 44940 43596 44996
rect 43652 44940 46508 44996
rect 46564 44940 47180 44996
rect 47236 44940 47246 44996
rect 52658 44940 52668 44996
rect 52724 44940 56700 44996
rect 56756 44940 56766 44996
rect 60386 44940 60396 44996
rect 60452 44940 60462 44996
rect 16930 44828 16940 44884
rect 16996 44828 17500 44884
rect 17556 44828 21644 44884
rect 21700 44828 23660 44884
rect 23716 44828 24108 44884
rect 24164 44828 24174 44884
rect 29362 44828 29372 44884
rect 29428 44828 32620 44884
rect 32676 44828 32686 44884
rect 52322 44828 52332 44884
rect 52388 44828 58828 44884
rect 58884 44828 58894 44884
rect 60396 44772 60452 44940
rect 54114 44716 54124 44772
rect 54180 44716 60452 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 29810 44380 29820 44436
rect 29876 44380 32284 44436
rect 32340 44380 33740 44436
rect 33796 44380 33806 44436
rect 49858 44380 49868 44436
rect 49924 44380 51100 44436
rect 51156 44380 51166 44436
rect 52994 44380 53004 44436
rect 53060 44380 61516 44436
rect 61572 44380 61582 44436
rect 31490 44268 31500 44324
rect 31556 44268 32844 44324
rect 32900 44268 36428 44324
rect 36484 44268 36988 44324
rect 37044 44268 37054 44324
rect 46610 44268 46620 44324
rect 46676 44268 46686 44324
rect 49746 44268 49756 44324
rect 49812 44268 57596 44324
rect 57652 44268 57662 44324
rect 41682 44156 41692 44212
rect 41748 44156 43596 44212
rect 43652 44156 45388 44212
rect 45444 44156 45454 44212
rect 46620 44100 46676 44268
rect 55458 44156 55468 44212
rect 55524 44156 58268 44212
rect 58324 44156 58334 44212
rect 60050 44156 60060 44212
rect 60116 44156 62524 44212
rect 62580 44156 62590 44212
rect 25778 44044 25788 44100
rect 25844 44044 28364 44100
rect 28420 44044 28430 44100
rect 33618 44044 33628 44100
rect 33684 44044 35980 44100
rect 36036 44044 36046 44100
rect 46620 44044 57596 44100
rect 57652 44044 57662 44100
rect 37650 43932 37660 43988
rect 37716 43932 42812 43988
rect 42868 43932 42878 43988
rect 45378 43932 45388 43988
rect 45444 43932 46396 43988
rect 46452 43932 46462 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 24210 43820 24220 43876
rect 24276 43820 24780 43876
rect 24836 43820 24846 43876
rect 40898 43820 40908 43876
rect 40964 43820 45948 43876
rect 46004 43820 46014 43876
rect 49074 43820 49084 43876
rect 49140 43820 49756 43876
rect 49812 43820 49822 43876
rect 48934 43708 48972 43764
rect 49028 43708 50316 43764
rect 50372 43708 52780 43764
rect 52836 43708 52846 43764
rect 56018 43708 56028 43764
rect 56084 43708 56812 43764
rect 56868 43708 58492 43764
rect 58548 43708 59500 43764
rect 59556 43708 59566 43764
rect 48972 43652 49028 43708
rect 14802 43596 14812 43652
rect 14868 43596 20860 43652
rect 20916 43596 20926 43652
rect 28690 43596 28700 43652
rect 28756 43596 33068 43652
rect 33124 43596 33134 43652
rect 47730 43596 47740 43652
rect 47796 43596 48188 43652
rect 48244 43596 49028 43652
rect 49522 43596 49532 43652
rect 49588 43596 49980 43652
rect 50036 43596 50876 43652
rect 50932 43596 51548 43652
rect 51604 43596 51614 43652
rect 51762 43596 51772 43652
rect 51828 43596 54908 43652
rect 54964 43596 54974 43652
rect 56130 43596 56140 43652
rect 56196 43596 61404 43652
rect 61460 43596 61470 43652
rect 36530 43484 36540 43540
rect 36596 43484 41020 43540
rect 41076 43484 41086 43540
rect 47394 43484 47404 43540
rect 47460 43484 50988 43540
rect 51044 43484 51054 43540
rect 51426 43484 51436 43540
rect 51492 43484 52612 43540
rect 52770 43484 52780 43540
rect 52836 43484 54684 43540
rect 54740 43484 56700 43540
rect 56756 43484 56766 43540
rect 52556 43428 52612 43484
rect 32386 43372 32396 43428
rect 32452 43372 33292 43428
rect 33348 43372 33358 43428
rect 45154 43372 45164 43428
rect 45220 43372 48860 43428
rect 48916 43372 49196 43428
rect 49252 43372 49262 43428
rect 50194 43372 50204 43428
rect 50260 43372 51548 43428
rect 51604 43372 51614 43428
rect 52556 43372 55132 43428
rect 55188 43372 57148 43428
rect 57204 43372 59276 43428
rect 59332 43372 59342 43428
rect 60386 43372 60396 43428
rect 60452 43372 60462 43428
rect 60396 43316 60452 43372
rect 53218 43260 53228 43316
rect 53284 43260 60452 43316
rect 48290 43148 48300 43204
rect 48356 43148 58828 43204
rect 58884 43148 58894 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 18386 42924 18396 42980
rect 18452 42924 21196 42980
rect 21252 42924 21262 42980
rect 23090 42812 23100 42868
rect 23156 42812 28252 42868
rect 28308 42812 28318 42868
rect 41458 42812 41468 42868
rect 41524 42812 42588 42868
rect 42644 42812 42654 42868
rect 57026 42812 57036 42868
rect 57092 42812 61516 42868
rect 61572 42812 61582 42868
rect 29250 42700 29260 42756
rect 29316 42700 31388 42756
rect 31444 42700 31454 42756
rect 36866 42700 36876 42756
rect 36932 42700 39004 42756
rect 39060 42700 39070 42756
rect 44930 42700 44940 42756
rect 44996 42700 47740 42756
rect 47796 42700 47806 42756
rect 15922 42588 15932 42644
rect 15988 42588 23772 42644
rect 23828 42588 23838 42644
rect 48402 42588 48412 42644
rect 48468 42588 55468 42644
rect 56242 42588 56252 42644
rect 56308 42588 62524 42644
rect 62580 42588 62590 42644
rect 27906 42476 27916 42532
rect 27972 42476 28476 42532
rect 28532 42476 28542 42532
rect 46498 42476 46508 42532
rect 46564 42476 47628 42532
rect 47684 42476 47694 42532
rect 55412 42420 55468 42588
rect 55412 42364 58828 42420
rect 58884 42364 58894 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 22082 42252 22092 42308
rect 22148 42252 25004 42308
rect 25060 42252 25070 42308
rect 25890 42252 25900 42308
rect 25956 42252 30268 42308
rect 30324 42252 30334 42308
rect 55346 42140 55356 42196
rect 55412 42140 59276 42196
rect 59332 42140 59342 42196
rect 16146 42028 16156 42084
rect 16212 42028 16940 42084
rect 16996 42028 17006 42084
rect 17826 42028 17836 42084
rect 17892 42028 21756 42084
rect 21812 42028 21822 42084
rect 26562 42028 26572 42084
rect 26628 42028 29372 42084
rect 29428 42028 29438 42084
rect 36306 42028 36316 42084
rect 36372 42028 41804 42084
rect 41860 42028 41870 42084
rect 56242 42028 56252 42084
rect 56308 42028 61404 42084
rect 61460 42028 61470 42084
rect 15810 41916 15820 41972
rect 15876 41916 20636 41972
rect 20692 41916 20702 41972
rect 21522 41916 21532 41972
rect 21588 41916 23996 41972
rect 24052 41916 24062 41972
rect 25452 41916 27132 41972
rect 27188 41916 28140 41972
rect 28196 41916 28206 41972
rect 38994 41916 39004 41972
rect 39060 41916 39564 41972
rect 39620 41916 40796 41972
rect 40852 41916 40862 41972
rect 45266 41916 45276 41972
rect 45332 41916 55468 41972
rect 56690 41916 56700 41972
rect 56756 41916 59500 41972
rect 59556 41916 59566 41972
rect 25452 41860 25508 41916
rect 55412 41860 55468 41916
rect 18722 41804 18732 41860
rect 18788 41804 20972 41860
rect 21028 41804 21038 41860
rect 23650 41804 23660 41860
rect 23716 41804 24332 41860
rect 24388 41804 24780 41860
rect 24836 41804 25452 41860
rect 25508 41804 25518 41860
rect 25666 41804 25676 41860
rect 25732 41804 32620 41860
rect 32676 41804 32686 41860
rect 55412 41804 57596 41860
rect 57652 41804 57662 41860
rect 59378 41804 59388 41860
rect 59444 41804 62188 41860
rect 62244 41804 62254 41860
rect 25778 41692 25788 41748
rect 25844 41692 26460 41748
rect 26516 41692 26526 41748
rect 28018 41692 28028 41748
rect 28084 41692 31164 41748
rect 31220 41692 31230 41748
rect 32386 41692 32396 41748
rect 32452 41692 34076 41748
rect 34132 41692 34972 41748
rect 35028 41692 36092 41748
rect 36148 41692 36988 41748
rect 37044 41692 37054 41748
rect 59602 41692 59612 41748
rect 59668 41692 62412 41748
rect 62468 41692 62972 41748
rect 63028 41692 63038 41748
rect 16818 41580 16828 41636
rect 16884 41580 17724 41636
rect 17780 41580 17790 41636
rect 18722 41580 18732 41636
rect 18788 41580 27916 41636
rect 27972 41580 27982 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 19730 41244 19740 41300
rect 19796 41244 21812 41300
rect 21970 41244 21980 41300
rect 22036 41244 24444 41300
rect 24500 41244 24510 41300
rect 26674 41244 26684 41300
rect 26740 41244 26908 41300
rect 36642 41244 36652 41300
rect 36708 41244 38220 41300
rect 38276 41244 38286 41300
rect 40002 41244 40012 41300
rect 40068 41244 43372 41300
rect 43428 41244 43438 41300
rect 43922 41244 43932 41300
rect 43988 41244 45500 41300
rect 45556 41244 45566 41300
rect 46162 41244 46172 41300
rect 46228 41244 46844 41300
rect 46900 41244 46910 41300
rect 51426 41244 51436 41300
rect 51492 41244 52108 41300
rect 52164 41244 55580 41300
rect 55636 41244 56812 41300
rect 56868 41244 56878 41300
rect 21756 41076 21812 41244
rect 26852 41188 26908 41244
rect 26852 41132 32732 41188
rect 32788 41132 32798 41188
rect 42466 41132 42476 41188
rect 42532 41132 47908 41188
rect 48066 41132 48076 41188
rect 48132 41132 60396 41188
rect 60452 41132 60462 41188
rect 47852 41076 47908 41132
rect 15922 41020 15932 41076
rect 15988 41020 21084 41076
rect 21140 41020 21150 41076
rect 21756 41020 29484 41076
rect 29540 41020 29550 41076
rect 38546 41020 38556 41076
rect 38612 41020 40124 41076
rect 40180 41020 43708 41076
rect 43764 41020 43774 41076
rect 45154 41020 45164 41076
rect 45220 41020 45230 41076
rect 47852 41020 58492 41076
rect 58548 41020 58558 41076
rect 45164 40964 45220 41020
rect 20738 40908 20748 40964
rect 20804 40908 23548 40964
rect 23604 40908 27132 40964
rect 27188 40908 27198 40964
rect 35186 40908 35196 40964
rect 35252 40908 37100 40964
rect 37156 40908 37166 40964
rect 43138 40908 43148 40964
rect 43204 40908 45220 40964
rect 51090 40908 51100 40964
rect 51156 40908 61404 40964
rect 61460 40908 61470 40964
rect 43698 40796 43708 40852
rect 43764 40796 44044 40852
rect 44100 40796 45724 40852
rect 45780 40796 45790 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 28466 40684 28476 40740
rect 28532 40684 30604 40740
rect 30660 40684 30670 40740
rect 56130 40684 56140 40740
rect 56196 40684 62524 40740
rect 62580 40684 62590 40740
rect 10770 40572 10780 40628
rect 10836 40572 11676 40628
rect 11732 40572 11742 40628
rect 12002 40572 12012 40628
rect 12068 40572 17276 40628
rect 17332 40572 17342 40628
rect 22866 40572 22876 40628
rect 22932 40572 25788 40628
rect 25844 40572 25854 40628
rect 33954 40572 33964 40628
rect 34020 40572 37212 40628
rect 37268 40572 37278 40628
rect 47954 40572 47964 40628
rect 48020 40572 57092 40628
rect 57036 40516 57092 40572
rect 16594 40460 16604 40516
rect 16660 40460 17836 40516
rect 17892 40460 17902 40516
rect 22306 40460 22316 40516
rect 22372 40460 25564 40516
rect 25620 40460 25630 40516
rect 28690 40460 28700 40516
rect 28756 40460 30604 40516
rect 30660 40460 31724 40516
rect 31780 40460 32284 40516
rect 32340 40460 32350 40516
rect 42802 40460 42812 40516
rect 42868 40460 55468 40516
rect 55524 40460 55534 40516
rect 57036 40460 58828 40516
rect 58884 40460 58894 40516
rect 9986 40348 9996 40404
rect 10052 40348 12236 40404
rect 12292 40348 12302 40404
rect 16258 40348 16268 40404
rect 16324 40348 17500 40404
rect 17556 40348 17566 40404
rect 17714 40348 17724 40404
rect 17780 40348 24108 40404
rect 24164 40348 24174 40404
rect 24658 40348 24668 40404
rect 24724 40348 28588 40404
rect 28644 40348 28924 40404
rect 28980 40348 31164 40404
rect 31220 40348 31948 40404
rect 32004 40348 32014 40404
rect 38546 40348 38556 40404
rect 38612 40348 42700 40404
rect 42756 40348 42766 40404
rect 44930 40348 44940 40404
rect 44996 40348 47012 40404
rect 53106 40348 53116 40404
rect 53172 40348 61516 40404
rect 61572 40348 61582 40404
rect 46956 40292 47012 40348
rect 19842 40236 19852 40292
rect 19908 40236 25340 40292
rect 25396 40236 25406 40292
rect 32162 40236 32172 40292
rect 32228 40236 33516 40292
rect 33572 40236 33582 40292
rect 34514 40236 34524 40292
rect 34580 40236 38444 40292
rect 38500 40236 38510 40292
rect 46956 40236 54012 40292
rect 54068 40236 54078 40292
rect 21746 40124 21756 40180
rect 21812 40124 24780 40180
rect 24836 40124 24846 40180
rect 50306 40124 50316 40180
rect 50372 40124 51436 40180
rect 51492 40124 51502 40180
rect 53666 40124 53676 40180
rect 53732 40124 61740 40180
rect 61796 40124 61806 40180
rect 50194 40012 50204 40068
rect 50260 40012 60396 40068
rect 60452 40012 60462 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 11890 39900 11900 39956
rect 11956 39900 13916 39956
rect 13972 39900 13982 39956
rect 16706 39900 16716 39956
rect 16772 39900 24780 39956
rect 24836 39900 24846 39956
rect 30930 39900 30940 39956
rect 30996 39900 32060 39956
rect 32116 39900 32126 39956
rect 48402 39900 48412 39956
rect 48468 39900 58940 39956
rect 58996 39900 59006 39956
rect 29922 39788 29932 39844
rect 29988 39788 32620 39844
rect 32676 39788 32686 39844
rect 40908 39788 57596 39844
rect 57652 39788 57662 39844
rect 9090 39676 9100 39732
rect 9156 39676 14700 39732
rect 14756 39676 14766 39732
rect 16818 39676 16828 39732
rect 16884 39676 20188 39732
rect 27906 39676 27916 39732
rect 27972 39676 29148 39732
rect 29204 39676 29214 39732
rect 20132 39620 20188 39676
rect 40908 39620 40964 39788
rect 44482 39676 44492 39732
rect 44548 39676 49196 39732
rect 49252 39676 52444 39732
rect 52500 39676 53004 39732
rect 53060 39676 53788 39732
rect 53844 39676 53854 39732
rect 54002 39676 54012 39732
rect 54068 39676 57932 39732
rect 57988 39676 57998 39732
rect 11890 39564 11900 39620
rect 11956 39564 17724 39620
rect 17780 39564 17790 39620
rect 20132 39564 24332 39620
rect 24388 39564 24398 39620
rect 40898 39564 40908 39620
rect 40964 39564 40974 39620
rect 41682 39564 41692 39620
rect 41748 39564 43708 39620
rect 43764 39564 43774 39620
rect 45378 39564 45388 39620
rect 45444 39564 57596 39620
rect 57652 39564 57662 39620
rect 20178 39452 20188 39508
rect 20244 39452 21308 39508
rect 21364 39452 21374 39508
rect 21634 39452 21644 39508
rect 21700 39452 22428 39508
rect 22484 39452 22876 39508
rect 22932 39452 22942 39508
rect 10770 39340 10780 39396
rect 10836 39340 20972 39396
rect 21028 39340 21038 39396
rect 56690 39340 56700 39396
rect 56756 39340 61404 39396
rect 61460 39340 61470 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 40898 39116 40908 39172
rect 40964 39116 41244 39172
rect 41300 39116 41804 39172
rect 41860 39116 41870 39172
rect 12002 39004 12012 39060
rect 12068 39004 22204 39060
rect 22260 39004 22270 39060
rect 41570 39004 41580 39060
rect 41636 39004 45388 39060
rect 45444 39004 57484 39060
rect 57540 39004 57550 39060
rect 10994 38892 11004 38948
rect 11060 38892 20748 38948
rect 20804 38892 20814 38948
rect 28802 38892 28812 38948
rect 28868 38892 31948 38948
rect 32004 38892 32014 38948
rect 33282 38892 33292 38948
rect 33348 38892 37436 38948
rect 37492 38892 40236 38948
rect 40292 38892 43708 38948
rect 47058 38892 47068 38948
rect 47124 38892 47134 38948
rect 53218 38892 53228 38948
rect 53284 38892 62524 38948
rect 62580 38892 62590 38948
rect 43652 38836 43708 38892
rect 13010 38780 13020 38836
rect 13076 38780 13804 38836
rect 13860 38780 13870 38836
rect 31154 38780 31164 38836
rect 31220 38780 38668 38836
rect 42690 38780 42700 38836
rect 42756 38780 42766 38836
rect 43652 38780 44380 38836
rect 44436 38780 45052 38836
rect 45108 38780 45118 38836
rect 38612 38724 38668 38780
rect 42700 38724 42756 38780
rect 47068 38724 47124 38892
rect 53778 38780 53788 38836
rect 53844 38780 56700 38836
rect 56756 38780 56766 38836
rect 13458 38668 13468 38724
rect 13524 38668 15148 38724
rect 15204 38668 15820 38724
rect 15876 38668 17164 38724
rect 17220 38668 18396 38724
rect 18452 38668 18462 38724
rect 20132 38668 20300 38724
rect 20356 38668 22764 38724
rect 22820 38668 22830 38724
rect 28018 38668 28028 38724
rect 28084 38668 33292 38724
rect 33348 38668 33358 38724
rect 38612 38668 42756 38724
rect 43026 38668 43036 38724
rect 43092 38668 47124 38724
rect 47394 38668 47404 38724
rect 47460 38668 48972 38724
rect 49028 38668 49038 38724
rect 20132 38612 20188 38668
rect 15026 38556 15036 38612
rect 15092 38556 20188 38612
rect 39666 38444 39676 38500
rect 39732 38444 49644 38500
rect 49700 38444 49710 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 7970 38332 7980 38388
rect 8036 38332 9884 38388
rect 9940 38332 9950 38388
rect 19394 38332 19404 38388
rect 19460 38332 27692 38388
rect 27748 38332 27758 38388
rect 49186 38332 49196 38388
rect 49252 38332 60396 38388
rect 60452 38332 60462 38388
rect 18834 38220 18844 38276
rect 18900 38220 28364 38276
rect 28420 38220 28430 38276
rect 35074 38220 35084 38276
rect 35140 38220 42924 38276
rect 42980 38220 42990 38276
rect 45378 38220 45388 38276
rect 45444 38220 57596 38276
rect 57652 38220 57662 38276
rect 6962 38108 6972 38164
rect 7028 38108 12908 38164
rect 12964 38108 12974 38164
rect 22642 38108 22652 38164
rect 22708 38108 30940 38164
rect 30996 38108 31006 38164
rect 37426 38108 37436 38164
rect 37492 38108 37996 38164
rect 38052 38108 38062 38164
rect 53330 38108 53340 38164
rect 53396 38108 61516 38164
rect 61572 38108 61582 38164
rect 19506 37996 19516 38052
rect 19572 37996 21140 38052
rect 21298 37996 21308 38052
rect 21364 37996 23996 38052
rect 24052 37996 24668 38052
rect 24724 37996 24734 38052
rect 41794 37996 41804 38052
rect 41860 37996 52780 38052
rect 52836 37996 52846 38052
rect 58818 37996 58828 38052
rect 58884 37996 58894 38052
rect 21084 37940 21140 37996
rect 58828 37940 58884 37996
rect 19618 37884 19628 37940
rect 19684 37884 20412 37940
rect 20468 37884 20478 37940
rect 21084 37884 24556 37940
rect 24612 37884 24622 37940
rect 29138 37884 29148 37940
rect 29204 37884 30828 37940
rect 30884 37884 30894 37940
rect 31154 37884 31164 37940
rect 31220 37884 33404 37940
rect 33460 37884 33470 37940
rect 42130 37884 42140 37940
rect 42196 37884 42924 37940
rect 42980 37884 42990 37940
rect 43138 37884 43148 37940
rect 43204 37884 43820 37940
rect 43876 37884 45500 37940
rect 45556 37884 45566 37940
rect 50372 37884 58884 37940
rect 50372 37828 50428 37884
rect 8082 37772 8092 37828
rect 8148 37772 13020 37828
rect 13076 37772 13086 37828
rect 19628 37772 19740 37828
rect 19796 37772 20636 37828
rect 20692 37772 21644 37828
rect 21700 37772 21710 37828
rect 48402 37772 48412 37828
rect 48468 37772 50428 37828
rect 52210 37772 52220 37828
rect 52276 37772 61404 37828
rect 61460 37772 61470 37828
rect 19628 37492 19684 37772
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 10994 37436 11004 37492
rect 11060 37436 19180 37492
rect 19236 37436 19246 37492
rect 19628 37436 19740 37492
rect 19796 37436 19806 37492
rect 38612 37436 39452 37492
rect 39508 37436 39518 37492
rect 47842 37436 47852 37492
rect 47908 37436 48972 37492
rect 49028 37436 49038 37492
rect 6962 37324 6972 37380
rect 7028 37324 11900 37380
rect 11956 37324 11966 37380
rect 24210 37324 24220 37380
rect 24276 37324 25228 37380
rect 25284 37324 25294 37380
rect 33394 37324 33404 37380
rect 33460 37324 34188 37380
rect 34244 37324 37436 37380
rect 37492 37324 37502 37380
rect 5170 37212 5180 37268
rect 5236 37212 8652 37268
rect 8708 37212 8718 37268
rect 9314 37212 9324 37268
rect 9380 37212 13244 37268
rect 13300 37212 13310 37268
rect 16258 37212 16268 37268
rect 16324 37212 17388 37268
rect 17444 37212 17454 37268
rect 20132 37212 21644 37268
rect 21700 37212 21710 37268
rect 27794 37212 27804 37268
rect 27860 37212 29484 37268
rect 29540 37212 29550 37268
rect 38546 37212 38556 37268
rect 38612 37212 38668 37436
rect 45490 37324 45500 37380
rect 45556 37324 47292 37380
rect 47348 37324 47964 37380
rect 48020 37324 48524 37380
rect 48580 37324 48590 37380
rect 48850 37324 48860 37380
rect 48916 37324 49532 37380
rect 49588 37324 49598 37380
rect 53106 37324 53116 37380
rect 53172 37324 53900 37380
rect 53956 37324 53966 37380
rect 54674 37324 54684 37380
rect 54740 37324 55580 37380
rect 55636 37324 56700 37380
rect 56756 37324 56766 37380
rect 54226 37212 54236 37268
rect 54292 37212 55468 37268
rect 55524 37212 55534 37268
rect 20132 37156 20188 37212
rect 7970 37100 7980 37156
rect 8036 37100 8428 37156
rect 12002 37100 12012 37156
rect 12068 37100 20188 37156
rect 40338 37100 40348 37156
rect 40404 37100 43148 37156
rect 43204 37100 43214 37156
rect 44818 37100 44828 37156
rect 44884 37100 46732 37156
rect 46788 37100 48188 37156
rect 48244 37100 48254 37156
rect 50642 37100 50652 37156
rect 50708 37100 60396 37156
rect 60452 37100 60462 37156
rect 8372 37044 8428 37100
rect 8372 36988 13916 37044
rect 13972 36988 13982 37044
rect 41692 36988 42196 37044
rect 48402 36988 48412 37044
rect 48468 36988 58828 37044
rect 58884 36988 58894 37044
rect 41692 36932 41748 36988
rect 42140 36932 42196 36988
rect 25330 36876 25340 36932
rect 25396 36876 29596 36932
rect 29652 36876 29662 36932
rect 38612 36876 41748 36932
rect 41906 36876 41916 36932
rect 41972 36876 41982 36932
rect 42140 36876 43036 36932
rect 43092 36876 43102 36932
rect 50372 36876 57596 36932
rect 57652 36876 57662 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 10210 36764 10220 36820
rect 10276 36764 12796 36820
rect 12852 36764 14028 36820
rect 14084 36764 14812 36820
rect 14868 36764 14878 36820
rect 38612 36708 38668 36876
rect 41916 36820 41972 36876
rect 50372 36820 50428 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 7074 36652 7084 36708
rect 7140 36652 11116 36708
rect 11172 36652 11182 36708
rect 12450 36652 12460 36708
rect 12516 36652 15820 36708
rect 15876 36652 15886 36708
rect 36530 36652 36540 36708
rect 36596 36652 38668 36708
rect 38780 36764 41972 36820
rect 45266 36764 45276 36820
rect 45332 36764 50428 36820
rect 56242 36764 56252 36820
rect 56308 36764 62188 36820
rect 38780 36596 38836 36764
rect 62132 36708 62188 36764
rect 41682 36652 41692 36708
rect 41748 36652 50876 36708
rect 50932 36652 50942 36708
rect 53004 36652 58492 36708
rect 58548 36652 58558 36708
rect 62132 36652 62524 36708
rect 62580 36652 62590 36708
rect 53004 36596 53060 36652
rect 8082 36540 8092 36596
rect 8148 36540 18228 36596
rect 22642 36540 22652 36596
rect 22708 36540 31164 36596
rect 31220 36540 31230 36596
rect 33506 36540 33516 36596
rect 33572 36540 38836 36596
rect 38892 36540 39676 36596
rect 39732 36540 41020 36596
rect 41076 36540 42028 36596
rect 42084 36540 42812 36596
rect 42868 36540 44828 36596
rect 44884 36540 44894 36596
rect 46386 36540 46396 36596
rect 46452 36540 53060 36596
rect 53218 36540 53228 36596
rect 53284 36540 61516 36596
rect 61572 36540 61582 36596
rect 18172 36484 18228 36540
rect 38892 36484 38948 36540
rect 7970 36428 7980 36484
rect 8036 36428 9884 36484
rect 9940 36428 9950 36484
rect 18162 36428 18172 36484
rect 18228 36428 18238 36484
rect 18946 36428 18956 36484
rect 19012 36428 24556 36484
rect 24612 36428 24622 36484
rect 26450 36428 26460 36484
rect 26516 36428 32732 36484
rect 32788 36428 32798 36484
rect 33058 36428 33068 36484
rect 33124 36428 34860 36484
rect 34916 36428 35644 36484
rect 35700 36428 37772 36484
rect 37828 36428 38892 36484
rect 38948 36428 38958 36484
rect 44370 36428 44380 36484
rect 44436 36428 47068 36484
rect 47124 36428 48076 36484
rect 48132 36428 48142 36484
rect 50418 36428 50428 36484
rect 50484 36428 52556 36484
rect 52612 36428 56588 36484
rect 56644 36428 56654 36484
rect 0 36372 800 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 12450 36316 12460 36372
rect 12516 36316 13692 36372
rect 13748 36316 13758 36372
rect 19506 36316 19516 36372
rect 19572 36316 20412 36372
rect 20468 36316 22092 36372
rect 22148 36316 22158 36372
rect 35970 36316 35980 36372
rect 36036 36316 36988 36372
rect 37044 36316 37054 36372
rect 40114 36316 40124 36372
rect 40180 36316 40908 36372
rect 40964 36316 40974 36372
rect 53666 36316 53676 36372
rect 53732 36316 62524 36372
rect 62580 36316 62590 36372
rect 0 36288 800 36316
rect 10882 36204 10892 36260
rect 10948 36204 29932 36260
rect 29988 36204 29998 36260
rect 7074 36092 7084 36148
rect 7140 36092 17052 36148
rect 17108 36092 17118 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 12674 35980 12684 36036
rect 12740 35980 14588 36036
rect 14644 35980 14654 36036
rect 35522 35980 35532 36036
rect 35588 35980 45836 36036
rect 45892 35980 45902 36036
rect 2034 35868 2044 35924
rect 2100 35868 23212 35924
rect 23268 35868 23278 35924
rect 31826 35868 31836 35924
rect 31892 35812 31948 35924
rect 44482 35868 44492 35924
rect 44548 35868 50428 35924
rect 53666 35868 53676 35924
rect 53732 35868 54460 35924
rect 54516 35868 54526 35924
rect 50372 35812 50428 35868
rect 4162 35756 4172 35812
rect 4228 35756 12796 35812
rect 12852 35756 12862 35812
rect 14802 35756 14812 35812
rect 14868 35756 16044 35812
rect 16100 35756 16716 35812
rect 16772 35756 17612 35812
rect 17668 35756 18172 35812
rect 18228 35756 18238 35812
rect 31892 35756 33068 35812
rect 33124 35756 33134 35812
rect 33394 35756 33404 35812
rect 33460 35756 34076 35812
rect 34132 35756 34142 35812
rect 50372 35756 58828 35812
rect 58884 35756 58894 35812
rect 33404 35700 33460 35756
rect 3042 35644 3052 35700
rect 3108 35644 11228 35700
rect 11284 35644 11294 35700
rect 20132 35644 22876 35700
rect 22932 35644 24220 35700
rect 24276 35644 24286 35700
rect 24434 35644 24444 35700
rect 24500 35644 25340 35700
rect 25396 35644 26012 35700
rect 26068 35644 26078 35700
rect 32386 35644 32396 35700
rect 32452 35644 33460 35700
rect 41458 35644 41468 35700
rect 41524 35644 54348 35700
rect 54404 35644 54414 35700
rect 20132 35588 20188 35644
rect 9874 35532 9884 35588
rect 9940 35532 11452 35588
rect 11508 35532 11518 35588
rect 17154 35532 17164 35588
rect 17220 35532 18956 35588
rect 19012 35532 20188 35588
rect 47618 35532 47628 35588
rect 47684 35532 60396 35588
rect 60452 35532 60462 35588
rect 6962 35420 6972 35476
rect 7028 35420 15148 35476
rect 15204 35420 15214 35476
rect 54898 35420 54908 35476
rect 54964 35420 55580 35476
rect 55636 35420 59388 35476
rect 59444 35420 59454 35476
rect 5170 35308 5180 35364
rect 5236 35308 13020 35364
rect 13076 35308 13086 35364
rect 16482 35308 16492 35364
rect 16548 35308 18396 35364
rect 18452 35308 18462 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 54908 35252 54964 35420
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 21522 35196 21532 35252
rect 21588 35196 31836 35252
rect 31892 35196 31902 35252
rect 50418 35196 50428 35252
rect 50484 35196 50988 35252
rect 51044 35196 51324 35252
rect 51380 35196 52108 35252
rect 52164 35196 54572 35252
rect 54628 35196 54964 35252
rect 41122 35084 41132 35140
rect 41188 35084 50428 35140
rect 56354 35084 56364 35140
rect 56420 35084 61404 35140
rect 61460 35084 61470 35140
rect 50372 35028 50428 35084
rect 7298 34972 7308 35028
rect 7364 34972 17780 35028
rect 24210 34972 24220 35028
rect 24276 34972 26348 35028
rect 26404 34972 28028 35028
rect 28084 34972 28094 35028
rect 38546 34972 38556 35028
rect 17724 34916 17780 34972
rect 3042 34860 3052 34916
rect 3108 34860 12236 34916
rect 12292 34860 12302 34916
rect 15250 34860 15260 34916
rect 15316 34860 17164 34916
rect 17220 34860 17230 34916
rect 17714 34860 17724 34916
rect 17780 34860 17790 34916
rect 31892 34860 35196 34916
rect 35252 34860 37884 34916
rect 37940 34860 37950 34916
rect 31892 34804 31948 34860
rect 6290 34748 6300 34804
rect 6356 34748 20188 34804
rect 28466 34748 28476 34804
rect 28532 34748 31948 34804
rect 38612 34804 38668 35028
rect 50372 34972 57596 35028
rect 57652 34972 57662 35028
rect 38612 34748 41804 34804
rect 41860 34748 42924 34804
rect 42980 34748 43596 34804
rect 43652 34748 43662 34804
rect 56130 34748 56140 34804
rect 56196 34748 58828 34804
rect 58884 34748 58894 34804
rect 62514 34748 62524 34804
rect 62580 34748 62590 34804
rect 20132 34692 20188 34748
rect 62524 34692 62580 34748
rect 11666 34636 11676 34692
rect 11732 34636 13468 34692
rect 13524 34636 13534 34692
rect 20132 34636 20972 34692
rect 21028 34636 21038 34692
rect 50642 34636 50652 34692
rect 50708 34636 55188 34692
rect 55346 34636 55356 34692
rect 55412 34636 59500 34692
rect 59556 34636 59566 34692
rect 62132 34636 62580 34692
rect 55132 34580 55188 34636
rect 62132 34580 62188 34636
rect 51884 34524 53956 34580
rect 55132 34524 62188 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 36082 34412 36092 34468
rect 36148 34412 36540 34468
rect 36596 34412 48748 34468
rect 48804 34412 48814 34468
rect 51884 34356 51940 34524
rect 53900 34468 53956 34524
rect 7970 34300 7980 34356
rect 8036 34300 17836 34356
rect 17892 34300 17902 34356
rect 31266 34300 31276 34356
rect 31332 34300 31948 34356
rect 49298 34300 49308 34356
rect 49364 34300 51940 34356
rect 51996 34412 53676 34468
rect 53732 34412 53742 34468
rect 53900 34412 61516 34468
rect 61572 34412 61582 34468
rect 31892 34244 31948 34300
rect 51996 34244 52052 34412
rect 52322 34300 52332 34356
rect 52388 34300 61404 34356
rect 61460 34300 61470 34356
rect 6962 34188 6972 34244
rect 7028 34188 20860 34244
rect 20916 34188 20926 34244
rect 31892 34188 32060 34244
rect 32116 34188 32126 34244
rect 41468 34188 52052 34244
rect 52668 34188 58828 34244
rect 58884 34188 58894 34244
rect 41468 34132 41524 34188
rect 4162 34076 4172 34132
rect 4228 34076 9100 34132
rect 9156 34076 9166 34132
rect 14130 34076 14140 34132
rect 14196 34076 14206 34132
rect 20738 34076 20748 34132
rect 20804 34076 21980 34132
rect 22036 34076 22046 34132
rect 37426 34076 37436 34132
rect 37492 34076 41132 34132
rect 41188 34076 41198 34132
rect 41458 34076 41468 34132
rect 41524 34076 41534 34132
rect 48850 34076 48860 34132
rect 48916 34076 52444 34132
rect 52500 34076 52510 34132
rect 7970 33964 7980 34020
rect 8036 33964 13580 34020
rect 13636 33964 13646 34020
rect 14140 33908 14196 34076
rect 52668 34020 52724 34188
rect 14690 33964 14700 34020
rect 14756 33964 15820 34020
rect 15876 33964 16268 34020
rect 16324 33964 16334 34020
rect 44482 33964 44492 34020
rect 44548 33964 52724 34020
rect 57586 33964 57596 34020
rect 57652 33964 57662 34020
rect 57596 33908 57652 33964
rect 5170 33852 5180 33908
rect 5236 33852 14196 33908
rect 21746 33852 21756 33908
rect 21812 33852 32956 33908
rect 33012 33852 33022 33908
rect 40450 33852 40460 33908
rect 40516 33852 40526 33908
rect 47058 33852 47068 33908
rect 47124 33852 57652 33908
rect 7858 33740 7868 33796
rect 7924 33740 21644 33796
rect 21700 33740 21710 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 40460 33684 40516 33852
rect 43922 33740 43932 33796
rect 43988 33740 45052 33796
rect 45108 33740 46060 33796
rect 46116 33740 47964 33796
rect 48020 33740 51436 33796
rect 51492 33740 51502 33796
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 40460 33628 48804 33684
rect 53106 33628 53116 33684
rect 53172 33628 53844 33684
rect 4274 33516 4284 33572
rect 4340 33516 8316 33572
rect 8372 33516 8382 33572
rect 10546 33516 10556 33572
rect 10612 33516 11340 33572
rect 11396 33516 13804 33572
rect 13860 33516 15036 33572
rect 15092 33516 15102 33572
rect 22754 33516 22764 33572
rect 22820 33516 23548 33572
rect 23604 33516 23614 33572
rect 41906 33516 41916 33572
rect 41972 33516 47068 33572
rect 47124 33516 47134 33572
rect 48748 33460 48804 33628
rect 53788 33572 53844 33628
rect 53788 33516 61516 33572
rect 61572 33516 61582 33572
rect 4050 33404 4060 33460
rect 4116 33404 13692 33460
rect 13748 33404 13758 33460
rect 20402 33404 20412 33460
rect 20468 33404 21420 33460
rect 21476 33404 21486 33460
rect 32498 33404 32508 33460
rect 32564 33404 35084 33460
rect 35140 33404 35644 33460
rect 35700 33404 36428 33460
rect 36484 33404 36494 33460
rect 39890 33404 39900 33460
rect 39956 33404 42924 33460
rect 42980 33404 42990 33460
rect 43250 33404 43260 33460
rect 43316 33404 43932 33460
rect 43988 33404 43998 33460
rect 48748 33404 54684 33460
rect 54740 33404 54750 33460
rect 3826 33292 3836 33348
rect 3892 33292 12124 33348
rect 12180 33292 12190 33348
rect 20066 33292 20076 33348
rect 20132 33292 22540 33348
rect 22596 33292 22606 33348
rect 25778 33292 25788 33348
rect 25844 33292 27692 33348
rect 27748 33292 27758 33348
rect 30594 33292 30604 33348
rect 30660 33292 31836 33348
rect 31892 33292 36540 33348
rect 36596 33292 40348 33348
rect 40404 33292 41244 33348
rect 41300 33292 41310 33348
rect 45378 33292 45388 33348
rect 45444 33292 45454 33348
rect 49186 33292 49196 33348
rect 49252 33292 60396 33348
rect 60452 33292 60462 33348
rect 30146 33180 30156 33236
rect 30212 33180 34524 33236
rect 34580 33180 36092 33236
rect 36148 33180 37324 33236
rect 37380 33180 37390 33236
rect 45388 33124 45444 33292
rect 46274 33180 46284 33236
rect 46340 33180 47628 33236
rect 47684 33180 47694 33236
rect 48738 33180 48748 33236
rect 48804 33180 52052 33236
rect 62514 33180 62524 33236
rect 62580 33180 62590 33236
rect 3042 33068 3052 33124
rect 3108 33068 16156 33124
rect 16212 33068 16222 33124
rect 39890 33068 39900 33124
rect 39956 33068 43820 33124
rect 43876 33068 43886 33124
rect 45388 33068 51940 33124
rect 4162 32956 4172 33012
rect 4228 32956 17052 33012
rect 17108 32956 17118 33012
rect 24546 32956 24556 33012
rect 24612 32956 28700 33012
rect 28756 32956 28766 33012
rect 39330 32956 39340 33012
rect 39396 32956 47180 33012
rect 47236 32956 47246 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 51884 32900 51940 33068
rect 51996 33012 52052 33180
rect 52210 33068 52220 33124
rect 52276 33068 61404 33124
rect 61460 33068 61470 33124
rect 62524 33012 62580 33180
rect 51996 32956 56476 33012
rect 56532 32956 56542 33012
rect 62132 32956 62580 33012
rect 62132 32900 62188 32956
rect 42914 32844 42924 32900
rect 42980 32844 43708 32900
rect 43764 32844 43774 32900
rect 51884 32844 53900 32900
rect 53956 32844 53966 32900
rect 54226 32844 54236 32900
rect 54292 32844 62188 32900
rect 6626 32732 6636 32788
rect 6692 32732 21196 32788
rect 21252 32732 21262 32788
rect 36092 32732 44212 32788
rect 44930 32732 44940 32788
rect 44996 32732 46396 32788
rect 46452 32732 46462 32788
rect 48402 32732 48412 32788
rect 48468 32732 50428 32788
rect 51202 32732 51212 32788
rect 51268 32732 60396 32788
rect 60452 32732 60462 32788
rect 6962 32620 6972 32676
rect 7028 32620 20860 32676
rect 20916 32620 20926 32676
rect 36092 32564 36148 32732
rect 44156 32676 44212 32732
rect 50372 32676 50428 32732
rect 37436 32620 38668 32676
rect 44156 32620 49812 32676
rect 50372 32620 58828 32676
rect 58884 32620 58894 32676
rect 37436 32564 37492 32620
rect 38612 32564 38668 32620
rect 9090 32508 9100 32564
rect 9156 32508 9884 32564
rect 9940 32508 16716 32564
rect 16772 32508 16782 32564
rect 17266 32508 17276 32564
rect 17332 32508 18396 32564
rect 18452 32508 23548 32564
rect 23604 32508 23614 32564
rect 25890 32508 25900 32564
rect 25956 32508 27132 32564
rect 27188 32508 28476 32564
rect 28532 32508 28542 32564
rect 36082 32508 36092 32564
rect 36148 32508 36158 32564
rect 37426 32508 37436 32564
rect 37492 32508 37502 32564
rect 38612 32508 45388 32564
rect 45444 32508 45454 32564
rect 45602 32508 45612 32564
rect 45668 32508 48076 32564
rect 48132 32508 48142 32564
rect 49756 32452 49812 32620
rect 53890 32508 53900 32564
rect 53956 32508 57708 32564
rect 57764 32508 57774 32564
rect 15026 32396 15036 32452
rect 15092 32396 16828 32452
rect 16884 32396 17612 32452
rect 17668 32396 17678 32452
rect 19506 32396 19516 32452
rect 19572 32396 21084 32452
rect 21140 32396 21150 32452
rect 21634 32396 21644 32452
rect 21700 32396 22316 32452
rect 22372 32396 23324 32452
rect 23380 32396 23772 32452
rect 23828 32396 24668 32452
rect 24724 32396 26684 32452
rect 26740 32396 26750 32452
rect 44706 32396 44716 32452
rect 44772 32396 45724 32452
rect 45780 32396 48524 32452
rect 48580 32396 48590 32452
rect 49746 32396 49756 32452
rect 49812 32396 49822 32452
rect 57586 32396 57596 32452
rect 57652 32396 57662 32452
rect 9202 32284 9212 32340
rect 9268 32284 10668 32340
rect 10724 32284 10734 32340
rect 38658 32284 38668 32340
rect 38724 32284 46172 32340
rect 46228 32284 46238 32340
rect 47058 32284 47068 32340
rect 47124 32284 50764 32340
rect 50820 32284 50830 32340
rect 57596 32228 57652 32396
rect 5170 32172 5180 32228
rect 5236 32172 17724 32228
rect 17780 32172 17790 32228
rect 45378 32172 45388 32228
rect 45444 32172 57652 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 20066 31948 20076 32004
rect 20132 31948 22988 32004
rect 23044 31948 23054 32004
rect 40450 31948 40460 32004
rect 40516 31948 53788 32004
rect 53844 31948 53854 32004
rect 4050 31836 4060 31892
rect 4116 31836 8428 31892
rect 9090 31836 9100 31892
rect 9156 31836 9436 31892
rect 9492 31836 9996 31892
rect 10052 31836 12012 31892
rect 12068 31836 12460 31892
rect 12516 31836 12526 31892
rect 13570 31836 13580 31892
rect 13636 31836 20188 31892
rect 22194 31836 22204 31892
rect 22260 31836 26628 31892
rect 28130 31836 28140 31892
rect 28196 31836 29372 31892
rect 29428 31836 29438 31892
rect 31154 31836 31164 31892
rect 31220 31836 33460 31892
rect 33730 31836 33740 31892
rect 33796 31836 36988 31892
rect 37044 31836 37054 31892
rect 48290 31836 48300 31892
rect 48356 31836 50428 31892
rect 53218 31836 53228 31892
rect 53284 31836 61516 31892
rect 61572 31836 61582 31892
rect 8372 31780 8428 31836
rect 20132 31780 20188 31836
rect 8372 31724 17724 31780
rect 17780 31724 17790 31780
rect 20132 31724 20972 31780
rect 21028 31724 21700 31780
rect 23986 31724 23996 31780
rect 24052 31724 24668 31780
rect 24724 31724 24734 31780
rect 21644 31668 21700 31724
rect 26572 31668 26628 31836
rect 33404 31780 33460 31836
rect 50372 31780 50428 31836
rect 29250 31724 29260 31780
rect 29316 31724 32172 31780
rect 32228 31724 32238 31780
rect 33394 31724 33404 31780
rect 33460 31724 33470 31780
rect 36530 31724 36540 31780
rect 36596 31724 47068 31780
rect 47124 31724 47134 31780
rect 50372 31724 57036 31780
rect 57092 31724 57102 31780
rect 3042 31612 3052 31668
rect 3108 31612 5292 31668
rect 5348 31612 5358 31668
rect 7074 31612 7084 31668
rect 7140 31612 20860 31668
rect 20916 31612 20926 31668
rect 21644 31612 24220 31668
rect 24276 31612 24286 31668
rect 26562 31612 26572 31668
rect 26628 31612 27804 31668
rect 27860 31612 31948 31668
rect 37314 31612 37324 31668
rect 37380 31612 38332 31668
rect 38388 31612 38398 31668
rect 41122 31612 41132 31668
rect 41188 31612 41916 31668
rect 41972 31612 41982 31668
rect 43148 31612 58492 31668
rect 58548 31612 58558 31668
rect 3938 31500 3948 31556
rect 4004 31500 9884 31556
rect 9940 31500 9950 31556
rect 18834 31500 18844 31556
rect 18900 31500 25004 31556
rect 25060 31500 25070 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 31892 31332 31948 31612
rect 43148 31556 43204 31612
rect 41682 31500 41692 31556
rect 41748 31500 43204 31556
rect 43362 31500 43372 31556
rect 43428 31500 43708 31556
rect 43764 31500 43774 31556
rect 47842 31500 47852 31556
rect 47908 31500 51548 31556
rect 51604 31500 51614 31556
rect 56242 31500 56252 31556
rect 56308 31500 65548 31556
rect 65604 31500 65614 31556
rect 57138 31388 57148 31444
rect 57204 31388 64316 31444
rect 64372 31388 64382 31444
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 31892 31276 37324 31332
rect 37380 31276 37772 31332
rect 37828 31276 45612 31332
rect 45668 31276 45678 31332
rect 56130 31276 56140 31332
rect 56196 31276 62524 31332
rect 62580 31276 62590 31332
rect 11330 31164 11340 31220
rect 11396 31164 13132 31220
rect 13188 31164 13198 31220
rect 25442 31164 25452 31220
rect 25508 31164 28588 31220
rect 28644 31164 28654 31220
rect 36082 31164 36092 31220
rect 36148 31164 39900 31220
rect 39956 31164 39966 31220
rect 41468 31164 50428 31220
rect 57026 31164 57036 31220
rect 57092 31164 60508 31220
rect 60564 31164 60574 31220
rect 2146 31052 2156 31108
rect 2212 31052 16940 31108
rect 16996 31052 17006 31108
rect 41468 30996 41524 31164
rect 50372 31108 50428 31164
rect 50372 31052 57484 31108
rect 57540 31052 57550 31108
rect 67200 30996 68000 31024
rect 12002 30940 12012 30996
rect 12068 30940 13244 30996
rect 13300 30940 14700 30996
rect 14756 30940 14766 30996
rect 20290 30940 20300 30996
rect 20356 30940 21308 30996
rect 21364 30940 21374 30996
rect 38322 30940 38332 30996
rect 38388 30940 39788 30996
rect 39844 30940 39854 30996
rect 41458 30940 41468 30996
rect 41524 30940 41534 30996
rect 49298 30940 49308 30996
rect 49364 30940 55972 30996
rect 60162 30940 60172 30996
rect 60228 30940 64988 30996
rect 65044 30940 65054 30996
rect 66098 30940 66108 30996
rect 66164 30940 68000 30996
rect 55916 30884 55972 30940
rect 67200 30912 68000 30940
rect 3154 30828 3164 30884
rect 3220 30828 9884 30884
rect 9940 30828 9950 30884
rect 16370 30828 16380 30884
rect 16436 30828 17836 30884
rect 17892 30828 17902 30884
rect 23538 30828 23548 30884
rect 23604 30828 26012 30884
rect 26068 30828 27132 30884
rect 27188 30828 29036 30884
rect 29092 30828 29102 30884
rect 32162 30828 32172 30884
rect 32228 30828 33180 30884
rect 33236 30828 33246 30884
rect 38658 30828 38668 30884
rect 38724 30828 52556 30884
rect 52612 30828 52622 30884
rect 55916 30828 61516 30884
rect 61572 30828 61582 30884
rect 2818 30716 2828 30772
rect 2884 30716 4396 30772
rect 4452 30716 4462 30772
rect 8194 30716 8204 30772
rect 8260 30716 14308 30772
rect 36642 30716 36652 30772
rect 36708 30716 38668 30772
rect 44482 30716 44492 30772
rect 44548 30716 46060 30772
rect 46116 30716 46126 30772
rect 52322 30716 52332 30772
rect 52388 30716 62412 30772
rect 62468 30716 62478 30772
rect 7074 30604 7084 30660
rect 7140 30604 13916 30660
rect 13972 30604 13982 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 14252 30548 14308 30716
rect 16706 30604 16716 30660
rect 16772 30604 18508 30660
rect 18564 30604 25900 30660
rect 25956 30604 25966 30660
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 38612 30548 38668 30716
rect 45154 30604 45164 30660
rect 45220 30604 57484 30660
rect 57540 30604 57550 30660
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 14252 30492 20188 30548
rect 20244 30492 20254 30548
rect 38612 30492 50876 30548
rect 50932 30492 50942 30548
rect 5058 30380 5068 30436
rect 5124 30380 23212 30436
rect 23268 30380 23278 30436
rect 24322 30380 24332 30436
rect 24388 30380 26348 30436
rect 26404 30380 26414 30436
rect 8978 30268 8988 30324
rect 9044 30268 10220 30324
rect 10276 30268 10286 30324
rect 14690 30268 14700 30324
rect 14756 30268 16828 30324
rect 16884 30268 16894 30324
rect 20290 30268 20300 30324
rect 20356 30268 20748 30324
rect 20804 30268 21308 30324
rect 21364 30268 23996 30324
rect 24052 30268 24062 30324
rect 33058 30268 33068 30324
rect 33124 30268 35644 30324
rect 35700 30268 35710 30324
rect 48066 30268 48076 30324
rect 48132 30268 48748 30324
rect 48804 30268 48814 30324
rect 52658 30268 52668 30324
rect 52724 30268 55468 30324
rect 55524 30268 55916 30324
rect 55972 30268 56476 30324
rect 56532 30268 56542 30324
rect 4050 30156 4060 30212
rect 4116 30156 11340 30212
rect 11396 30156 11406 30212
rect 12338 30156 12348 30212
rect 12404 30156 13692 30212
rect 13748 30156 13758 30212
rect 14018 30156 14028 30212
rect 14084 30156 15036 30212
rect 15092 30156 15102 30212
rect 18610 30156 18620 30212
rect 18676 30156 18686 30212
rect 21634 30156 21644 30212
rect 21700 30156 22316 30212
rect 22372 30156 22382 30212
rect 26226 30156 26236 30212
rect 26292 30156 27244 30212
rect 27300 30156 28252 30212
rect 28308 30156 29260 30212
rect 29316 30156 29326 30212
rect 33506 30156 33516 30212
rect 33572 30156 33582 30212
rect 38210 30156 38220 30212
rect 38276 30156 40684 30212
rect 40740 30156 40750 30212
rect 43586 30156 43596 30212
rect 43652 30156 46284 30212
rect 46340 30156 46732 30212
rect 46788 30156 52220 30212
rect 52276 30156 53900 30212
rect 53956 30156 53966 30212
rect 18620 30100 18676 30156
rect 3042 30044 3052 30100
rect 3108 30044 4508 30100
rect 4564 30044 4574 30100
rect 9874 30044 9884 30100
rect 9940 30044 18676 30100
rect 33516 30100 33572 30156
rect 33516 30044 41972 30100
rect 47730 30044 47740 30100
rect 47796 30044 50428 30100
rect 50484 30044 50494 30100
rect 51986 30044 51996 30100
rect 52052 30044 52780 30100
rect 52836 30044 52846 30100
rect 55570 30044 55580 30100
rect 55636 30044 61404 30100
rect 61460 30044 61470 30100
rect 41916 29988 41972 30044
rect 12338 29932 12348 29988
rect 12404 29932 14028 29988
rect 14084 29932 14094 29988
rect 25106 29932 25116 29988
rect 25172 29932 27580 29988
rect 27636 29932 27646 29988
rect 32162 29932 32172 29988
rect 32228 29932 33068 29988
rect 33124 29932 33134 29988
rect 40002 29932 40012 29988
rect 40068 29932 40908 29988
rect 40964 29932 40974 29988
rect 41916 29932 49644 29988
rect 49700 29932 49710 29988
rect 53218 29820 53228 29876
rect 53284 29820 61516 29876
rect 61572 29820 61582 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 3154 29708 3164 29764
rect 3220 29708 13244 29764
rect 13300 29708 13310 29764
rect 41682 29708 41692 29764
rect 41748 29708 43932 29764
rect 43988 29708 43998 29764
rect 8194 29596 8204 29652
rect 8260 29596 8428 29652
rect 16818 29596 16828 29652
rect 16884 29596 17500 29652
rect 17556 29596 17948 29652
rect 18004 29596 19068 29652
rect 19124 29596 20300 29652
rect 20356 29596 20366 29652
rect 32050 29596 32060 29652
rect 32116 29596 33740 29652
rect 33796 29596 33806 29652
rect 41570 29596 41580 29652
rect 41636 29596 41916 29652
rect 41972 29596 44156 29652
rect 44212 29596 44222 29652
rect 44706 29596 44716 29652
rect 44772 29596 46284 29652
rect 46340 29596 46844 29652
rect 46900 29596 46910 29652
rect 8372 29540 8428 29596
rect 6178 29484 6188 29540
rect 6244 29484 7868 29540
rect 7924 29484 7934 29540
rect 8372 29484 20188 29540
rect 29698 29484 29708 29540
rect 29764 29484 30492 29540
rect 30548 29484 30558 29540
rect 45378 29484 45388 29540
rect 45444 29484 57596 29540
rect 57652 29484 57662 29540
rect 20132 29428 20188 29484
rect 8082 29372 8092 29428
rect 8148 29372 8764 29428
rect 8820 29372 9100 29428
rect 9156 29372 9660 29428
rect 9716 29372 11564 29428
rect 11620 29372 11630 29428
rect 20132 29372 21644 29428
rect 21700 29372 21710 29428
rect 25330 29372 25340 29428
rect 25396 29372 26236 29428
rect 26292 29372 26302 29428
rect 31154 29372 31164 29428
rect 31220 29372 31948 29428
rect 32050 29372 32060 29428
rect 32116 29372 33292 29428
rect 33348 29372 33358 29428
rect 36194 29372 36204 29428
rect 36260 29372 38444 29428
rect 38500 29372 38892 29428
rect 38948 29372 38958 29428
rect 40674 29372 40684 29428
rect 40740 29372 42252 29428
rect 42308 29372 44156 29428
rect 44212 29372 44222 29428
rect 49298 29372 49308 29428
rect 49364 29372 50428 29428
rect 31892 29316 31948 29372
rect 50372 29316 50428 29372
rect 5282 29260 5292 29316
rect 5348 29260 15596 29316
rect 15652 29260 15662 29316
rect 19842 29260 19852 29316
rect 19908 29260 24556 29316
rect 24612 29260 24622 29316
rect 31892 29260 32620 29316
rect 32676 29260 33068 29316
rect 33124 29260 34636 29316
rect 34692 29260 37100 29316
rect 37156 29260 38556 29316
rect 38612 29260 38622 29316
rect 50372 29260 60396 29316
rect 60452 29260 60462 29316
rect 4162 29148 4172 29204
rect 4228 29148 4900 29204
rect 22530 29148 22540 29204
rect 22596 29148 28924 29204
rect 28980 29148 28990 29204
rect 45938 29148 45948 29204
rect 46004 29148 50428 29204
rect 52322 29148 52332 29204
rect 52388 29148 62188 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 4844 28980 4900 29148
rect 50372 29092 50428 29148
rect 6066 29036 6076 29092
rect 6132 29036 23548 29092
rect 23604 29036 23614 29092
rect 24434 29036 24444 29092
rect 24500 29036 25788 29092
rect 25844 29036 25854 29092
rect 50372 29036 58828 29092
rect 58884 29036 58894 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 62132 28980 62188 29148
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 4844 28924 17724 28980
rect 17780 28924 17790 28980
rect 48178 28924 48188 28980
rect 48244 28924 49756 28980
rect 49812 28924 51100 28980
rect 51156 28924 51166 28980
rect 62132 28924 62524 28980
rect 62580 28924 62590 28980
rect 4498 28812 4508 28868
rect 4564 28812 25788 28868
rect 25844 28812 25854 28868
rect 40562 28812 40572 28868
rect 40628 28812 45612 28868
rect 45668 28812 45678 28868
rect 48514 28812 48524 28868
rect 48580 28812 61404 28868
rect 61460 28812 61470 28868
rect 5170 28700 5180 28756
rect 5236 28700 6860 28756
rect 6916 28700 6926 28756
rect 12898 28700 12908 28756
rect 12964 28700 13916 28756
rect 13972 28700 15708 28756
rect 15764 28700 16380 28756
rect 16436 28700 16446 28756
rect 30706 28700 30716 28756
rect 30772 28700 33404 28756
rect 33460 28700 33964 28756
rect 34020 28700 36316 28756
rect 36372 28700 38332 28756
rect 38388 28700 38398 28756
rect 47730 28700 47740 28756
rect 47796 28700 51660 28756
rect 51716 28700 51726 28756
rect 51986 28700 51996 28756
rect 52052 28700 54348 28756
rect 54404 28700 54414 28756
rect 2034 28588 2044 28644
rect 2100 28588 5404 28644
rect 5460 28588 5470 28644
rect 6514 28588 6524 28644
rect 6580 28588 7196 28644
rect 7252 28588 7644 28644
rect 7700 28588 8764 28644
rect 8820 28588 9884 28644
rect 9940 28588 9950 28644
rect 12908 28532 12964 28700
rect 28242 28588 28252 28644
rect 28308 28588 29708 28644
rect 29764 28588 29774 28644
rect 45490 28588 45500 28644
rect 45556 28588 47908 28644
rect 49970 28588 49980 28644
rect 50036 28588 52668 28644
rect 52724 28588 52734 28644
rect 56018 28588 56028 28644
rect 56084 28588 59276 28644
rect 59332 28588 59342 28644
rect 47852 28532 47908 28588
rect 3042 28476 3052 28532
rect 3108 28476 4508 28532
rect 4564 28476 4574 28532
rect 11442 28476 11452 28532
rect 11508 28476 12964 28532
rect 28578 28476 28588 28532
rect 28644 28476 29932 28532
rect 29988 28476 31500 28532
rect 31556 28476 32396 28532
rect 32452 28476 32462 28532
rect 47852 28476 57596 28532
rect 57652 28476 57662 28532
rect 62514 28476 62524 28532
rect 62580 28476 62590 28532
rect 62524 28420 62580 28476
rect 6402 28364 6412 28420
rect 6468 28364 7420 28420
rect 7476 28364 7486 28420
rect 15026 28364 15036 28420
rect 15092 28364 16492 28420
rect 16548 28364 16558 28420
rect 30146 28364 30156 28420
rect 30212 28364 30940 28420
rect 30996 28364 31006 28420
rect 31714 28364 31724 28420
rect 31780 28364 33628 28420
rect 33684 28364 33694 28420
rect 37650 28364 37660 28420
rect 37716 28364 39900 28420
rect 39956 28364 39966 28420
rect 44370 28364 44380 28420
rect 44436 28364 50316 28420
rect 50372 28364 50382 28420
rect 51090 28364 51100 28420
rect 51156 28364 51996 28420
rect 52052 28364 52062 28420
rect 52434 28364 52444 28420
rect 52500 28364 62580 28420
rect 3938 28252 3948 28308
rect 4004 28252 10220 28308
rect 10276 28252 10286 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 24210 28140 24220 28196
rect 24276 28140 26572 28196
rect 26628 28140 26638 28196
rect 37538 28140 37548 28196
rect 37604 28140 38780 28196
rect 38836 28140 38846 28196
rect 4722 28028 4732 28084
rect 4788 28028 8428 28084
rect 8484 28028 8494 28084
rect 14018 28028 14028 28084
rect 14084 28028 17948 28084
rect 18004 28028 18014 28084
rect 26002 28028 26012 28084
rect 26068 28028 27244 28084
rect 27300 28028 27310 28084
rect 31826 28028 31836 28084
rect 31892 28028 32508 28084
rect 32564 28028 32574 28084
rect 49634 28028 49644 28084
rect 49700 28028 51212 28084
rect 51268 28028 53004 28084
rect 53060 28028 53070 28084
rect 54338 28028 54348 28084
rect 54404 28028 55300 28084
rect 55244 27972 55300 28028
rect 8306 27916 8316 27972
rect 8372 27916 10556 27972
rect 10612 27916 10622 27972
rect 12674 27916 12684 27972
rect 12740 27916 13692 27972
rect 13748 27916 13758 27972
rect 23762 27916 23772 27972
rect 23828 27916 29596 27972
rect 29652 27916 29662 27972
rect 39676 27916 40236 27972
rect 40292 27916 41916 27972
rect 41972 27916 41982 27972
rect 48402 27916 48412 27972
rect 48468 27916 50428 27972
rect 53106 27916 53116 27972
rect 53172 27916 54908 27972
rect 54964 27916 54974 27972
rect 55234 27916 55244 27972
rect 55300 27916 56028 27972
rect 56084 27916 56094 27972
rect 56242 27916 56252 27972
rect 56308 27916 61404 27972
rect 61460 27916 61470 27972
rect 39676 27860 39732 27916
rect 50372 27860 50428 27916
rect 4050 27804 4060 27860
rect 4116 27804 5964 27860
rect 6020 27804 6030 27860
rect 9874 27804 9884 27860
rect 9940 27804 10892 27860
rect 10948 27804 11452 27860
rect 11508 27804 11518 27860
rect 22306 27804 22316 27860
rect 22372 27804 23212 27860
rect 23268 27804 23660 27860
rect 23716 27804 24108 27860
rect 24164 27804 26236 27860
rect 26292 27804 26302 27860
rect 32386 27804 32396 27860
rect 32452 27804 33852 27860
rect 33908 27804 35084 27860
rect 35140 27804 35756 27860
rect 35812 27804 35822 27860
rect 39666 27804 39676 27860
rect 39732 27804 39742 27860
rect 44818 27804 44828 27860
rect 44884 27804 48748 27860
rect 48804 27804 49980 27860
rect 50036 27804 50046 27860
rect 50372 27804 58492 27860
rect 58548 27804 58558 27860
rect 16370 27692 16380 27748
rect 16436 27692 17612 27748
rect 17668 27692 18172 27748
rect 18228 27692 19740 27748
rect 19796 27692 19806 27748
rect 20738 27692 20748 27748
rect 20804 27692 24220 27748
rect 24276 27692 24286 27748
rect 24658 27692 24668 27748
rect 24724 27692 25228 27748
rect 25284 27692 25294 27748
rect 40002 27692 40012 27748
rect 40068 27692 41468 27748
rect 41524 27692 41534 27748
rect 47842 27692 47852 27748
rect 47908 27692 49196 27748
rect 49252 27692 49262 27748
rect 49522 27692 49532 27748
rect 49588 27692 49756 27748
rect 49812 27692 49822 27748
rect 53218 27692 53228 27748
rect 53284 27692 60396 27748
rect 60452 27692 60462 27748
rect 3042 27580 3052 27636
rect 3108 27580 8092 27636
rect 8148 27580 8158 27636
rect 8372 27580 11900 27636
rect 11956 27580 11966 27636
rect 23090 27580 23100 27636
rect 23156 27580 27468 27636
rect 27524 27580 27534 27636
rect 55570 27580 55580 27636
rect 55636 27580 59276 27636
rect 59332 27580 59342 27636
rect 8372 27524 8428 27580
rect 6626 27468 6636 27524
rect 6692 27468 8428 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 50642 27356 50652 27412
rect 50708 27356 60284 27412
rect 60340 27356 60350 27412
rect 3490 27244 3500 27300
rect 3556 27244 11116 27300
rect 11172 27244 11182 27300
rect 20290 27244 20300 27300
rect 20356 27244 21308 27300
rect 21364 27244 21374 27300
rect 43922 27244 43932 27300
rect 43988 27244 53564 27300
rect 53620 27244 53630 27300
rect 4050 27132 4060 27188
rect 4116 27132 10108 27188
rect 10164 27132 10174 27188
rect 22428 27132 24668 27188
rect 24724 27132 24734 27188
rect 31378 27132 31388 27188
rect 31444 27132 33964 27188
rect 34020 27132 34030 27188
rect 45388 27132 57484 27188
rect 57540 27132 57550 27188
rect 22428 27076 22484 27132
rect 45388 27076 45444 27132
rect 13794 27020 13804 27076
rect 13860 27020 14812 27076
rect 14868 27020 15932 27076
rect 15988 27020 15998 27076
rect 19730 27020 19740 27076
rect 19796 27020 21532 27076
rect 21588 27020 22428 27076
rect 22484 27020 22494 27076
rect 23650 27020 23660 27076
rect 23716 27020 28028 27076
rect 28084 27020 28094 27076
rect 37090 27020 37100 27076
rect 37156 27020 38556 27076
rect 38612 27020 40684 27076
rect 40740 27020 40750 27076
rect 41346 27020 41356 27076
rect 41412 27020 44156 27076
rect 44212 27020 44222 27076
rect 45378 27020 45388 27076
rect 45444 27020 45454 27076
rect 49074 27020 49084 27076
rect 49140 27020 50764 27076
rect 50820 27020 50830 27076
rect 53218 27020 53228 27076
rect 53284 27020 61516 27076
rect 61572 27020 61582 27076
rect 5730 26908 5740 26964
rect 5796 26908 7196 26964
rect 7252 26908 7262 26964
rect 14690 26908 14700 26964
rect 14756 26908 15372 26964
rect 15428 26908 16380 26964
rect 16436 26908 16446 26964
rect 20066 26908 20076 26964
rect 20132 26908 23884 26964
rect 23940 26908 23950 26964
rect 34514 26908 34524 26964
rect 34580 26908 36092 26964
rect 36148 26908 36158 26964
rect 7196 26852 7252 26908
rect 7196 26796 8316 26852
rect 8372 26796 8382 26852
rect 11554 26796 11564 26852
rect 11620 26796 15596 26852
rect 15652 26796 15662 26852
rect 19954 26796 19964 26852
rect 20020 26796 21588 26852
rect 26674 26796 26684 26852
rect 26740 26796 28364 26852
rect 28420 26796 28430 26852
rect 32722 26796 32732 26852
rect 32788 26796 33628 26852
rect 33684 26796 33694 26852
rect 45042 26796 45052 26852
rect 45108 26796 58492 26852
rect 58548 26796 58558 26852
rect 21532 26740 21588 26796
rect 21522 26684 21532 26740
rect 21588 26684 21598 26740
rect 28578 26684 28588 26740
rect 28644 26684 29372 26740
rect 29428 26684 29438 26740
rect 34738 26684 34748 26740
rect 34804 26684 36876 26740
rect 36932 26684 36942 26740
rect 56354 26684 56364 26740
rect 56420 26684 61404 26740
rect 61460 26684 61470 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 3938 26460 3948 26516
rect 4004 26460 8652 26516
rect 8708 26460 8718 26516
rect 11666 26460 11676 26516
rect 11732 26460 13580 26516
rect 13636 26460 16380 26516
rect 16436 26460 16446 26516
rect 18274 26460 18284 26516
rect 18340 26460 20860 26516
rect 20916 26460 20926 26516
rect 28242 26460 28252 26516
rect 28308 26460 29372 26516
rect 29428 26460 29438 26516
rect 33730 26460 33740 26516
rect 33796 26460 34748 26516
rect 34804 26460 34814 26516
rect 44482 26460 44492 26516
rect 44548 26460 49084 26516
rect 49140 26460 49150 26516
rect 53666 26460 53676 26516
rect 53732 26460 55468 26516
rect 55412 26404 55468 26460
rect 21746 26348 21756 26404
rect 21812 26348 23996 26404
rect 24052 26348 24062 26404
rect 50306 26348 50316 26404
rect 50372 26348 54572 26404
rect 54628 26348 54638 26404
rect 55412 26348 58828 26404
rect 58884 26348 58894 26404
rect 1810 26236 1820 26292
rect 1876 26236 4508 26292
rect 4564 26236 5404 26292
rect 5460 26236 5470 26292
rect 5954 26236 5964 26292
rect 6020 26236 6524 26292
rect 6580 26236 9772 26292
rect 9828 26236 10892 26292
rect 10948 26236 10958 26292
rect 19506 26236 19516 26292
rect 19572 26236 21644 26292
rect 21700 26236 21710 26292
rect 25218 26236 25228 26292
rect 25284 26236 25676 26292
rect 25732 26236 25742 26292
rect 45490 26124 45500 26180
rect 45556 26124 57596 26180
rect 57652 26124 57662 26180
rect 2930 26012 2940 26068
rect 2996 26012 9100 26068
rect 9156 26012 9166 26068
rect 15474 26012 15484 26068
rect 15540 26012 17276 26068
rect 17332 26012 17342 26068
rect 44034 26012 44044 26068
rect 44100 26012 46956 26068
rect 47012 26012 48748 26068
rect 48804 26012 48814 26068
rect 52322 26012 52332 26068
rect 52388 26012 62524 26068
rect 62580 26012 62590 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 16370 25788 16380 25844
rect 16436 25788 17276 25844
rect 17332 25788 17342 25844
rect 38434 25788 38444 25844
rect 38500 25788 39900 25844
rect 39956 25788 39966 25844
rect 7522 25676 7532 25732
rect 7588 25676 9324 25732
rect 9380 25676 9390 25732
rect 18050 25676 18060 25732
rect 18116 25676 19404 25732
rect 19460 25676 19470 25732
rect 29474 25676 29484 25732
rect 29540 25676 30380 25732
rect 30436 25676 30446 25732
rect 45378 25676 45388 25732
rect 45444 25676 49196 25732
rect 49252 25676 49262 25732
rect 7746 25564 7756 25620
rect 7812 25564 12684 25620
rect 12740 25564 12750 25620
rect 29698 25564 29708 25620
rect 29764 25564 30828 25620
rect 30884 25564 30894 25620
rect 39554 25564 39564 25620
rect 39620 25564 41916 25620
rect 41972 25564 42700 25620
rect 42756 25564 43148 25620
rect 43204 25564 44044 25620
rect 44100 25564 44110 25620
rect 48402 25564 48412 25620
rect 48468 25564 58716 25620
rect 58772 25564 58782 25620
rect 8978 25452 8988 25508
rect 9044 25452 10220 25508
rect 10276 25452 11452 25508
rect 11508 25452 11518 25508
rect 20178 25452 20188 25508
rect 20244 25452 20636 25508
rect 20692 25452 20702 25508
rect 29250 25452 29260 25508
rect 29316 25452 31388 25508
rect 31444 25452 31454 25508
rect 36418 25452 36428 25508
rect 36484 25452 38444 25508
rect 38500 25452 38510 25508
rect 48962 25452 48972 25508
rect 49028 25452 57876 25508
rect 58930 25452 58940 25508
rect 58996 25452 59006 25508
rect 57820 25396 57876 25452
rect 58940 25396 58996 25452
rect 8306 25340 8316 25396
rect 8372 25340 9436 25396
rect 9492 25340 9502 25396
rect 19282 25340 19292 25396
rect 19348 25340 21420 25396
rect 21476 25340 21486 25396
rect 28130 25340 28140 25396
rect 28196 25340 30380 25396
rect 30436 25340 30446 25396
rect 41570 25340 41580 25396
rect 41636 25340 42364 25396
rect 42420 25340 42430 25396
rect 49298 25340 49308 25396
rect 49364 25340 57596 25396
rect 57652 25340 57662 25396
rect 57820 25340 58996 25396
rect 3826 25228 3836 25284
rect 3892 25228 9548 25284
rect 9604 25228 9614 25284
rect 9762 25228 9772 25284
rect 9828 25228 15820 25284
rect 15876 25228 15886 25284
rect 17378 25228 17388 25284
rect 17444 25228 20300 25284
rect 20356 25228 20748 25284
rect 20804 25228 20814 25284
rect 25106 25228 25116 25284
rect 25172 25228 27468 25284
rect 27524 25228 29148 25284
rect 29204 25228 30044 25284
rect 30100 25228 30940 25284
rect 30996 25228 31006 25284
rect 37314 25228 37324 25284
rect 37380 25228 39004 25284
rect 39060 25228 39070 25284
rect 45602 25228 45612 25284
rect 45668 25228 47628 25284
rect 47684 25228 47694 25284
rect 55906 25228 55916 25284
rect 55972 25228 59612 25284
rect 59668 25228 59678 25284
rect 19180 25172 19236 25228
rect 19170 25116 19180 25172
rect 19236 25116 19246 25172
rect 19618 25116 19628 25172
rect 19684 25116 19694 25172
rect 51762 25116 51772 25172
rect 51828 25116 55132 25172
rect 55188 25116 55198 25172
rect 19628 25060 19684 25116
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 4050 25004 4060 25060
rect 4116 25004 5068 25060
rect 5124 25004 5134 25060
rect 17938 25004 17948 25060
rect 18004 25004 19684 25060
rect 40898 25004 40908 25060
rect 40964 25004 43148 25060
rect 43204 25004 43214 25060
rect 0 24948 800 24976
rect 19628 24948 19684 25004
rect 0 24892 1708 24948
rect 1764 24892 1774 24948
rect 4722 24892 4732 24948
rect 4788 24892 6188 24948
rect 6244 24892 6254 24948
rect 19628 24892 20748 24948
rect 20804 24892 21308 24948
rect 21364 24892 21374 24948
rect 24322 24892 24332 24948
rect 24388 24892 27244 24948
rect 27300 24892 27310 24948
rect 41122 24892 41132 24948
rect 41188 24892 42140 24948
rect 42196 24892 42206 24948
rect 47730 24892 47740 24948
rect 47796 24892 50204 24948
rect 50260 24892 50270 24948
rect 53442 24892 53452 24948
rect 53508 24892 60396 24948
rect 60452 24892 60462 24948
rect 0 24864 800 24892
rect 21308 24836 21364 24892
rect 2706 24780 2716 24836
rect 2772 24780 12684 24836
rect 12740 24780 12750 24836
rect 19170 24780 19180 24836
rect 19236 24780 19628 24836
rect 19684 24780 19694 24836
rect 21308 24780 24668 24836
rect 24724 24780 24734 24836
rect 31378 24780 31388 24836
rect 31444 24780 34076 24836
rect 34132 24780 34142 24836
rect 49186 24780 49196 24836
rect 49252 24780 50876 24836
rect 50932 24780 51996 24836
rect 52052 24780 52062 24836
rect 56466 24780 56476 24836
rect 56532 24780 58828 24836
rect 58884 24780 58894 24836
rect 13346 24668 13356 24724
rect 13412 24668 15148 24724
rect 17602 24668 17612 24724
rect 17668 24668 17948 24724
rect 18004 24668 18014 24724
rect 23314 24668 23324 24724
rect 23380 24668 24556 24724
rect 24612 24668 24622 24724
rect 25218 24668 25228 24724
rect 25284 24668 26124 24724
rect 26180 24668 30940 24724
rect 30996 24668 31006 24724
rect 48850 24668 48860 24724
rect 48916 24668 51212 24724
rect 51268 24668 52444 24724
rect 52500 24668 52892 24724
rect 52948 24668 52958 24724
rect 8306 24556 8316 24612
rect 8372 24556 10668 24612
rect 10724 24556 10734 24612
rect 15092 24500 15148 24668
rect 28914 24556 28924 24612
rect 28980 24556 30044 24612
rect 30100 24556 30110 24612
rect 39106 24556 39116 24612
rect 39172 24556 40348 24612
rect 40404 24556 41692 24612
rect 41748 24556 41758 24612
rect 42354 24556 42364 24612
rect 42420 24556 49420 24612
rect 49476 24556 49486 24612
rect 15092 24444 15708 24500
rect 15764 24444 16828 24500
rect 16884 24444 16894 24500
rect 18834 24444 18844 24500
rect 18900 24444 19852 24500
rect 19908 24444 19918 24500
rect 54898 24444 54908 24500
rect 54964 24444 61404 24500
rect 61460 24444 61470 24500
rect 40674 24332 40684 24388
rect 40740 24332 41132 24388
rect 41188 24332 41198 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 28690 24220 28700 24276
rect 28756 24220 29708 24276
rect 29764 24220 29774 24276
rect 37426 24220 37436 24276
rect 37492 24220 40124 24276
rect 40180 24220 40190 24276
rect 45266 24220 45276 24276
rect 45332 24220 57708 24276
rect 57764 24220 57774 24276
rect 43698 24108 43708 24164
rect 43764 24108 46508 24164
rect 46564 24108 46574 24164
rect 5058 23996 5068 24052
rect 5124 23996 5404 24052
rect 5460 23996 5470 24052
rect 16370 23996 16380 24052
rect 16436 23996 19068 24052
rect 19124 23996 19134 24052
rect 27906 23996 27916 24052
rect 27972 23996 29148 24052
rect 29204 23996 29214 24052
rect 42914 23996 42924 24052
rect 42980 23996 50092 24052
rect 50148 23996 50158 24052
rect 55458 23996 55468 24052
rect 55524 23996 55916 24052
rect 55972 23996 58604 24052
rect 58660 23996 59500 24052
rect 59556 23996 59566 24052
rect 10882 23884 10892 23940
rect 10948 23884 11900 23940
rect 11956 23884 12684 23940
rect 12740 23884 12908 23940
rect 12964 23884 12974 23940
rect 20290 23884 20300 23940
rect 20356 23884 21196 23940
rect 21252 23884 23324 23940
rect 23380 23884 23390 23940
rect 34290 23884 34300 23940
rect 34356 23884 35084 23940
rect 35140 23884 36428 23940
rect 36484 23884 36494 23940
rect 37090 23884 37100 23940
rect 37156 23884 38724 23940
rect 53106 23884 53116 23940
rect 53172 23884 53900 23940
rect 53956 23884 56476 23940
rect 56532 23884 56542 23940
rect 38668 23828 38724 23884
rect 3042 23772 3052 23828
rect 3108 23772 6748 23828
rect 6804 23772 6814 23828
rect 38668 23772 40348 23828
rect 40404 23772 40796 23828
rect 40852 23772 41020 23828
rect 41076 23772 41086 23828
rect 46050 23772 46060 23828
rect 46116 23772 51100 23828
rect 51156 23772 51166 23828
rect 51762 23772 51772 23828
rect 51828 23772 58268 23828
rect 58324 23772 58334 23828
rect 10210 23660 10220 23716
rect 10276 23660 12572 23716
rect 12628 23660 12638 23716
rect 24322 23660 24332 23716
rect 24388 23660 24892 23716
rect 24948 23660 24958 23716
rect 32050 23660 32060 23716
rect 32116 23660 34076 23716
rect 34132 23660 34142 23716
rect 38994 23660 39004 23716
rect 39060 23660 41580 23716
rect 41636 23660 41646 23716
rect 3042 23548 3052 23604
rect 3108 23548 5292 23604
rect 5348 23548 5358 23604
rect 9314 23548 9324 23604
rect 9380 23548 12124 23604
rect 12180 23548 12908 23604
rect 12964 23548 13356 23604
rect 13412 23548 13422 23604
rect 29586 23548 29596 23604
rect 29652 23548 30604 23604
rect 30660 23548 30670 23604
rect 32946 23548 32956 23604
rect 33012 23548 34412 23604
rect 34468 23548 34478 23604
rect 36082 23548 36092 23604
rect 36148 23548 37100 23604
rect 37156 23548 37166 23604
rect 40450 23548 40460 23604
rect 40516 23548 42700 23604
rect 42756 23548 42766 23604
rect 47954 23548 47964 23604
rect 48020 23548 49756 23604
rect 49812 23548 49822 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 44370 23436 44380 23492
rect 44436 23436 46060 23492
rect 46116 23436 46126 23492
rect 10098 23324 10108 23380
rect 10164 23324 10892 23380
rect 10948 23324 10958 23380
rect 32386 23324 32396 23380
rect 32452 23324 33740 23380
rect 33796 23324 33806 23380
rect 48850 23324 48860 23380
rect 48916 23324 49644 23380
rect 49700 23324 49710 23380
rect 32050 23212 32060 23268
rect 32116 23212 33068 23268
rect 33124 23212 33134 23268
rect 56242 23212 56252 23268
rect 56308 23212 58828 23268
rect 58884 23212 58894 23268
rect 4162 23100 4172 23156
rect 4228 23100 5964 23156
rect 6020 23100 6030 23156
rect 19506 23100 19516 23156
rect 19572 23100 20300 23156
rect 20356 23100 20366 23156
rect 24770 23100 24780 23156
rect 24836 23100 25116 23156
rect 25172 23100 25182 23156
rect 27906 23100 27916 23156
rect 27972 23100 29148 23156
rect 29204 23100 29932 23156
rect 29988 23100 29998 23156
rect 35756 23100 38108 23156
rect 38164 23100 38444 23156
rect 38500 23100 38892 23156
rect 38948 23100 39564 23156
rect 39620 23100 39630 23156
rect 46050 23100 46060 23156
rect 46116 23100 46956 23156
rect 47012 23100 48860 23156
rect 48916 23100 48926 23156
rect 49298 23100 49308 23156
rect 49364 23100 50204 23156
rect 50260 23100 50270 23156
rect 35756 23044 35812 23100
rect 30482 22988 30492 23044
rect 30548 22988 33292 23044
rect 33348 22988 33964 23044
rect 34020 22988 35756 23044
rect 35812 22988 35822 23044
rect 37324 22932 37380 23100
rect 37650 22988 37660 23044
rect 37716 22988 39788 23044
rect 39844 22988 39854 23044
rect 51874 22988 51884 23044
rect 51940 22988 57596 23044
rect 57652 22988 57662 23044
rect 10882 22876 10892 22932
rect 10948 22876 13244 22932
rect 13300 22876 13310 22932
rect 37314 22876 37324 22932
rect 37380 22876 37390 22932
rect 52322 22876 52332 22932
rect 52388 22876 58492 22932
rect 58548 22876 58558 22932
rect 29138 22764 29148 22820
rect 29204 22764 30156 22820
rect 30212 22764 30222 22820
rect 41318 22764 41356 22820
rect 41412 22764 41422 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 44790 22652 44828 22708
rect 44884 22652 44894 22708
rect 45826 22652 45836 22708
rect 45892 22652 53676 22708
rect 53732 22652 53742 22708
rect 22082 22540 22092 22596
rect 22148 22540 22764 22596
rect 22820 22540 22830 22596
rect 27346 22540 27356 22596
rect 27412 22540 29148 22596
rect 29204 22540 29214 22596
rect 40562 22540 40572 22596
rect 40628 22540 42924 22596
rect 42980 22540 42990 22596
rect 48290 22540 48300 22596
rect 48356 22540 50428 22596
rect 50484 22540 50494 22596
rect 54338 22540 54348 22596
rect 54404 22540 55580 22596
rect 55636 22540 55646 22596
rect 25330 22428 25340 22484
rect 25396 22428 26460 22484
rect 26516 22428 26526 22484
rect 50372 22428 57484 22484
rect 57540 22428 57550 22484
rect 50372 22372 50428 22428
rect 13570 22316 13580 22372
rect 13636 22316 15820 22372
rect 15876 22316 17164 22372
rect 17220 22316 17500 22372
rect 17556 22316 20748 22372
rect 20804 22316 20814 22372
rect 22754 22316 22764 22372
rect 22820 22316 25228 22372
rect 25284 22316 26908 22372
rect 26964 22316 26974 22372
rect 33058 22316 33068 22372
rect 33124 22316 34300 22372
rect 34356 22316 34972 22372
rect 35028 22316 35038 22372
rect 49074 22316 49084 22372
rect 49140 22316 50428 22372
rect 4050 22204 4060 22260
rect 4116 22204 5852 22260
rect 5908 22204 5918 22260
rect 28578 22204 28588 22260
rect 28644 22204 30156 22260
rect 30212 22204 30492 22260
rect 30548 22204 30558 22260
rect 43922 22204 43932 22260
rect 43988 22204 46284 22260
rect 46340 22204 46350 22260
rect 48402 22204 48412 22260
rect 48468 22204 53900 22260
rect 53956 22204 53966 22260
rect 55682 22204 55692 22260
rect 55748 22204 59612 22260
rect 59668 22204 59678 22260
rect 9202 22092 9212 22148
rect 9268 22092 10780 22148
rect 10836 22092 10846 22148
rect 16370 22092 16380 22148
rect 16436 22092 17052 22148
rect 17108 22092 17118 22148
rect 23986 22092 23996 22148
rect 24052 22092 25116 22148
rect 25172 22092 25182 22148
rect 32274 22092 32284 22148
rect 32340 22092 35532 22148
rect 35588 22092 35598 22148
rect 44930 22092 44940 22148
rect 44996 22092 48860 22148
rect 48916 22092 48926 22148
rect 49634 22092 49644 22148
rect 49700 22092 51884 22148
rect 51940 22092 51950 22148
rect 7858 21980 7868 22036
rect 7924 21980 9772 22036
rect 9828 21980 9838 22036
rect 12562 21980 12572 22036
rect 12628 21980 17612 22036
rect 17668 21980 17678 22036
rect 25778 21980 25788 22036
rect 25844 21980 27356 22036
rect 27412 21980 27422 22036
rect 45378 21980 45388 22036
rect 45444 21980 45454 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 7634 21868 7644 21924
rect 7700 21868 8652 21924
rect 8708 21868 8718 21924
rect 11890 21868 11900 21924
rect 11956 21868 13916 21924
rect 13972 21868 13982 21924
rect 25330 21868 25340 21924
rect 25396 21868 27468 21924
rect 27524 21868 27534 21924
rect 34626 21868 34636 21924
rect 34692 21868 35756 21924
rect 35812 21868 35822 21924
rect 36530 21868 36540 21924
rect 36596 21868 38220 21924
rect 38276 21868 38286 21924
rect 45388 21812 45444 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 45602 21868 45612 21924
rect 45668 21868 46060 21924
rect 46116 21868 46126 21924
rect 4834 21756 4844 21812
rect 4900 21756 5964 21812
rect 6020 21756 6030 21812
rect 9202 21756 9212 21812
rect 9268 21756 9278 21812
rect 9426 21756 9436 21812
rect 9492 21756 10556 21812
rect 10612 21756 10622 21812
rect 12450 21756 12460 21812
rect 12516 21756 13804 21812
rect 13860 21756 13870 21812
rect 17266 21756 17276 21812
rect 17332 21756 19068 21812
rect 19124 21756 19134 21812
rect 32386 21756 32396 21812
rect 32452 21756 34524 21812
rect 34580 21756 34590 21812
rect 34850 21756 34860 21812
rect 34916 21756 38444 21812
rect 38500 21756 38510 21812
rect 45388 21756 48524 21812
rect 48580 21756 48590 21812
rect 9212 21700 9268 21756
rect 5628 21644 7756 21700
rect 7812 21644 9268 21700
rect 10994 21644 11004 21700
rect 11060 21644 16268 21700
rect 16324 21644 16334 21700
rect 24658 21644 24668 21700
rect 24724 21644 25788 21700
rect 25844 21644 25854 21700
rect 35186 21644 35196 21700
rect 35252 21644 35868 21700
rect 35924 21644 35934 21700
rect 41346 21644 41356 21700
rect 41412 21644 49644 21700
rect 49700 21644 49710 21700
rect 52882 21644 52892 21700
rect 52948 21644 54012 21700
rect 54068 21644 54078 21700
rect 56130 21644 56140 21700
rect 56196 21644 58828 21700
rect 58884 21644 58894 21700
rect 5628 21588 5684 21644
rect 5618 21532 5628 21588
rect 5684 21532 5694 21588
rect 5852 21532 8988 21588
rect 9044 21532 9054 21588
rect 23874 21532 23884 21588
rect 23940 21532 27580 21588
rect 27636 21532 27646 21588
rect 29474 21532 29484 21588
rect 29540 21532 31612 21588
rect 31668 21532 31678 21588
rect 32386 21532 32396 21588
rect 32452 21532 33404 21588
rect 33460 21532 33470 21588
rect 39442 21532 39452 21588
rect 39508 21532 39788 21588
rect 39844 21532 41020 21588
rect 41076 21532 41086 21588
rect 42242 21532 42252 21588
rect 42308 21532 45724 21588
rect 45780 21532 45790 21588
rect 45938 21532 45948 21588
rect 46004 21532 49756 21588
rect 49812 21532 49822 21588
rect 5852 21476 5908 21532
rect 3154 21420 3164 21476
rect 3220 21420 5908 21476
rect 8194 21420 8204 21476
rect 8260 21420 9660 21476
rect 9716 21420 9726 21476
rect 24770 21420 24780 21476
rect 24836 21420 25900 21476
rect 25956 21420 25966 21476
rect 32498 21420 32508 21476
rect 32564 21420 34076 21476
rect 34132 21420 34142 21476
rect 42578 21420 42588 21476
rect 42644 21420 46060 21476
rect 46116 21420 46126 21476
rect 53218 21420 53228 21476
rect 53284 21420 57596 21476
rect 57652 21420 57662 21476
rect 33394 21308 33404 21364
rect 33460 21308 35756 21364
rect 35812 21308 35822 21364
rect 15586 21196 15596 21252
rect 15652 21196 16156 21252
rect 16212 21196 16222 21252
rect 49522 21196 49532 21252
rect 49588 21196 53676 21252
rect 53732 21196 53742 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 9874 21084 9884 21140
rect 9940 21084 13020 21140
rect 13076 21084 13086 21140
rect 48402 20972 48412 21028
rect 48468 20972 54796 21028
rect 54852 20972 54862 21028
rect 12674 20860 12684 20916
rect 12740 20860 13468 20916
rect 13524 20860 13534 20916
rect 15250 20860 15260 20916
rect 15316 20860 16716 20916
rect 16772 20860 16782 20916
rect 19282 20860 19292 20916
rect 19348 20860 19740 20916
rect 19796 20860 20412 20916
rect 20468 20860 21756 20916
rect 21812 20860 21822 20916
rect 35970 20860 35980 20916
rect 36036 20860 36988 20916
rect 37044 20860 37054 20916
rect 7970 20748 7980 20804
rect 8036 20748 8428 20804
rect 8484 20748 8494 20804
rect 15698 20748 15708 20804
rect 15764 20748 16380 20804
rect 16436 20748 16446 20804
rect 11778 20636 11788 20692
rect 11844 20636 13692 20692
rect 13748 20636 13758 20692
rect 37986 20636 37996 20692
rect 38052 20636 38892 20692
rect 38948 20636 38958 20692
rect 52210 20636 52220 20692
rect 52276 20636 54684 20692
rect 54740 20636 54750 20692
rect 16370 20524 16380 20580
rect 16436 20524 16828 20580
rect 16884 20524 16894 20580
rect 18162 20524 18172 20580
rect 18228 20524 18732 20580
rect 18788 20524 18798 20580
rect 32610 20412 32620 20468
rect 32676 20412 33740 20468
rect 33796 20412 33806 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 9202 20300 9212 20356
rect 9268 20300 9660 20356
rect 9716 20300 9726 20356
rect 11732 20300 12684 20356
rect 12740 20300 12750 20356
rect 17826 20300 17836 20356
rect 17892 20300 18620 20356
rect 18676 20300 18686 20356
rect 28802 20300 28812 20356
rect 28868 20300 31276 20356
rect 31332 20300 31342 20356
rect 40002 20300 40012 20356
rect 40068 20300 41804 20356
rect 41860 20300 41870 20356
rect 5170 20188 5180 20244
rect 5236 20188 5572 20244
rect 5516 20020 5572 20188
rect 5516 19964 6636 20020
rect 6692 19964 6702 20020
rect 11732 19908 11788 20300
rect 18050 20188 18060 20244
rect 18116 20188 18508 20244
rect 18564 20188 18574 20244
rect 23202 20188 23212 20244
rect 23268 20188 24220 20244
rect 24276 20188 24286 20244
rect 29586 20188 29596 20244
rect 29652 20188 31164 20244
rect 31220 20188 31230 20244
rect 36642 20188 36652 20244
rect 36708 20188 37996 20244
rect 38052 20188 38062 20244
rect 41010 20188 41020 20244
rect 41076 20188 42364 20244
rect 42420 20188 42430 20244
rect 48626 20188 48636 20244
rect 48692 20188 49140 20244
rect 49084 20132 49140 20188
rect 17490 20076 17500 20132
rect 17556 20076 19068 20132
rect 19124 20076 20636 20132
rect 20692 20076 20702 20132
rect 45042 20076 45052 20132
rect 45108 20076 46732 20132
rect 46788 20076 46798 20132
rect 47058 20076 47068 20132
rect 47124 20076 47516 20132
rect 47572 20076 47582 20132
rect 48178 20076 48188 20132
rect 48244 20076 48860 20132
rect 48916 20076 48926 20132
rect 49084 20076 50764 20132
rect 50820 20076 50830 20132
rect 55412 20076 55916 20132
rect 55972 20076 55982 20132
rect 55412 20020 55468 20076
rect 16818 19964 16828 20020
rect 16884 19964 17836 20020
rect 17892 19964 18844 20020
rect 18900 19964 19292 20020
rect 19348 19964 19358 20020
rect 23538 19964 23548 20020
rect 23604 19964 24668 20020
rect 24724 19964 25340 20020
rect 25396 19964 25406 20020
rect 44706 19964 44716 20020
rect 44772 19964 48636 20020
rect 48692 19964 48702 20020
rect 51426 19964 51436 20020
rect 51492 19964 54460 20020
rect 54516 19964 55468 20020
rect 7970 19852 7980 19908
rect 8036 19852 8988 19908
rect 9044 19852 11788 19908
rect 15092 19852 15484 19908
rect 15540 19852 17388 19908
rect 17444 19852 17454 19908
rect 45378 19852 45388 19908
rect 45444 19852 52556 19908
rect 52612 19852 52622 19908
rect 15092 19684 15148 19852
rect 44818 19740 44828 19796
rect 44884 19740 49644 19796
rect 49700 19740 49710 19796
rect 14914 19628 14924 19684
rect 14980 19628 15148 19684
rect 43698 19628 43708 19684
rect 43764 19628 44268 19684
rect 44324 19628 46396 19684
rect 46452 19628 46462 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 18498 19516 18508 19572
rect 18564 19516 19516 19572
rect 19572 19516 19582 19572
rect 2258 19292 2268 19348
rect 2324 19292 8316 19348
rect 8372 19292 8382 19348
rect 16818 19292 16828 19348
rect 16884 19292 17724 19348
rect 17780 19292 17790 19348
rect 20626 19292 20636 19348
rect 20692 19292 21420 19348
rect 21476 19292 22540 19348
rect 22596 19292 23212 19348
rect 23268 19292 23884 19348
rect 23940 19292 26572 19348
rect 26628 19292 26638 19348
rect 42354 19292 42364 19348
rect 42420 19292 44380 19348
rect 44436 19292 45052 19348
rect 45108 19292 45118 19348
rect 19506 19180 19516 19236
rect 19572 19180 22092 19236
rect 22148 19180 22158 19236
rect 23762 19068 23772 19124
rect 23828 19068 25452 19124
rect 25508 19068 25518 19124
rect 40786 19068 40796 19124
rect 40852 19068 42588 19124
rect 42644 19068 42654 19124
rect 44482 19068 44492 19124
rect 44548 19068 47068 19124
rect 47124 19068 47134 19124
rect 52658 19068 52668 19124
rect 52724 19068 55020 19124
rect 55076 19068 55086 19124
rect 17490 18956 17500 19012
rect 17556 18956 20300 19012
rect 20356 18956 20366 19012
rect 41234 18956 41244 19012
rect 41300 18956 45836 19012
rect 45892 18956 45902 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 44594 18620 44604 18676
rect 44660 18620 44670 18676
rect 19058 18508 19068 18564
rect 19124 18508 23996 18564
rect 24052 18508 24062 18564
rect 28466 18508 28476 18564
rect 28532 18508 30156 18564
rect 30212 18508 30222 18564
rect 34626 18508 34636 18564
rect 34692 18508 35756 18564
rect 35812 18508 35822 18564
rect 44604 18452 44660 18620
rect 46834 18508 46844 18564
rect 46900 18508 47852 18564
rect 47908 18508 47918 18564
rect 7186 18396 7196 18452
rect 7252 18396 11340 18452
rect 11396 18396 11406 18452
rect 21522 18396 21532 18452
rect 21588 18396 23660 18452
rect 23716 18396 23726 18452
rect 41346 18396 41356 18452
rect 41412 18396 42588 18452
rect 42644 18396 42654 18452
rect 44604 18396 47068 18452
rect 47124 18396 47134 18452
rect 16482 18284 16492 18340
rect 16548 18284 21868 18340
rect 21924 18284 21934 18340
rect 26114 18172 26124 18228
rect 26180 18172 31836 18228
rect 31892 18172 31902 18228
rect 42802 18060 42812 18116
rect 42868 18060 44716 18116
rect 44772 18060 44782 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 6178 17724 6188 17780
rect 6244 17724 8652 17780
rect 8708 17724 8718 17780
rect 24098 17724 24108 17780
rect 24164 17724 28252 17780
rect 28308 17724 28318 17780
rect 45938 17500 45948 17556
rect 46004 17500 49644 17556
rect 49700 17500 49710 17556
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 32722 16940 32732 16996
rect 32788 16940 35308 16996
rect 35364 16940 35374 16996
rect 20402 16716 20412 16772
rect 20468 16716 24332 16772
rect 24388 16716 24398 16772
rect 19730 16604 19740 16660
rect 19796 16604 20300 16660
rect 20356 16604 20366 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 9874 15932 9884 15988
rect 9940 15932 10892 15988
rect 10948 15932 10958 15988
rect 24546 15932 24556 15988
rect 24612 15932 27244 15988
rect 27300 15932 27310 15988
rect 41682 15932 41692 15988
rect 41748 15932 43708 15988
rect 43764 15932 43774 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 54012 40236 54068 40292
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 54012 39676 54068 39732
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 41356 22764 41412 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 44828 22652 44884 22708
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 41356 21644 41412 21700
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 44828 19740 44884 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 63532 4768 64348
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 64316 20128 64348
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 63532 35488 64348
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 50528 64316 50848 64348
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 65888 63532 66208 64348
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 54012 40292 54068 40302
rect 54012 39732 54068 40236
rect 54012 39666 54068 39676
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 41356 22820 41412 22830
rect 41356 21700 41412 22764
rect 41356 21634 41412 21644
rect 44828 22708 44884 22718
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 44828 19796 44884 22652
rect 44828 19730 44884 19740
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _294_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37520 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _295_
timestamp 1698431365
transform -1 0 30352 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _296_
timestamp 1698431365
transform -1 0 34272 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _297_
timestamp 1698431365
transform -1 0 30912 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _298_
timestamp 1698431365
transform -1 0 33600 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _299_
timestamp 1698431365
transform 1 0 39648 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _300_
timestamp 1698431365
transform -1 0 36624 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _301_
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _302_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _303_
timestamp 1698431365
transform -1 0 43456 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _304_
timestamp 1698431365
transform 1 0 42448 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _305_
timestamp 1698431365
transform -1 0 45248 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _306_
timestamp 1698431365
transform 1 0 45808 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _307_
timestamp 1698431365
transform -1 0 44128 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _308_
timestamp 1698431365
transform -1 0 42448 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _309_
timestamp 1698431365
transform 1 0 43120 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _310_
timestamp 1698431365
transform -1 0 45696 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _311_
timestamp 1698431365
transform 1 0 51296 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _312_
timestamp 1698431365
transform -1 0 50960 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _313_
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _314_
timestamp 1698431365
transform 1 0 48160 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _315_
timestamp 1698431365
transform 1 0 55328 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _316_
timestamp 1698431365
transform 1 0 51072 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _317_
timestamp 1698431365
transform -1 0 54432 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _318_
timestamp 1698431365
transform 1 0 54656 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _319_
timestamp 1698431365
transform 1 0 55328 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _320_
timestamp 1698431365
transform -1 0 50512 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _321_
timestamp 1698431365
transform 1 0 50736 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _322_
timestamp 1698431365
transform -1 0 52304 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _323_
timestamp 1698431365
transform -1 0 54880 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _324_
timestamp 1698431365
transform 1 0 59248 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _325_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _326_
timestamp 1698431365
transform -1 0 49728 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _327_
timestamp 1698431365
transform 1 0 49728 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _328_
timestamp 1698431365
transform 1 0 51184 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _329_
timestamp 1698431365
transform -1 0 58800 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _330_
timestamp 1698431365
transform -1 0 62720 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _331_
timestamp 1698431365
transform -1 0 59808 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _332_
timestamp 1698431365
transform -1 0 56224 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _333_
timestamp 1698431365
transform -1 0 51968 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _334_
timestamp 1698431365
transform 1 0 51744 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _335_
timestamp 1698431365
transform 1 0 54432 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _336_
timestamp 1698431365
transform 1 0 44576 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _337_
timestamp 1698431365
transform -1 0 42000 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _338_
timestamp 1698431365
transform 1 0 43456 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _339_
timestamp 1698431365
transform -1 0 45696 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _340_
timestamp 1698431365
transform -1 0 38752 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _341_
timestamp 1698431365
transform -1 0 43904 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _342_
timestamp 1698431365
transform -1 0 40320 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _343_
timestamp 1698431365
transform -1 0 44240 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _344_
timestamp 1698431365
transform -1 0 46032 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _345_
timestamp 1698431365
transform 1 0 46032 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _346_
timestamp 1698431365
transform 1 0 46704 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _347_
timestamp 1698431365
transform 1 0 45472 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _348_
timestamp 1698431365
transform -1 0 50176 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _349_
timestamp 1698431365
transform -1 0 52192 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _350_
timestamp 1698431365
transform -1 0 54656 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _351_
timestamp 1698431365
transform 1 0 55216 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _352_
timestamp 1698431365
transform -1 0 59920 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _353_
timestamp 1698431365
transform -1 0 59808 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _354_
timestamp 1698431365
transform -1 0 59472 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _355_
timestamp 1698431365
transform 1 0 49728 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _356_
timestamp 1698431365
transform 1 0 51296 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _357_
timestamp 1698431365
transform -1 0 55440 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _358_
timestamp 1698431365
transform 1 0 41216 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _359_
timestamp 1698431365
transform -1 0 41440 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _360_
timestamp 1698431365
transform -1 0 42448 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _361_
timestamp 1698431365
transform -1 0 40544 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _362_
timestamp 1698431365
transform -1 0 43120 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _363_
timestamp 1698431365
transform 1 0 43120 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _364_
timestamp 1698431365
transform -1 0 47376 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _365_
timestamp 1698431365
transform 1 0 47040 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _366_
timestamp 1698431365
transform -1 0 46704 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _367_
timestamp 1698431365
transform 1 0 46368 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _368_
timestamp 1698431365
transform 1 0 47376 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _369_
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _370_
timestamp 1698431365
transform -1 0 30016 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _371_
timestamp 1698431365
transform -1 0 32144 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _372_
timestamp 1698431365
transform -1 0 30464 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _373_
timestamp 1698431365
transform -1 0 29792 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _374_
timestamp 1698431365
transform 1 0 30576 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _375_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _376_
timestamp 1698431365
transform 1 0 33712 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _377_
timestamp 1698431365
transform 1 0 35840 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _378_
timestamp 1698431365
transform 1 0 32032 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _379_
timestamp 1698431365
transform 1 0 35840 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _380_
timestamp 1698431365
transform -1 0 28000 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _381_
timestamp 1698431365
transform -1 0 24528 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _382_
timestamp 1698431365
transform -1 0 24976 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _383_
timestamp 1698431365
transform 1 0 26992 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _384_
timestamp 1698431365
transform 1 0 28112 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _385_
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _386_
timestamp 1698431365
transform 1 0 21504 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _387_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _388_
timestamp 1698431365
transform -1 0 26208 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _389_
timestamp 1698431365
transform -1 0 25760 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _390_
timestamp 1698431365
transform 1 0 28000 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _391_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _392_
timestamp 1698431365
transform -1 0 32480 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _393_
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _394_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _395_
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _396_
timestamp 1698431365
transform -1 0 30800 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _397_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _398_
timestamp 1698431365
transform -1 0 33600 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _399_
timestamp 1698431365
transform -1 0 32704 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _400_
timestamp 1698431365
transform -1 0 35280 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _401_
timestamp 1698431365
transform -1 0 36512 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _402_
timestamp 1698431365
transform -1 0 47600 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _403_
timestamp 1698431365
transform -1 0 40544 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _404_
timestamp 1698431365
transform -1 0 43456 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _405_
timestamp 1698431365
transform 1 0 43008 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _406_
timestamp 1698431365
transform -1 0 48160 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _407_
timestamp 1698431365
transform 1 0 47152 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _408_
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _409_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _410_
timestamp 1698431365
transform -1 0 43232 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _411_
timestamp 1698431365
transform -1 0 44128 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _412_
timestamp 1698431365
transform -1 0 45360 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _413_
timestamp 1698431365
transform -1 0 40544 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _414_
timestamp 1698431365
transform -1 0 32592 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _415_
timestamp 1698431365
transform -1 0 34272 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _416_
timestamp 1698431365
transform -1 0 31360 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _417_
timestamp 1698431365
transform -1 0 33600 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _418_
timestamp 1698431365
transform -1 0 33600 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _419_
timestamp 1698431365
transform 1 0 34048 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _420_
timestamp 1698431365
transform -1 0 37520 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _421_
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _422_
timestamp 1698431365
transform -1 0 37520 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _423_
timestamp 1698431365
transform 1 0 37968 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _424_
timestamp 1698431365
transform 1 0 25200 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _425_
timestamp 1698431365
transform -1 0 17136 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _426_
timestamp 1698431365
transform -1 0 15120 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _427_
timestamp 1698431365
transform 1 0 18032 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _428_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _429_
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _430_
timestamp 1698431365
transform -1 0 14224 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _431_
timestamp 1698431365
transform -1 0 16352 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _432_
timestamp 1698431365
transform -1 0 10416 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _433_
timestamp 1698431365
transform -1 0 16688 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _434_
timestamp 1698431365
transform -1 0 17920 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _435_
timestamp 1698431365
transform -1 0 18032 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _436_
timestamp 1698431365
transform -1 0 24080 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _437_
timestamp 1698431365
transform 1 0 19600 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _438_
timestamp 1698431365
transform -1 0 21840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _439_
timestamp 1698431365
transform 1 0 22736 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _440_
timestamp 1698431365
transform -1 0 22736 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _441_
timestamp 1698431365
transform 1 0 25648 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _442_
timestamp 1698431365
transform -1 0 26096 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _443_
timestamp 1698431365
transform 1 0 26320 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _444_
timestamp 1698431365
transform 1 0 19600 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _445_
timestamp 1698431365
transform -1 0 20944 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _446_
timestamp 1698431365
transform -1 0 25760 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _447_
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _448_
timestamp 1698431365
transform -1 0 21840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _449_
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _450_
timestamp 1698431365
transform -1 0 27440 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _451_
timestamp 1698431365
transform -1 0 24864 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _452_
timestamp 1698431365
transform -1 0 21840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _453_
timestamp 1698431365
transform 1 0 22176 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _454_
timestamp 1698431365
transform -1 0 23520 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _455_
timestamp 1698431365
transform 1 0 23520 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _456_
timestamp 1698431365
transform -1 0 26880 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _457_
timestamp 1698431365
transform 1 0 27328 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _458_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _459_
timestamp 1698431365
transform -1 0 11088 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _460_
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _461_
timestamp 1698431365
transform -1 0 14224 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _462_
timestamp 1698431365
transform 1 0 16240 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _463_
timestamp 1698431365
transform -1 0 8960 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _464_
timestamp 1698431365
transform -1 0 10080 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _465_
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _466_
timestamp 1698431365
transform -1 0 6720 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _467_
timestamp 1698431365
transform -1 0 7392 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _468_
timestamp 1698431365
transform 1 0 7392 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _469_
timestamp 1698431365
transform 1 0 9520 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _470_
timestamp 1698431365
transform -1 0 10752 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _471_
timestamp 1698431365
transform 1 0 12096 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _472_
timestamp 1698431365
transform -1 0 14224 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _473_
timestamp 1698431365
transform 1 0 14896 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _474_
timestamp 1698431365
transform -1 0 17024 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _475_
timestamp 1698431365
transform 1 0 17584 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _476_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _477_
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _478_
timestamp 1698431365
transform -1 0 14000 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _479_
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _480_
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _481_
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _482_
timestamp 1698431365
transform -1 0 30240 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _483_
timestamp 1698431365
transform -1 0 29680 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _484_
timestamp 1698431365
transform 1 0 31360 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _485_
timestamp 1698431365
transform -1 0 34160 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _486_
timestamp 1698431365
transform -1 0 29680 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _487_
timestamp 1698431365
transform -1 0 30688 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _488_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _489_
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _490_
timestamp 1698431365
transform -1 0 35392 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _491_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _492_
timestamp 1698431365
transform -1 0 38416 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _493_
timestamp 1698431365
transform 1 0 38752 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _494_
timestamp 1698431365
transform 1 0 39424 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _495_
timestamp 1698431365
transform -1 0 36064 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _496_
timestamp 1698431365
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _497_
timestamp 1698431365
transform -1 0 38752 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _498_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _499_
timestamp 1698431365
transform 1 0 30464 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _500_
timestamp 1698431365
transform -1 0 33600 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _501_
timestamp 1698431365
transform -1 0 34272 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _502_
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _503_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _504_
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _505_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _506_
timestamp 1698431365
transform -1 0 22064 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _507_
timestamp 1698431365
transform -1 0 22064 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _508_
timestamp 1698431365
transform -1 0 18704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _509_
timestamp 1698431365
transform 1 0 17808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _510_
timestamp 1698431365
transform -1 0 20160 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _511_
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _512_
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _513_
timestamp 1698431365
transform -1 0 15232 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _514_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _515_
timestamp 1698431365
transform -1 0 6720 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _516_
timestamp 1698431365
transform -1 0 10080 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _517_
timestamp 1698431365
transform -1 0 11200 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _518_
timestamp 1698431365
transform 1 0 11760 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _519_
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _520_
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _521_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _522_
timestamp 1698431365
transform -1 0 11200 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _523_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _524_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _525_
timestamp 1698431365
transform -1 0 15456 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _526_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _527_
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _528_
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _529_
timestamp 1698431365
transform -1 0 19040 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _530_
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _531_
timestamp 1698431365
transform 1 0 21728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _532_
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _533_
timestamp 1698431365
transform -1 0 19600 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _534_
timestamp 1698431365
transform 1 0 21280 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _535_
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _536_
timestamp 1698431365
transform -1 0 24416 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _537_
timestamp 1698431365
transform 1 0 20272 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _538_
timestamp 1698431365
transform -1 0 23072 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _539_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _540_
timestamp 1698431365
transform 1 0 25424 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _541_
timestamp 1698431365
transform 1 0 48608 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _542_
timestamp 1698431365
transform -1 0 55440 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _543_
timestamp 1698431365
transform -1 0 52192 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _544_
timestamp 1698431365
transform -1 0 48384 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _545_
timestamp 1698431365
transform -1 0 49728 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _546_
timestamp 1698431365
transform -1 0 52192 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _547_
timestamp 1698431365
transform -1 0 52080 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _548_
timestamp 1698431365
transform 1 0 52640 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _549_
timestamp 1698431365
transform 1 0 54096 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _550_
timestamp 1698431365
transform -1 0 56224 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _551_
timestamp 1698431365
transform 1 0 59136 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _552_
timestamp 1698431365
transform 1 0 49056 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _553_
timestamp 1698431365
transform 1 0 51296 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _554_
timestamp 1698431365
transform -1 0 51296 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _555_
timestamp 1698431365
transform -1 0 58800 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _556_
timestamp 1698431365
transform 1 0 54208 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _557_
timestamp 1698431365
transform 1 0 59248 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _558_
timestamp 1698431365
transform -1 0 56112 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _559_
timestamp 1698431365
transform 1 0 59360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _560_
timestamp 1698431365
transform -1 0 55664 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _561_
timestamp 1698431365
transform 1 0 55216 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _562_
timestamp 1698431365
transform -1 0 59808 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _563_
timestamp 1698431365
transform -1 0 51408 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _564_
timestamp 1698431365
transform -1 0 48160 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _565_
timestamp 1698431365
transform 1 0 49952 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _566_
timestamp 1698431365
transform -1 0 46592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _567_
timestamp 1698431365
transform -1 0 49952 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _568_
timestamp 1698431365
transform -1 0 43904 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _569_
timestamp 1698431365
transform -1 0 44464 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _570_
timestamp 1698431365
transform -1 0 47264 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _571_
timestamp 1698431365
transform 1 0 46704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _572_
timestamp 1698431365
transform 1 0 47264 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _573_
timestamp 1698431365
transform 1 0 47712 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _574_
timestamp 1698431365
transform 1 0 45136 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _575_
timestamp 1698431365
transform -1 0 41440 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _576_
timestamp 1698431365
transform -1 0 42112 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _577_
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _578_
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _579_
timestamp 1698431365
transform -1 0 40432 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _580_
timestamp 1698431365
transform -1 0 39760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _581_
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _582_
timestamp 1698431365
transform -1 0 42896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _583_
timestamp 1698431365
transform -1 0 44240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _584_
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _585_
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _586_
timestamp 1698431365
transform -1 0 34832 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _587_
timestamp 1698431365
transform -1 0 36400 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _588_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49952 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _589_
timestamp 1698431365
transform 1 0 44576 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _590_
timestamp 1698431365
transform 1 0 45248 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _591_
timestamp 1698431365
transform 1 0 44800 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _592_
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _593_
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _594_
timestamp 1698431365
transform -1 0 56224 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _595_
timestamp 1698431365
transform 1 0 52416 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _596_
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _597_
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _598_
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _599_
timestamp 1698431365
transform 1 0 48496 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _600_
timestamp 1698431365
transform 1 0 48832 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _601_
timestamp 1698431365
transform 1 0 52416 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _602_
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _603_
timestamp 1698431365
transform 1 0 51184 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _604_
timestamp 1698431365
transform 1 0 52752 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _605_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _606_
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _607_
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _608_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _609_
timestamp 1698431365
transform 1 0 44576 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _610_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _611_
timestamp 1698431365
transform -1 0 45360 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _612_
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _613_
timestamp 1698431365
transform 1 0 40656 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _614_
timestamp 1698431365
transform 1 0 42112 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _615_
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _616_
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _617_
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _618_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _619_
timestamp 1698431365
transform -1 0 44464 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _620_
timestamp 1698431365
transform 1 0 40656 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _621_
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _622_
timestamp 1698431365
transform -1 0 40656 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _623_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _624_
timestamp 1698431365
transform 1 0 36736 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _625_
timestamp 1698431365
transform 1 0 38416 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _626_
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _627_
timestamp 1698431365
transform 1 0 41328 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _628_
timestamp 1698431365
transform -1 0 36736 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _629_
timestamp 1698431365
transform 1 0 32816 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _630_
timestamp 1698431365
transform -1 0 36736 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _631_
timestamp 1698431365
transform -1 0 32480 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _632_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _633_
timestamp 1698431365
transform -1 0 32704 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _634_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _635_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _636_
timestamp 1698431365
transform 1 0 32816 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _637_
timestamp 1698431365
transform 1 0 34160 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _638_
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _639_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _640_
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _641_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _642_
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _643_
timestamp 1698431365
transform 1 0 37968 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _644_
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _645_
timestamp 1698431365
transform 1 0 42224 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _646_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _647_
timestamp 1698431365
transform 1 0 44576 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _648_
timestamp 1698431365
transform 1 0 52976 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _649_
timestamp 1698431365
transform 1 0 48496 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _650_
timestamp 1698431365
transform 1 0 49952 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _651_
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _652_
timestamp 1698431365
transform 1 0 52640 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _653_
timestamp 1698431365
transform 1 0 46928 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _654_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _655_
timestamp 1698431365
transform 1 0 48496 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _656_
timestamp 1698431365
transform 1 0 50512 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _657_
timestamp 1698431365
transform 1 0 52416 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _658_
timestamp 1698431365
transform 1 0 45920 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _659_
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _660_
timestamp 1698431365
transform 1 0 48496 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _661_
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _662_
timestamp 1698431365
transform 1 0 56336 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _663_
timestamp 1698431365
transform 1 0 52416 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _664_
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _665_
timestamp 1698431365
transform 1 0 47376 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _666_
timestamp 1698431365
transform 1 0 49504 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _667_
timestamp 1698431365
transform 1 0 52416 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _668_
timestamp 1698431365
transform 1 0 36736 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _669_
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _670_
timestamp 1698431365
transform -1 0 46144 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _671_
timestamp 1698431365
transform -1 0 39648 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _672_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _673_
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _674_
timestamp 1698431365
transform 1 0 40656 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _675_
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _676_
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _677_
timestamp 1698431365
transform 1 0 44576 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _678_
timestamp 1698431365
transform -1 0 52416 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _679_
timestamp 1698431365
transform 1 0 48496 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _680_
timestamp 1698431365
transform 1 0 50176 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _681_
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _682_
timestamp 1698431365
transform -1 0 56224 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _683_
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _684_
timestamp 1698431365
transform 1 0 52416 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _685_
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _686_
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _687_
timestamp 1698431365
transform -1 0 54768 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _688_
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _689_
timestamp 1698431365
transform -1 0 41216 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _690_
timestamp 1698431365
transform 1 0 36736 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _691_
timestamp 1698431365
transform 1 0 37968 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _692_
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _693_
timestamp 1698431365
transform 1 0 42224 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _694_
timestamp 1698431365
transform -1 0 48384 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _695_
timestamp 1698431365
transform 1 0 41664 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _696_
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _697_
timestamp 1698431365
transform 1 0 44912 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _698_
timestamp 1698431365
transform 1 0 24976 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _699_
timestamp 1698431365
transform -1 0 32816 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _700_
timestamp 1698431365
transform 1 0 24976 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _701_
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _702_
timestamp 1698431365
transform 1 0 27888 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _703_
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _704_
timestamp 1698431365
transform 1 0 31472 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _705_
timestamp 1698431365
transform 1 0 32816 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _706_
timestamp 1698431365
transform -1 0 36736 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _707_
timestamp 1698431365
transform 1 0 32816 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _708_
timestamp 1698431365
transform -1 0 24528 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _709_
timestamp 1698431365
transform -1 0 24976 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _710_
timestamp 1698431365
transform 1 0 24304 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _711_
timestamp 1698431365
transform -1 0 28784 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _712_
timestamp 1698431365
transform -1 0 20944 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _713_
timestamp 1698431365
transform 1 0 20720 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _714_
timestamp 1698431365
transform -1 0 20944 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _715_
timestamp 1698431365
transform 1 0 20720 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _716_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _717_
timestamp 1698431365
transform 1 0 24192 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _718_
timestamp 1698431365
transform -1 0 31808 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _719_
timestamp 1698431365
transform 1 0 28896 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _720_
timestamp 1698431365
transform 1 0 32144 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _721_
timestamp 1698431365
transform 1 0 33488 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _722_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _723_
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _724_
timestamp 1698431365
transform -1 0 31696 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _725_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _726_
timestamp 1698431365
transform 1 0 31472 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _727_
timestamp 1698431365
transform -1 0 36624 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _728_
timestamp 1698431365
transform 1 0 37968 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _729_
timestamp 1698431365
transform 1 0 38976 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _730_
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _731_
timestamp 1698431365
transform 1 0 44576 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _732_
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _733_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _734_
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _735_
timestamp 1698431365
transform -1 0 41552 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _736_
timestamp 1698431365
transform 1 0 38752 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _737_
timestamp 1698431365
transform 1 0 40880 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _738_
timestamp 1698431365
transform 1 0 28112 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _739_
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _740_
timestamp 1698431365
transform -1 0 32144 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _741_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _742_
timestamp 1698431365
transform 1 0 28896 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _743_
timestamp 1698431365
transform 1 0 31360 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _744_
timestamp 1698431365
transform 1 0 32816 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _745_
timestamp 1698431365
transform 1 0 34832 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _746_
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _747_
timestamp 1698431365
transform 1 0 35616 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _748_
timestamp 1698431365
transform -1 0 15680 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _749_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _750_
timestamp 1698431365
transform -1 0 18928 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _751_
timestamp 1698431365
transform -1 0 14896 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _752_
timestamp 1698431365
transform 1 0 9296 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _753_
timestamp 1698431365
transform 1 0 9296 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _754_
timestamp 1698431365
transform -1 0 15456 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _755_
timestamp 1698431365
transform 1 0 13216 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _756_
timestamp 1698431365
transform 1 0 13216 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _757_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _758_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _759_
timestamp 1698431365
transform 1 0 17136 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _760_
timestamp 1698431365
transform 1 0 20048 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _761_
timestamp 1698431365
transform -1 0 24864 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _762_
timestamp 1698431365
transform 1 0 23744 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _763_
timestamp 1698431365
transform -1 0 24864 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _764_
timestamp 1698431365
transform 1 0 23968 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _765_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _766_
timestamp 1698431365
transform -1 0 22960 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _767_
timestamp 1698431365
transform 1 0 21056 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _768_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _769_
timestamp 1698431365
transform -1 0 28784 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _770_
timestamp 1698431365
transform 1 0 23968 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _771_
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _772_
timestamp 1698431365
transform 1 0 17136 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _773_
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _774_
timestamp 1698431365
transform 1 0 17136 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _775_
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _776_
timestamp 1698431365
transform -1 0 27328 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _777_
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _778_
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _779_
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _780_
timestamp 1698431365
transform -1 0 15680 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _781_
timestamp 1698431365
transform 1 0 12096 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _782_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _783_
timestamp 1698431365
transform -1 0 10528 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _784_
timestamp 1698431365
transform 1 0 8960 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _785_
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _786_
timestamp 1698431365
transform -1 0 8176 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _787_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _788_
timestamp 1698431365
transform -1 0 11872 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _789_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _790_
timestamp 1698431365
transform 1 0 9296 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _791_
timestamp 1698431365
transform 1 0 12432 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _792_
timestamp 1698431365
transform 1 0 13216 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _793_
timestamp 1698431365
transform -1 0 19376 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _794_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _795_
timestamp 1698431365
transform -1 0 12880 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _796_
timestamp 1698431365
transform 1 0 8512 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _797_
timestamp 1698431365
transform -1 0 12096 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _798_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _799_
timestamp 1698431365
transform -1 0 31248 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _800_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _801_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _802_
timestamp 1698431365
transform -1 0 34720 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _803_
timestamp 1698431365
transform 1 0 24752 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _804_
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _805_
timestamp 1698431365
transform 1 0 28896 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _806_
timestamp 1698431365
transform 1 0 31360 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _807_
timestamp 1698431365
transform -1 0 36736 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _808_
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _809_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _810_
timestamp 1698431365
transform -1 0 40656 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _811_
timestamp 1698431365
transform -1 0 35280 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _812_
timestamp 1698431365
transform 1 0 32816 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _813_
timestamp 1698431365
transform -1 0 39536 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _814_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _815_
timestamp 1698431365
transform 1 0 27776 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _816_
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _817_
timestamp 1698431365
transform -1 0 35392 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _818_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _819_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _820_
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _821_
timestamp 1698431365
transform -1 0 23744 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _822_
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _823_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _824_
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _825_
timestamp 1698431365
transform -1 0 21056 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _826_
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _827_
timestamp 1698431365
transform -1 0 27776 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _828_
timestamp 1698431365
transform -1 0 13216 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _829_
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _830_
timestamp 1698431365
transform 1 0 5376 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _831_
timestamp 1698431365
transform 1 0 5376 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _832_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _833_
timestamp 1698431365
transform -1 0 7840 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _834_
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _835_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _836_
timestamp 1698431365
transform -1 0 13216 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _837_
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _838_
timestamp 1698431365
transform -1 0 17024 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _839_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _840_
timestamp 1698431365
transform 1 0 13216 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _841_
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _842_
timestamp 1698431365
transform -1 0 21056 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _843_
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _844_
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _845_
timestamp 1698431365
transform -1 0 24192 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _846_
timestamp 1698431365
transform 1 0 13216 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _847_
timestamp 1698431365
transform 1 0 21056 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _848_
timestamp 1698431365
transform -1 0 23632 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _849_
timestamp 1698431365
transform 1 0 17136 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _850_
timestamp 1698431365
transform -1 0 24976 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _851_
timestamp 1698431365
transform 1 0 17136 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1698431365
transform -1 0 48160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__I
timestamp 1698431365
transform 1 0 48832 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__I
timestamp 1698431365
transform 1 0 50624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__I
timestamp 1698431365
transform -1 0 51968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__I
timestamp 1698431365
transform 1 0 50736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__I
timestamp 1698431365
transform 1 0 59696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__I
timestamp 1698431365
transform 1 0 62944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__I
timestamp 1698431365
transform 1 0 59472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__I
timestamp 1698431365
transform 1 0 59472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__I
timestamp 1698431365
transform 1 0 52080 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__I
timestamp 1698431365
transform 1 0 56672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__I
timestamp 1698431365
transform 1 0 56672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I
timestamp 1698431365
transform 1 0 44912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__I
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1698431365
transform -1 0 49504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__I
timestamp 1698431365
transform 1 0 52752 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I
timestamp 1698431365
transform -1 0 55104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__I
timestamp 1698431365
transform 1 0 55552 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I
timestamp 1698431365
transform 1 0 59360 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__I
timestamp 1698431365
transform 1 0 60592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1698431365
transform 1 0 59472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__I
timestamp 1698431365
transform 1 0 51072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I
timestamp 1698431365
transform 1 0 48160 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I
timestamp 1698431365
transform 1 0 57120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__I
timestamp 1698431365
transform 1 0 40992 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__I
timestamp 1698431365
transform -1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__I
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__I
timestamp 1698431365
transform 1 0 24080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__I
timestamp 1698431365
transform 1 0 28112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__I
timestamp 1698431365
transform 1 0 25424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__I
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__I
timestamp 1698431365
transform 1 0 17920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__I
timestamp 1698431365
transform 1 0 22400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__I
timestamp 1698431365
transform -1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__I
timestamp 1698431365
transform 1 0 25312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__I
timestamp 1698431365
transform -1 0 26208 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__I
timestamp 1698431365
transform -1 0 28000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__I
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__I
timestamp 1698431365
transform -1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__I
timestamp 1698431365
transform 1 0 37408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1698431365
transform 1 0 18480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__I
timestamp 1698431365
transform 1 0 28448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__I
timestamp 1698431365
transform 1 0 15904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__I
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__I
timestamp 1698431365
transform 1 0 27216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__I
timestamp 1698431365
transform 1 0 26992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__I
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__I
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__I
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__I
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__I
timestamp 1698431365
transform 1 0 19712 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__I
timestamp 1698431365
transform 1 0 17584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__I
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__I
timestamp 1698431365
transform -1 0 14784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__I
timestamp 1698431365
transform 1 0 17584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__I
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__I
timestamp 1698431365
transform 1 0 25424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__I
timestamp 1698431365
transform 1 0 15456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__I
timestamp 1698431365
transform -1 0 20384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__I
timestamp 1698431365
transform -1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__I
timestamp 1698431365
transform 1 0 26656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__I
timestamp 1698431365
transform -1 0 19600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__I
timestamp 1698431365
transform 1 0 22176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__I
timestamp 1698431365
transform 1 0 23184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__I
timestamp 1698431365
transform -1 0 49392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__I
timestamp 1698431365
transform 1 0 51968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__I
timestamp 1698431365
transform 1 0 50848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__I
timestamp 1698431365
transform -1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__I
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__CLK
timestamp 1698431365
transform -1 0 52864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__CLK
timestamp 1698431365
transform -1 0 49280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__CLK
timestamp 1698431365
transform 1 0 49616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__CLK
timestamp 1698431365
transform 1 0 49168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__CLK
timestamp 1698431365
transform 1 0 57120 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__CLK
timestamp 1698431365
transform 1 0 57008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__CLK
timestamp 1698431365
transform 1 0 56560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__CLK
timestamp 1698431365
transform 1 0 60480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__607__CLK
timestamp 1698431365
transform 1 0 56560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__CLK
timestamp 1698431365
transform 1 0 53088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__CLK
timestamp 1698431365
transform 1 0 46032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__CLK
timestamp 1698431365
transform -1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__CLK
timestamp 1698431365
transform -1 0 45584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__613__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__CLK
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__CLK
timestamp 1698431365
transform -1 0 45136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__619__CLK
timestamp 1698431365
transform 1 0 47152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__CLK
timestamp 1698431365
transform 1 0 46256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__CLK
timestamp 1698431365
transform 1 0 44912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__CLK
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__CLK
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__D
timestamp 1698431365
transform -1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__CLK
timestamp 1698431365
transform 1 0 35056 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__CLK
timestamp 1698431365
transform -1 0 35728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__D
timestamp 1698431365
transform -1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__CLK
timestamp 1698431365
transform 1 0 46704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__641__CLK
timestamp 1698431365
transform 1 0 49280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__D
timestamp 1698431365
transform -1 0 45472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__643__CLK
timestamp 1698431365
transform 1 0 45696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__CLK
timestamp 1698431365
transform 1 0 48720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__CLK
timestamp 1698431365
transform 1 0 51184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__648__CLK
timestamp 1698431365
transform 1 0 57008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__CLK
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__CLK
timestamp 1698431365
transform 1 0 53760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__CLK
timestamp 1698431365
transform 1 0 56560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__CLK
timestamp 1698431365
transform -1 0 56896 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__CLK
timestamp 1698431365
transform 1 0 52752 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__CLK
timestamp 1698431365
transform -1 0 56896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__660__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__661__CLK
timestamp 1698431365
transform 1 0 59472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__662__CLK
timestamp 1698431365
transform 1 0 56560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__CLK
timestamp 1698431365
transform 1 0 57120 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__CLK
timestamp 1698431365
transform 1 0 57008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__CLK
timestamp 1698431365
transform -1 0 56784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__667__CLK
timestamp 1698431365
transform 1 0 57120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__676__CLK
timestamp 1698431365
transform 1 0 47712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__CLK
timestamp 1698431365
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__CLK
timestamp 1698431365
transform 1 0 53088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__CLK
timestamp 1698431365
transform -1 0 55552 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__CLK
timestamp 1698431365
transform 1 0 56560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__CLK
timestamp 1698431365
transform 1 0 57120 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__683__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__CLK
timestamp 1698431365
transform 1 0 57008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__CLK
timestamp 1698431365
transform 1 0 52640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__CLK
timestamp 1698431365
transform 1 0 57120 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__CLK
timestamp 1698431365
transform 1 0 42000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__CLK
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__CLK
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__CLK
timestamp 1698431365
transform 1 0 49280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__CLK
timestamp 1698431365
transform 1 0 49504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__CLK
timestamp 1698431365
transform 1 0 48720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__CLK
timestamp 1698431365
transform 1 0 49168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__CLK
timestamp 1698431365
transform 1 0 41776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__D
timestamp 1698431365
transform 1 0 45360 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__CLK
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__CLK
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__745__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__747__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__748__CLK
timestamp 1698431365
transform 1 0 15232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__751__CLK
timestamp 1698431365
transform -1 0 10080 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__765__CLK
timestamp 1698431365
transform -1 0 23408 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__766__CLK
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__768__CLK
timestamp 1698431365
transform -1 0 16352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__769__CLK
timestamp 1698431365
transform -1 0 25536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__770__CLK
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__771__CLK
timestamp 1698431365
transform -1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__772__CLK
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__773__CLK
timestamp 1698431365
transform 1 0 23968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__774__CLK
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__775__CLK
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__776__CLK
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__777__CLK
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__778__CLK
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__779__CLK
timestamp 1698431365
transform 1 0 8064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__780__CLK
timestamp 1698431365
transform 1 0 11424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__782__CLK
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__783__CLK
timestamp 1698431365
transform 1 0 11424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__784__CLK
timestamp 1698431365
transform 1 0 8736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__785__CLK
timestamp 1698431365
transform 1 0 8288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__786__CLK
timestamp 1698431365
transform -1 0 8736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__787__CLK
timestamp 1698431365
transform 1 0 7616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__788__CLK
timestamp 1698431365
transform 1 0 11872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__789__CLK
timestamp 1698431365
transform 1 0 12208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__790__CLK
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__791__CLK
timestamp 1698431365
transform 1 0 14672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__792__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__793__CLK
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__794__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__795__CLK
timestamp 1698431365
transform 1 0 8848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__797__CLK
timestamp 1698431365
transform -1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__798__CLK
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__800__CLK
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__803__CLK
timestamp 1698431365
transform 1 0 30912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__804__CLK
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__805__CLK
timestamp 1698431365
transform 1 0 27440 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__809__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__810__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__813__CLK
timestamp 1698431365
transform 1 0 39760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__814__CLK
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__815__CLK
timestamp 1698431365
transform 1 0 27552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__816__CLK
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__818__CLK
timestamp 1698431365
transform -1 0 23968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__819__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__820__CLK
timestamp 1698431365
transform 1 0 26992 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__821__CLK
timestamp 1698431365
transform -1 0 24192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__822__CLK
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__823__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__825__CLK
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__826__CLK
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__827__CLK
timestamp 1698431365
transform -1 0 28224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__829__CLK
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__830__CLK
timestamp 1698431365
transform 1 0 5824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__831__CLK
timestamp 1698431365
transform -1 0 8512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__835__CLK
timestamp 1698431365
transform -1 0 8064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__839__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__841__CLK
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__842__CLK
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__843__CLK
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__844__CLK
timestamp 1698431365
transform -1 0 23968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__845__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__847__CLK
timestamp 1698431365
transform 1 0 24528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__848__CLK
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__849__CLK
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__850__CLK
timestamp 1698431365
transform 1 0 19264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__850__D
timestamp 1698431365
transform -1 0 20944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__851__CLK
timestamp 1698431365
transform 1 0 18928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform -1 0 30016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_prog_clk_I
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_prog_clk_I
timestamp 1698431365
transform 1 0 23520 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_prog_clk_I
timestamp 1698431365
transform 1 0 29232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_prog_clk_I
timestamp 1698431365
transform 1 0 20272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_prog_clk_I
timestamp 1698431365
transform 1 0 30912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_prog_clk_I
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_prog_clk_I
timestamp 1698431365
transform 1 0 40880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_prog_clk_I
timestamp 1698431365
transform 1 0 42896 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_prog_clk_I
timestamp 1698431365
transform 1 0 45696 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_prog_clk_I
timestamp 1698431365
transform 1 0 56672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_prog_clk_I
timestamp 1698431365
transform 1 0 52752 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_prog_clk_I
timestamp 1698431365
transform 1 0 41328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_prog_clk_I
timestamp 1698431365
transform 1 0 43568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_prog_clk_I
timestamp 1698431365
transform 1 0 46704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_prog_clk_I
timestamp 1698431365
transform 1 0 52192 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_prog_clk_I
timestamp 1698431365
transform -1 0 53088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_prog_clk_I
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_prog_clk_I
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_prog_clk_I
timestamp 1698431365
transform 1 0 38864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_prog_clk_I
timestamp 1698431365
transform 1 0 25984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_prog_clk_I
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_prog_clk_I
timestamp 1698431365
transform -1 0 26992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_prog_clk_I
timestamp 1698431365
transform 1 0 16352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold229_I
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold261_I
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_prog_clk
timestamp 1698431365
transform -1 0 12432 0 1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_prog_clk
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_prog_clk
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_prog_clk
timestamp 1698431365
transform 1 0 13664 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_prog_clk
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_prog_clk
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_prog_clk
timestamp 1698431365
transform 1 0 34944 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_prog_clk
timestamp 1698431365
transform -1 0 42672 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_prog_clk
timestamp 1698431365
transform -1 0 51520 0 1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_prog_clk
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_prog_clk
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_prog_clk
timestamp 1698431365
transform 1 0 41552 0 -1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_prog_clk
timestamp 1698431365
transform 1 0 37184 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_prog_clk
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_prog_clk
timestamp 1698431365
transform 1 0 53312 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_prog_clk
timestamp 1698431365
transform -1 0 58128 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_prog_clk
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_prog_clk
timestamp 1698431365
transform -1 0 39312 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_prog_clk
timestamp 1698431365
transform 1 0 34608 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_prog_clk
timestamp 1698431365
transform 1 0 26992 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_prog_clk
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_prog_clk
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_prog_clk
timestamp 1698431365
transform -1 0 18928 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_353
timestamp 1698431365
transform 1 0 40880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_359 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41552 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_367
timestamp 1698431365
transform 1 0 42448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_371
timestamp 1698431365
transform 1 0 42896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698431365
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_383
timestamp 1698431365
transform 1 0 44240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_389 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_420
timestamp 1698431365
transform 1 0 48384 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_425
timestamp 1698431365
transform 1 0 48944 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698431365
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_482
timestamp 1698431365
transform 1 0 55328 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_498
timestamp 1698431365
transform 1 0 57120 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_512
timestamp 1698431365
transform 1 0 58688 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_546
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_580
timestamp 1698431365
transform 1 0 66304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_556
timestamp 1698431365
transform 1 0 63616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_562
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_578
timestamp 1698431365
transform 1 0 66080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_580
timestamp 1698431365
transform 1 0 66304 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_521
timestamp 1698431365
transform 1 0 59696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_527
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_559
timestamp 1698431365
transform 1 0 63952 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_575
timestamp 1698431365
transform 1 0 65744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_579
timestamp 1698431365
transform 1 0 66192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_556
timestamp 1698431365
transform 1 0 63616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_562
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_578
timestamp 1698431365
transform 1 0 66080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_580
timestamp 1698431365
transform 1 0 66304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_559
timestamp 1698431365
transform 1 0 63952 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_575
timestamp 1698431365
transform 1 0 65744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_579
timestamp 1698431365
transform 1 0 66192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_556
timestamp 1698431365
transform 1 0 63616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_562
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_578
timestamp 1698431365
transform 1 0 66080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_580
timestamp 1698431365
transform 1 0 66304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_559
timestamp 1698431365
transform 1 0 63952 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_575
timestamp 1698431365
transform 1 0 65744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_579
timestamp 1698431365
transform 1 0 66192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_578
timestamp 1698431365
transform 1 0 66080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_580
timestamp 1698431365
transform 1 0 66304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_559
timestamp 1698431365
transform 1 0 63952 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_575
timestamp 1698431365
transform 1 0 65744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_579
timestamp 1698431365
transform 1 0 66192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_578
timestamp 1698431365
transform 1 0 66080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_580
timestamp 1698431365
transform 1 0 66304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_559
timestamp 1698431365
transform 1 0 63952 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_575
timestamp 1698431365
transform 1 0 65744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_579
timestamp 1698431365
transform 1 0 66192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_578
timestamp 1698431365
transform 1 0 66080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_580
timestamp 1698431365
transform 1 0 66304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_559
timestamp 1698431365
transform 1 0 63952 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_575
timestamp 1698431365
transform 1 0 65744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_579
timestamp 1698431365
transform 1 0 66192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_578
timestamp 1698431365
transform 1 0 66080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_580
timestamp 1698431365
transform 1 0 66304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_165
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_211
timestamp 1698431365
transform 1 0 24976 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_219
timestamp 1698431365
transform 1 0 25872 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_272
timestamp 1698431365
transform 1 0 31808 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_304
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698431365
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_559
timestamp 1698431365
transform 1 0 63952 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_575
timestamp 1698431365
transform 1 0 65744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_579
timestamp 1698431365
transform 1 0 66192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_166
timestamp 1698431365
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_228
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_236
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_238
timestamp 1698431365
transform 1 0 28000 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_255
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_263
timestamp 1698431365
transform 1 0 30800 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_302
timestamp 1698431365
transform 1 0 35168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_304
timestamp 1698431365
transform 1 0 35392 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_321
timestamp 1698431365
transform 1 0 37296 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_337
timestamp 1698431365
transform 1 0 39088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_578
timestamp 1698431365
transform 1 0 66080 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_580
timestamp 1698431365
transform 1 0 66304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_73
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_91
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_99
timestamp 1698431365
transform 1 0 12432 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_135
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_151
timestamp 1698431365
transform 1 0 18256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_153
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_205
timestamp 1698431365
transform 1 0 24304 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_237
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_271
timestamp 1698431365
transform 1 0 31696 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_288
timestamp 1698431365
transform 1 0 33600 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_305
timestamp 1698431365
transform 1 0 35504 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_341
timestamp 1698431365
transform 1 0 39536 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_357
timestamp 1698431365
transform 1 0 41328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_365
timestamp 1698431365
transform 1 0 42224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698431365
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_559
timestamp 1698431365
transform 1 0 63952 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_575
timestamp 1698431365
transform 1 0 65744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_579
timestamp 1698431365
transform 1 0 66192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698431365
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_120
timestamp 1698431365
transform 1 0 14784 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_164
timestamp 1698431365
transform 1 0 19712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_172
timestamp 1698431365
transform 1 0 20608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_189
timestamp 1698431365
transform 1 0 22512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698431365
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_264
timestamp 1698431365
transform 1 0 30912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_307
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_323
timestamp 1698431365
transform 1 0 37520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_341
timestamp 1698431365
transform 1 0 39536 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_377
timestamp 1698431365
transform 1 0 43568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_385
timestamp 1698431365
transform 1 0 44464 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_402
timestamp 1698431365
transform 1 0 46368 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_418
timestamp 1698431365
transform 1 0 48160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_578
timestamp 1698431365
transform 1 0 66080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_580
timestamp 1698431365
transform 1 0 66304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_61
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_63
timestamp 1698431365
transform 1 0 8400 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_96
timestamp 1698431365
transform 1 0 12096 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_131
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_133
timestamp 1698431365
transform 1 0 16240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_211
timestamp 1698431365
transform 1 0 24976 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_227
timestamp 1698431365
transform 1 0 26768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_263
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_281
timestamp 1698431365
transform 1 0 32816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_289
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_341
timestamp 1698431365
transform 1 0 39536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_361
timestamp 1698431365
transform 1 0 41776 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_377
timestamp 1698431365
transform 1 0 43568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_395
timestamp 1698431365
transform 1 0 45584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_412
timestamp 1698431365
transform 1 0 47488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_420
timestamp 1698431365
transform 1 0 48384 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_437
timestamp 1698431365
transform 1 0 50288 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_453
timestamp 1698431365
transform 1 0 52080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698431365
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_559
timestamp 1698431365
transform 1 0 63952 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_575
timestamp 1698431365
transform 1 0 65744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_579
timestamp 1698431365
transform 1 0 66192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_36
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_44
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_61
timestamp 1698431365
transform 1 0 8176 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_90
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_98
timestamp 1698431365
transform 1 0 12320 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_102
timestamp 1698431365
transform 1 0 12768 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_119
timestamp 1698431365
transform 1 0 14672 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_164
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_180
timestamp 1698431365
transform 1 0 21504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_198
timestamp 1698431365
transform 1 0 23520 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_202
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_228
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_265
timestamp 1698431365
transform 1 0 31024 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698431365
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_302
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_318
timestamp 1698431365
transform 1 0 36960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_336
timestamp 1698431365
transform 1 0 38976 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_344
timestamp 1698431365
transform 1 0 39872 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_377
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_385
timestamp 1698431365
transform 1 0 44464 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_402
timestamp 1698431365
transform 1 0 46368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_404
timestamp 1698431365
transform 1 0 46592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_411
timestamp 1698431365
transform 1 0 47376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_413
timestamp 1698431365
transform 1 0 47600 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_430
timestamp 1698431365
transform 1 0 49504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_434
timestamp 1698431365
transform 1 0 49952 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_451
timestamp 1698431365
transform 1 0 51856 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_483
timestamp 1698431365
transform 1 0 55440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_487
timestamp 1698431365
transform 1 0 55888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1698431365
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_578
timestamp 1698431365
transform 1 0 66080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_580
timestamp 1698431365
transform 1 0 66304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_77
timestamp 1698431365
transform 1 0 9968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_79
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_96
timestamp 1698431365
transform 1 0 12096 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698431365
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_141
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_149
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_166
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_170
timestamp 1698431365
transform 1 0 20384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_181
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_188
timestamp 1698431365
transform 1 0 22400 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_227
timestamp 1698431365
transform 1 0 26768 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_268
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_284
timestamp 1698431365
transform 1 0 33152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_302
timestamp 1698431365
transform 1 0 35168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_345
timestamp 1698431365
transform 1 0 39984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_357
timestamp 1698431365
transform 1 0 41328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_380
timestamp 1698431365
transform 1 0 43904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_382
timestamp 1698431365
transform 1 0 44128 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_391
timestamp 1698431365
transform 1 0 45136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_412
timestamp 1698431365
transform 1 0 47488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_420
timestamp 1698431365
transform 1 0 48384 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_437
timestamp 1698431365
transform 1 0 50288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_439
timestamp 1698431365
transform 1 0 50512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_446
timestamp 1698431365
transform 1 0 51296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1698431365
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_465
timestamp 1698431365
transform 1 0 53424 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_485
timestamp 1698431365
transform 1 0 55664 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_517
timestamp 1698431365
transform 1 0 59248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_559
timestamp 1698431365
transform 1 0 63952 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_575
timestamp 1698431365
transform 1 0 65744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_579
timestamp 1698431365
transform 1 0 66192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_22
timestamp 1698431365
transform 1 0 3808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_89
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_97
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_124
timestamp 1698431365
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_128
timestamp 1698431365
transform 1 0 15680 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_132
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_192
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_202
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_217
timestamp 1698431365
transform 1 0 25648 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_234
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_242
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_246
timestamp 1698431365
transform 1 0 28896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_248
timestamp 1698431365
transform 1 0 29120 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_298
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_332
timestamp 1698431365
transform 1 0 38528 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_348
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_360
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_426
timestamp 1698431365
transform 1 0 49056 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_430
timestamp 1698431365
transform 1 0 49504 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_447
timestamp 1698431365
transform 1 0 51408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_455
timestamp 1698431365
transform 1 0 52304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_478
timestamp 1698431365
transform 1 0 54880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698431365
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_578
timestamp 1698431365
transform 1 0 66080 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_580
timestamp 1698431365
transform 1 0 66304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_57
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_60
timestamp 1698431365
transform 1 0 8064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_96
timestamp 1698431365
transform 1 0 12096 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_113
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_121
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_197
timestamp 1698431365
transform 1 0 23408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_199
timestamp 1698431365
transform 1 0 23632 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_236
timestamp 1698431365
transform 1 0 27776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_267
timestamp 1698431365
transform 1 0 31248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_303
timestamp 1698431365
transform 1 0 35280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_323
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_331
timestamp 1698431365
transform 1 0 38416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_333
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_350
timestamp 1698431365
transform 1 0 40544 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_358
timestamp 1698431365
transform 1 0 41440 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_362
timestamp 1698431365
transform 1 0 41888 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_421
timestamp 1698431365
transform 1 0 48496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_425
timestamp 1698431365
transform 1 0 48944 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_428
timestamp 1698431365
transform 1 0 49280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_452
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_465
timestamp 1698431365
transform 1 0 53424 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_482
timestamp 1698431365
transform 1 0 55328 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_514
timestamp 1698431365
transform 1 0 58912 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_522
timestamp 1698431365
transform 1 0 59808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_524
timestamp 1698431365
transform 1 0 60032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_559
timestamp 1698431365
transform 1 0 63952 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_575
timestamp 1698431365
transform 1 0 65744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_579
timestamp 1698431365
transform 1 0 66192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_27
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_35
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_168
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_204
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_225
timestamp 1698431365
transform 1 0 26544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_229
timestamp 1698431365
transform 1 0 26992 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_233
timestamp 1698431365
transform 1 0 27440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698431365
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_341
timestamp 1698431365
transform 1 0 39536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_345
timestamp 1698431365
transform 1 0 39984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_358
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_393
timestamp 1698431365
transform 1 0 45360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_397
timestamp 1698431365
transform 1 0 45808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_401
timestamp 1698431365
transform 1 0 46256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_418
timestamp 1698431365
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_458
timestamp 1698431365
transform 1 0 52640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_462
timestamp 1698431365
transform 1 0 53088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_466
timestamp 1698431365
transform 1 0 53536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_489
timestamp 1698431365
transform 1 0 56112 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_500
timestamp 1698431365
transform 1 0 57344 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_517
timestamp 1698431365
transform 1 0 59248 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_549
timestamp 1698431365
transform 1 0 62832 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_557
timestamp 1698431365
transform 1 0 63728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_559
timestamp 1698431365
transform 1 0 63952 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_578
timestamp 1698431365
transform 1 0 66080 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_580
timestamp 1698431365
transform 1 0 66304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_231
timestamp 1698431365
transform 1 0 27216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698431365
transform 1 0 27664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_273
timestamp 1698431365
transform 1 0 31920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_491
timestamp 1698431365
transform 1 0 56336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_499
timestamp 1698431365
transform 1 0 57232 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_516
timestamp 1698431365
transform 1 0 59136 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_524
timestamp 1698431365
transform 1 0 60032 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_559
timestamp 1698431365
transform 1 0 63952 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_575
timestamp 1698431365
transform 1 0 65744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_579
timestamp 1698431365
transform 1 0 66192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_27
timestamp 1698431365
transform 1 0 4368 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_35
timestamp 1698431365
transform 1 0 5264 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_356
timestamp 1698431365
transform 1 0 41216 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_418
timestamp 1698431365
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_500
timestamp 1698431365
transform 1 0 57344 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_523
timestamp 1698431365
transform 1 0 59920 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_555
timestamp 1698431365
transform 1 0 63504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_559
timestamp 1698431365
transform 1 0 63952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_578
timestamp 1698431365
transform 1 0 66080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_580
timestamp 1698431365
transform 1 0 66304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_6
timestamp 1698431365
transform 1 0 2016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_39
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_88
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_163
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698431365
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_257
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_259
timestamp 1698431365
transform 1 0 30352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_266
timestamp 1698431365
transform 1 0 31136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_425
timestamp 1698431365
transform 1 0 48944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_429
timestamp 1698431365
transform 1 0 49392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_433
timestamp 1698431365
transform 1 0 49840 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_450
timestamp 1698431365
transform 1 0 51744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_454
timestamp 1698431365
transform 1 0 52192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_513
timestamp 1698431365
transform 1 0 58800 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_559
timestamp 1698431365
transform 1 0 63952 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_575
timestamp 1698431365
transform 1 0 65744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_579
timestamp 1698431365
transform 1 0 66192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_155
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698431365
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_288
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_339
timestamp 1698431365
transform 1 0 39312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_440
timestamp 1698431365
transform 1 0 50624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_444
timestamp 1698431365
transform 1 0 51072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_485
timestamp 1698431365
transform 1 0 55664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_489
timestamp 1698431365
transform 1 0 56112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_500
timestamp 1698431365
transform 1 0 57344 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_517
timestamp 1698431365
transform 1 0 59248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_525
timestamp 1698431365
transform 1 0 60144 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_542
timestamp 1698431365
transform 1 0 62048 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_558
timestamp 1698431365
transform 1 0 63840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_578
timestamp 1698431365
transform 1 0 66080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_580
timestamp 1698431365
transform 1 0 66304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_59
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_64
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_102
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_111
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_117
timestamp 1698431365
transform 1 0 14448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_200
timestamp 1698431365
transform 1 0 23744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_204
timestamp 1698431365
transform 1 0 24192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_206
timestamp 1698431365
transform 1 0 24416 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_253
timestamp 1698431365
transform 1 0 29680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_262
timestamp 1698431365
transform 1 0 30688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_266
timestamp 1698431365
transform 1 0 31136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_302
timestamp 1698431365
transform 1 0 35168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_391
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_493
timestamp 1698431365
transform 1 0 56560 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_501
timestamp 1698431365
transform 1 0 57456 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_524
timestamp 1698431365
transform 1 0 60032 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_559
timestamp 1698431365
transform 1 0 63952 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_575
timestamp 1698431365
transform 1 0 65744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_579
timestamp 1698431365
transform 1 0 66192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_19
timestamp 1698431365
transform 1 0 3472 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_27
timestamp 1698431365
transform 1 0 4368 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_78
timestamp 1698431365
transform 1 0 10080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_92
timestamp 1698431365
transform 1 0 11648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_130
timestamp 1698431365
transform 1 0 15904 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_356
timestamp 1698431365
transform 1 0 41216 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_417
timestamp 1698431365
transform 1 0 48048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_456
timestamp 1698431365
transform 1 0 52416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_460
timestamp 1698431365
transform 1 0 52864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_464
timestamp 1698431365
transform 1 0 53312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_487
timestamp 1698431365
transform 1 0 55888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_489
timestamp 1698431365
transform 1 0 56112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_500
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_517
timestamp 1698431365
transform 1 0 59248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_525
timestamp 1698431365
transform 1 0 60144 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_542
timestamp 1698431365
transform 1 0 62048 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_558
timestamp 1698431365
transform 1 0 63840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_578
timestamp 1698431365
transform 1 0 66080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_580
timestamp 1698431365
transform 1 0 66304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_227
timestamp 1698431365
transform 1 0 26768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_231
timestamp 1698431365
transform 1 0 27216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_235
timestamp 1698431365
transform 1 0 27664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_281
timestamp 1698431365
transform 1 0 32816 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_289
timestamp 1698431365
transform 1 0 33712 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_453
timestamp 1698431365
transform 1 0 52080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_491
timestamp 1698431365
transform 1 0 56336 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_499
timestamp 1698431365
transform 1 0 57232 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_522
timestamp 1698431365
transform 1 0 59808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_524
timestamp 1698431365
transform 1 0 60032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_535
timestamp 1698431365
transform 1 0 61264 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_552
timestamp 1698431365
transform 1 0 63168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_568
timestamp 1698431365
transform 1 0 64960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_576
timestamp 1698431365
transform 1 0 65856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_580
timestamp 1698431365
transform 1 0 66304 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_87
timestamp 1698431365
transform 1 0 11088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_128
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_132
timestamp 1698431365
transform 1 0 16128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_155
timestamp 1698431365
transform 1 0 18704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_159
timestamp 1698431365
transform 1 0 19152 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_162
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_228
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_230
timestamp 1698431365
transform 1 0 27104 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_267
timestamp 1698431365
transform 1 0 31248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_286
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_333
timestamp 1698431365
transform 1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_432
timestamp 1698431365
transform 1 0 49728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_468
timestamp 1698431365
transform 1 0 53760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_470
timestamp 1698431365
transform 1 0 53984 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_483
timestamp 1698431365
transform 1 0 55440 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_496
timestamp 1698431365
transform 1 0 56896 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_500
timestamp 1698431365
transform 1 0 57344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_517
timestamp 1698431365
transform 1 0 59248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_525
timestamp 1698431365
transform 1 0 60144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_542
timestamp 1698431365
transform 1 0 62048 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_558
timestamp 1698431365
transform 1 0 63840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_578
timestamp 1698431365
transform 1 0 66080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_580
timestamp 1698431365
transform 1 0 66304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_26
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_30
timestamp 1698431365
transform 1 0 4704 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_94
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_96
timestamp 1698431365
transform 1 0 12096 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_139
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_251
timestamp 1698431365
transform 1 0 29456 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_304
timestamp 1698431365
transform 1 0 35392 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_308
timestamp 1698431365
transform 1 0 35840 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_454
timestamp 1698431365
transform 1 0 52192 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_491
timestamp 1698431365
transform 1 0 56336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_495
timestamp 1698431365
transform 1 0 56784 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_499
timestamp 1698431365
transform 1 0 57232 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_522
timestamp 1698431365
transform 1 0 59808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_524
timestamp 1698431365
transform 1 0 60032 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_535
timestamp 1698431365
transform 1 0 61264 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_552
timestamp 1698431365
transform 1 0 63168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_568
timestamp 1698431365
transform 1 0 64960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_576
timestamp 1698431365
transform 1 0 65856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_580
timestamp 1698431365
transform 1 0 66304 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_10
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_27
timestamp 1698431365
transform 1 0 4368 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_35
timestamp 1698431365
transform 1 0 5264 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_171
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_175
timestamp 1698431365
transform 1 0 20944 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_294
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_296
timestamp 1698431365
transform 1 0 34496 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_347
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_364
timestamp 1698431365
transform 1 0 42112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_399
timestamp 1698431365
transform 1 0 46032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_403
timestamp 1698431365
transform 1 0 46480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_407
timestamp 1698431365
transform 1 0 46928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_411
timestamp 1698431365
transform 1 0 47376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_413
timestamp 1698431365
transform 1 0 47600 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_496
timestamp 1698431365
transform 1 0 56896 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_500
timestamp 1698431365
transform 1 0 57344 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_517
timestamp 1698431365
transform 1 0 59248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_525
timestamp 1698431365
transform 1 0 60144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_542
timestamp 1698431365
transform 1 0 62048 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_558
timestamp 1698431365
transform 1 0 63840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_578
timestamp 1698431365
transform 1 0 66080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_580
timestamp 1698431365
transform 1 0 66304 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_26
timestamp 1698431365
transform 1 0 4256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_30
timestamp 1698431365
transform 1 0 4704 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_55
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_58
timestamp 1698431365
transform 1 0 7840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_102
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_161
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_165
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_192
timestamp 1698431365
transform 1 0 22848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_196
timestamp 1698431365
transform 1 0 23296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_238
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_443
timestamp 1698431365
transform 1 0 50960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_447
timestamp 1698431365
transform 1 0 51408 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_514
timestamp 1698431365
transform 1 0 58912 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_522
timestamp 1698431365
transform 1 0 59808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_524
timestamp 1698431365
transform 1 0 60032 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_535
timestamp 1698431365
transform 1 0 61264 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_552
timestamp 1698431365
transform 1 0 63168 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_568
timestamp 1698431365
transform 1 0 64960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_576
timestamp 1698431365
transform 1 0 65856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_580
timestamp 1698431365
transform 1 0 66304 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_26
timestamp 1698431365
transform 1 0 4256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_61
timestamp 1698431365
transform 1 0 8176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_63
timestamp 1698431365
transform 1 0 8400 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_144
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_151
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_155
timestamp 1698431365
transform 1 0 18704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_196
timestamp 1698431365
transform 1 0 23296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_200
timestamp 1698431365
transform 1 0 23744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_204
timestamp 1698431365
transform 1 0 24192 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_208
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_216
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_348
timestamp 1698431365
transform 1 0 40320 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_526
timestamp 1698431365
transform 1 0 60256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_530
timestamp 1698431365
transform 1 0 60704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_534
timestamp 1698431365
transform 1 0 61152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_551
timestamp 1698431365
transform 1 0 63056 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_559
timestamp 1698431365
transform 1 0 63952 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_566
timestamp 1698431365
transform 1 0 64736 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_26
timestamp 1698431365
transform 1 0 4256 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_62
timestamp 1698431365
transform 1 0 8288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_66
timestamp 1698431365
transform 1 0 8736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_68
timestamp 1698431365
transform 1 0 8960 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_421
timestamp 1698431365
transform 1 0 48496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_425
timestamp 1698431365
transform 1 0 48944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_429
timestamp 1698431365
transform 1 0 49392 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_452
timestamp 1698431365
transform 1 0 51968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_491
timestamp 1698431365
transform 1 0 56336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_495
timestamp 1698431365
transform 1 0 56784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_499
timestamp 1698431365
transform 1 0 57232 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_516
timestamp 1698431365
transform 1 0 59136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_524
timestamp 1698431365
transform 1 0 60032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_535
timestamp 1698431365
transform 1 0 61264 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_552
timestamp 1698431365
transform 1 0 63168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_560
timestamp 1698431365
transform 1 0 64064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_577
timestamp 1698431365
transform 1 0 65968 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_18
timestamp 1698431365
transform 1 0 3360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_36
timestamp 1698431365
transform 1 0 5376 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_65
timestamp 1698431365
transform 1 0 8624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_133
timestamp 1698431365
transform 1 0 16240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_390
timestamp 1698431365
transform 1 0 45024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_394
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_398
timestamp 1698431365
transform 1 0 45920 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_415
timestamp 1698431365
transform 1 0 47824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_426
timestamp 1698431365
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_430
timestamp 1698431365
transform 1 0 49504 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_447
timestamp 1698431365
transform 1 0 51408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_451
timestamp 1698431365
transform 1 0 51856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_453
timestamp 1698431365
transform 1 0 52080 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_478
timestamp 1698431365
transform 1 0 54880 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_500
timestamp 1698431365
transform 1 0 57344 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_517
timestamp 1698431365
transform 1 0 59248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_525
timestamp 1698431365
transform 1 0 60144 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_542
timestamp 1698431365
transform 1 0 62048 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_558
timestamp 1698431365
transform 1 0 63840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_578
timestamp 1698431365
transform 1 0 66080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_580
timestamp 1698431365
transform 1 0 66304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_26
timestamp 1698431365
transform 1 0 4256 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_41
timestamp 1698431365
transform 1 0 5936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_43
timestamp 1698431365
transform 1 0 6160 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_60
timestamp 1698431365
transform 1 0 8064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_64
timestamp 1698431365
transform 1 0 8512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_66
timestamp 1698431365
transform 1 0 8736 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_103
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_183
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_194
timestamp 1698431365
transform 1 0 23072 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_299
timestamp 1698431365
transform 1 0 34832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_303
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_319
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_461
timestamp 1698431365
transform 1 0 52976 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_465
timestamp 1698431365
transform 1 0 53424 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_482
timestamp 1698431365
transform 1 0 55328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_490
timestamp 1698431365
transform 1 0 56224 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_507
timestamp 1698431365
transform 1 0 58128 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_523
timestamp 1698431365
transform 1 0 59920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_535
timestamp 1698431365
transform 1 0 61264 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_552
timestamp 1698431365
transform 1 0 63168 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_568
timestamp 1698431365
transform 1 0 64960 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_576
timestamp 1698431365
transform 1 0 65856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_580
timestamp 1698431365
transform 1 0 66304 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_18
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_36
timestamp 1698431365
transform 1 0 5376 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_44
timestamp 1698431365
transform 1 0 6272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_61
timestamp 1698431365
transform 1 0 8176 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_84
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_86
timestamp 1698431365
transform 1 0 10976 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_123
timestamp 1698431365
transform 1 0 15120 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_126
timestamp 1698431365
transform 1 0 15456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_130
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_392
timestamp 1698431365
transform 1 0 45248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_496
timestamp 1698431365
transform 1 0 56896 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_500
timestamp 1698431365
transform 1 0 57344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_517
timestamp 1698431365
transform 1 0 59248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_525
timestamp 1698431365
transform 1 0 60144 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_542
timestamp 1698431365
transform 1 0 62048 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_558
timestamp 1698431365
transform 1 0 63840 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_578
timestamp 1698431365
transform 1 0 66080 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_580
timestamp 1698431365
transform 1 0 66304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_26
timestamp 1698431365
transform 1 0 4256 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_55
timestamp 1698431365
transform 1 0 7504 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_63
timestamp 1698431365
transform 1 0 8400 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_98
timestamp 1698431365
transform 1 0 12320 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_253
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_306
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_310
timestamp 1698431365
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_323
timestamp 1698431365
transform 1 0 37520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_375
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_379
timestamp 1698431365
transform 1 0 43792 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_389
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_396
timestamp 1698431365
transform 1 0 45696 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_403
timestamp 1698431365
transform 1 0 46480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_447
timestamp 1698431365
transform 1 0 51408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_492
timestamp 1698431365
transform 1 0 56448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_496
timestamp 1698431365
transform 1 0 56896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_500
timestamp 1698431365
transform 1 0 57344 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_523
timestamp 1698431365
transform 1 0 59920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_535
timestamp 1698431365
transform 1 0 61264 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_552
timestamp 1698431365
transform 1 0 63168 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_568
timestamp 1698431365
transform 1 0 64960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_576
timestamp 1698431365
transform 1 0 65856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_580
timestamp 1698431365
transform 1 0 66304 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_6
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_36
timestamp 1698431365
transform 1 0 5376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_44
timestamp 1698431365
transform 1 0 6272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_61
timestamp 1698431365
transform 1 0 8176 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_148
timestamp 1698431365
transform 1 0 17920 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_155
timestamp 1698431365
transform 1 0 18704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_193
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_195
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_214
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_298
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_333
timestamp 1698431365
transform 1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_337
timestamp 1698431365
transform 1 0 39088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_345
timestamp 1698431365
transform 1 0 39984 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_426
timestamp 1698431365
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_430
timestamp 1698431365
transform 1 0 49504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_432
timestamp 1698431365
transform 1 0 49728 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_473
timestamp 1698431365
transform 1 0 54320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_475
timestamp 1698431365
transform 1 0 54544 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_488
timestamp 1698431365
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_496
timestamp 1698431365
transform 1 0 56896 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_500
timestamp 1698431365
transform 1 0 57344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_517
timestamp 1698431365
transform 1 0 59248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_525
timestamp 1698431365
transform 1 0 60144 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_542
timestamp 1698431365
transform 1 0 62048 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_558
timestamp 1698431365
transform 1 0 63840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_578
timestamp 1698431365
transform 1 0 66080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_580
timestamp 1698431365
transform 1 0 66304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_26
timestamp 1698431365
transform 1 0 4256 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_62
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_157
timestamp 1698431365
transform 1 0 18928 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_193
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_323
timestamp 1698431365
transform 1 0 37520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_361
timestamp 1698431365
transform 1 0 41776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_365
timestamp 1698431365
transform 1 0 42224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_369
timestamp 1698431365
transform 1 0 42672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_378
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_413
timestamp 1698431365
transform 1 0 47600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_415
timestamp 1698431365
transform 1 0 47824 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_450
timestamp 1698431365
transform 1 0 51744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_454
timestamp 1698431365
transform 1 0 52192 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_491
timestamp 1698431365
transform 1 0 56336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_495
timestamp 1698431365
transform 1 0 56784 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_499
timestamp 1698431365
transform 1 0 57232 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_516
timestamp 1698431365
transform 1 0 59136 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_524
timestamp 1698431365
transform 1 0 60032 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_535
timestamp 1698431365
transform 1 0 61264 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_552
timestamp 1698431365
transform 1 0 63168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_568
timestamp 1698431365
transform 1 0 64960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_576
timestamp 1698431365
transform 1 0 65856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_580
timestamp 1698431365
transform 1 0 66304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_36
timestamp 1698431365
transform 1 0 5376 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_61
timestamp 1698431365
transform 1 0 8176 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_97
timestamp 1698431365
transform 1 0 12208 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_105
timestamp 1698431365
transform 1 0 13104 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_288
timestamp 1698431365
transform 1 0 33600 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_340
timestamp 1698431365
transform 1 0 39424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_356
timestamp 1698431365
transform 1 0 41216 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_415
timestamp 1698431365
transform 1 0 47824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_417
timestamp 1698431365
transform 1 0 48048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_428
timestamp 1698431365
transform 1 0 49280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_432
timestamp 1698431365
transform 1 0 49728 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_480
timestamp 1698431365
transform 1 0 55104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_488
timestamp 1698431365
transform 1 0 56000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_496
timestamp 1698431365
transform 1 0 56896 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_500
timestamp 1698431365
transform 1 0 57344 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_517
timestamp 1698431365
transform 1 0 59248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_525
timestamp 1698431365
transform 1 0 60144 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_542
timestamp 1698431365
transform 1 0 62048 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_558
timestamp 1698431365
transform 1 0 63840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_578
timestamp 1698431365
transform 1 0 66080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_580
timestamp 1698431365
transform 1 0 66304 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_45
timestamp 1698431365
transform 1 0 6384 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_62
timestamp 1698431365
transform 1 0 8288 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_70
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_109
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_160
timestamp 1698431365
transform 1 0 19264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_162
timestamp 1698431365
transform 1 0 19488 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_197
timestamp 1698431365
transform 1 0 23408 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_201
timestamp 1698431365
transform 1 0 23856 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698431365
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_240
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_255
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_259
timestamp 1698431365
transform 1 0 30352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_261
timestamp 1698431365
transform 1 0 30576 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_302
timestamp 1698431365
transform 1 0 35168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_310
timestamp 1698431365
transform 1 0 36064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_335
timestamp 1698431365
transform 1 0 38864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_507
timestamp 1698431365
transform 1 0 58128 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_523
timestamp 1698431365
transform 1 0 59920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_535
timestamp 1698431365
transform 1 0 61264 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_552
timestamp 1698431365
transform 1 0 63168 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_568
timestamp 1698431365
transform 1 0 64960 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_576
timestamp 1698431365
transform 1 0 65856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_580
timestamp 1698431365
transform 1 0 66304 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_34
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_42
timestamp 1698431365
transform 1 0 6048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_44
timestamp 1698431365
transform 1 0 6272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_61
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_74
timestamp 1698431365
transform 1 0 9632 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_97
timestamp 1698431365
transform 1 0 12208 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_105
timestamp 1698431365
transform 1 0 13104 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_387
timestamp 1698431365
transform 1 0 44688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_391
timestamp 1698431365
transform 1 0 45136 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_395
timestamp 1698431365
transform 1 0 45584 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_428
timestamp 1698431365
transform 1 0 49280 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_464
timestamp 1698431365
transform 1 0 53312 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_470
timestamp 1698431365
transform 1 0 53984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_472
timestamp 1698431365
transform 1 0 54208 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_489
timestamp 1698431365
transform 1 0 56112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_496
timestamp 1698431365
transform 1 0 56896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_500
timestamp 1698431365
transform 1 0 57344 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_517
timestamp 1698431365
transform 1 0 59248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_525
timestamp 1698431365
transform 1 0 60144 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_542
timestamp 1698431365
transform 1 0 62048 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_558
timestamp 1698431365
transform 1 0 63840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_578
timestamp 1698431365
transform 1 0 66080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_580
timestamp 1698431365
transform 1 0 66304 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_53
timestamp 1698431365
transform 1 0 7280 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_71
timestamp 1698431365
transform 1 0 9296 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_79
timestamp 1698431365
transform 1 0 10192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_96
timestamp 1698431365
transform 1 0 12096 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_197
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_199
timestamp 1698431365
transform 1 0 23632 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_234
timestamp 1698431365
transform 1 0 27552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_236
timestamp 1698431365
transform 1 0 27776 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_303
timestamp 1698431365
transform 1 0 35280 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_321
timestamp 1698431365
transform 1 0 37296 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_324
timestamp 1698431365
transform 1 0 37632 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_359
timestamp 1698431365
transform 1 0 41552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_363
timestamp 1698431365
transform 1 0 42000 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_367
timestamp 1698431365
transform 1 0 42448 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_421
timestamp 1698431365
transform 1 0 48496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_425
timestamp 1698431365
transform 1 0 48944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_429
timestamp 1698431365
transform 1 0 49392 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_452
timestamp 1698431365
transform 1 0 51968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698431365
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_495
timestamp 1698431365
transform 1 0 56784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_499
timestamp 1698431365
transform 1 0 57232 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_503
timestamp 1698431365
transform 1 0 57680 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_520
timestamp 1698431365
transform 1 0 59584 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_524
timestamp 1698431365
transform 1 0 60032 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_527
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_535
timestamp 1698431365
transform 1 0 61264 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_552
timestamp 1698431365
transform 1 0 63168 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_568
timestamp 1698431365
transform 1 0 64960 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_576
timestamp 1698431365
transform 1 0 65856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_580
timestamp 1698431365
transform 1 0 66304 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_126
timestamp 1698431365
transform 1 0 15456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_130
timestamp 1698431365
transform 1 0 15904 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_137
timestamp 1698431365
transform 1 0 16688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_149
timestamp 1698431365
transform 1 0 18032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_167
timestamp 1698431365
transform 1 0 20048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_171
timestamp 1698431365
transform 1 0 20496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_175
timestamp 1698431365
transform 1 0 20944 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_214
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_237
timestamp 1698431365
transform 1 0 27888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_241
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_245
timestamp 1698431365
transform 1 0 28784 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_321
timestamp 1698431365
transform 1 0 37296 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_329
timestamp 1698431365
transform 1 0 38192 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_417
timestamp 1698431365
transform 1 0 48048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_448
timestamp 1698431365
transform 1 0 51520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_496
timestamp 1698431365
transform 1 0 56896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_500
timestamp 1698431365
transform 1 0 57344 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_517
timestamp 1698431365
transform 1 0 59248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_521
timestamp 1698431365
transform 1 0 59696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_525
timestamp 1698431365
transform 1 0 60144 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_542
timestamp 1698431365
transform 1 0 62048 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_558
timestamp 1698431365
transform 1 0 63840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_562
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_578
timestamp 1698431365
transform 1 0 66080 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_580
timestamp 1698431365
transform 1 0 66304 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_69
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_77
timestamp 1698431365
transform 1 0 9968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_79
timestamp 1698431365
transform 1 0 10192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_96
timestamp 1698431365
transform 1 0 12096 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_123
timestamp 1698431365
transform 1 0 15120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_141
timestamp 1698431365
transform 1 0 17136 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_149
timestamp 1698431365
transform 1 0 18032 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_166
timestamp 1698431365
transform 1 0 19936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_170
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_203
timestamp 1698431365
transform 1 0 24080 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_249
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_266
timestamp 1698431365
transform 1 0 31136 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_274
timestamp 1698431365
transform 1 0 32032 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_323
timestamp 1698431365
transform 1 0 37520 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_327
timestamp 1698431365
transform 1 0 37968 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_380
timestamp 1698431365
transform 1 0 43904 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_491
timestamp 1698431365
transform 1 0 56336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_495
timestamp 1698431365
transform 1 0 56784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_499
timestamp 1698431365
transform 1 0 57232 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_522
timestamp 1698431365
transform 1 0 59808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_524
timestamp 1698431365
transform 1 0 60032 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_527
timestamp 1698431365
transform 1 0 60368 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_535
timestamp 1698431365
transform 1 0 61264 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_552
timestamp 1698431365
transform 1 0 63168 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_568
timestamp 1698431365
transform 1 0 64960 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_576
timestamp 1698431365
transform 1 0 65856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_580
timestamp 1698431365
transform 1 0 66304 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_88
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_106
timestamp 1698431365
transform 1 0 13216 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_122
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_158
timestamp 1698431365
transform 1 0 19040 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_166
timestamp 1698431365
transform 1 0 19936 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_214
timestamp 1698431365
transform 1 0 25312 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_275
timestamp 1698431365
transform 1 0 32144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_496
timestamp 1698431365
transform 1 0 56896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_500
timestamp 1698431365
transform 1 0 57344 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_517
timestamp 1698431365
transform 1 0 59248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_521
timestamp 1698431365
transform 1 0 59696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_525
timestamp 1698431365
transform 1 0 60144 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_548
timestamp 1698431365
transform 1 0 62720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_552
timestamp 1698431365
transform 1 0 63168 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_562
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_578
timestamp 1698431365
transform 1 0 66080 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_580
timestamp 1698431365
transform 1 0 66304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_123
timestamp 1698431365
transform 1 0 15120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_141
timestamp 1698431365
transform 1 0 17136 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_145
timestamp 1698431365
transform 1 0 17584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_147
timestamp 1698431365
transform 1 0 17808 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_166
timestamp 1698431365
transform 1 0 19936 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_535
timestamp 1698431365
transform 1 0 61264 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_552
timestamp 1698431365
transform 1 0 63168 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_568
timestamp 1698431365
transform 1 0 64960 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_576
timestamp 1698431365
transform 1 0 65856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_580
timestamp 1698431365
transform 1 0 66304 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_104
timestamp 1698431365
transform 1 0 12992 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_112
timestamp 1698431365
transform 1 0 13888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_114
timestamp 1698431365
transform 1 0 14112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_131
timestamp 1698431365
transform 1 0 16016 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_164
timestamp 1698431365
transform 1 0 19712 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_172
timestamp 1698431365
transform 1 0 20608 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_228
timestamp 1698431365
transform 1 0 26880 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_232
timestamp 1698431365
transform 1 0 27328 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_234
timestamp 1698431365
transform 1 0 27552 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_271
timestamp 1698431365
transform 1 0 31696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_273
timestamp 1698431365
transform 1 0 31920 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_295
timestamp 1698431365
transform 1 0 34384 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_299
timestamp 1698431365
transform 1 0 34832 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_412
timestamp 1698431365
transform 1 0 47488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_438
timestamp 1698431365
transform 1 0 50400 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_440
timestamp 1698431365
transform 1 0 50624 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_483
timestamp 1698431365
transform 1 0 55440 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_496
timestamp 1698431365
transform 1 0 56896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_500
timestamp 1698431365
transform 1 0 57344 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_517
timestamp 1698431365
transform 1 0 59248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_521
timestamp 1698431365
transform 1 0 59696 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_525
timestamp 1698431365
transform 1 0 60144 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_542
timestamp 1698431365
transform 1 0 62048 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_558
timestamp 1698431365
transform 1 0 63840 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_578
timestamp 1698431365
transform 1 0 66080 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_580
timestamp 1698431365
transform 1 0 66304 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_135
timestamp 1698431365
transform 1 0 16464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_139
timestamp 1698431365
transform 1 0 16912 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_179
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_196
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_200
timestamp 1698431365
transform 1 0 23744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_202
timestamp 1698431365
transform 1 0 23968 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_249
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_256
timestamp 1698431365
transform 1 0 30016 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_263
timestamp 1698431365
transform 1 0 30800 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_267
timestamp 1698431365
transform 1 0 31248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_303
timestamp 1698431365
transform 1 0 35280 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_307
timestamp 1698431365
transform 1 0 35728 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_351
timestamp 1698431365
transform 1 0 40656 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_355
timestamp 1698431365
transform 1 0 41104 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_359
timestamp 1698431365
transform 1 0 41552 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_382
timestamp 1698431365
transform 1 0 44128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_389
timestamp 1698431365
transform 1 0 44912 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_396
timestamp 1698431365
transform 1 0 45696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_438
timestamp 1698431365
transform 1 0 50400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_442
timestamp 1698431365
transform 1 0 50848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_452
timestamp 1698431365
transform 1 0 51968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_519
timestamp 1698431365
transform 1 0 59472 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_523
timestamp 1698431365
transform 1 0 59920 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_535
timestamp 1698431365
transform 1 0 61264 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_552
timestamp 1698431365
transform 1 0 63168 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_568
timestamp 1698431365
transform 1 0 64960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_576
timestamp 1698431365
transform 1 0 65856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_580
timestamp 1698431365
transform 1 0 66304 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_164
timestamp 1698431365
transform 1 0 19712 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_172
timestamp 1698431365
transform 1 0 20608 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_207
timestamp 1698431365
transform 1 0 24528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_262
timestamp 1698431365
transform 1 0 30688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_266
timestamp 1698431365
transform 1 0 31136 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_356
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_363
timestamp 1698431365
transform 1 0 42000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_365
timestamp 1698431365
transform 1 0 42224 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_400
timestamp 1698431365
transform 1 0 46144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_414
timestamp 1698431365
transform 1 0 47712 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_496
timestamp 1698431365
transform 1 0 56896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_500
timestamp 1698431365
transform 1 0 57344 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_517
timestamp 1698431365
transform 1 0 59248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_521
timestamp 1698431365
transform 1 0 59696 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_525
timestamp 1698431365
transform 1 0 60144 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_542
timestamp 1698431365
transform 1 0 62048 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_558
timestamp 1698431365
transform 1 0 63840 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_578
timestamp 1698431365
transform 1 0 66080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_580
timestamp 1698431365
transform 1 0 66304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_139
timestamp 1698431365
transform 1 0 16912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_321
timestamp 1698431365
transform 1 0 37296 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_382
timestamp 1698431365
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_391
timestamp 1698431365
transform 1 0 45136 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_395
timestamp 1698431365
transform 1 0 45584 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_448
timestamp 1698431365
transform 1 0 51520 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_452
timestamp 1698431365
transform 1 0 51968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_454
timestamp 1698431365
transform 1 0 52192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_491
timestamp 1698431365
transform 1 0 56336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_495
timestamp 1698431365
transform 1 0 56784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_499
timestamp 1698431365
transform 1 0 57232 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_522
timestamp 1698431365
transform 1 0 59808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_524
timestamp 1698431365
transform 1 0 60032 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_527
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_531
timestamp 1698431365
transform 1 0 60816 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_563
timestamp 1698431365
transform 1 0 64400 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_579
timestamp 1698431365
transform 1 0 66192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_160
timestamp 1698431365
transform 1 0 19264 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_168
timestamp 1698431365
transform 1 0 20160 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_172
timestamp 1698431365
transform 1 0 20608 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_207
timestamp 1698431365
transform 1 0 24528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698431365
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_228
timestamp 1698431365
transform 1 0 26880 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_236
timestamp 1698431365
transform 1 0 27776 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_271
timestamp 1698431365
transform 1 0 31696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_273
timestamp 1698431365
transform 1 0 31920 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_341
timestamp 1698431365
transform 1 0 39536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_343
timestamp 1698431365
transform 1 0 39760 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_496
timestamp 1698431365
transform 1 0 56896 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_500
timestamp 1698431365
transform 1 0 57344 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_523
timestamp 1698431365
transform 1 0 59920 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_555
timestamp 1698431365
transform 1 0 63504 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_559
timestamp 1698431365
transform 1 0 63952 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_562
timestamp 1698431365
transform 1 0 64288 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_578
timestamp 1698431365
transform 1 0 66080 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_580
timestamp 1698431365
transform 1 0 66304 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_139
timestamp 1698431365
transform 1 0 16912 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_147
timestamp 1698431365
transform 1 0 17808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_149
timestamp 1698431365
transform 1 0 18032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_166
timestamp 1698431365
transform 1 0 19936 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_174
timestamp 1698431365
transform 1 0 20832 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_179
timestamp 1698431365
transform 1 0 21392 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_186
timestamp 1698431365
transform 1 0 22176 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_190
timestamp 1698431365
transform 1 0 22624 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_194
timestamp 1698431365
transform 1 0 23072 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_369
timestamp 1698431365
transform 1 0 42672 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_373
timestamp 1698431365
transform 1 0 43120 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_491
timestamp 1698431365
transform 1 0 56336 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_495
timestamp 1698431365
transform 1 0 56784 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_499
timestamp 1698431365
transform 1 0 57232 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_516
timestamp 1698431365
transform 1 0 59136 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_520
timestamp 1698431365
transform 1 0 59584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_524
timestamp 1698431365
transform 1 0 60032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_527
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_559
timestamp 1698431365
transform 1 0 63952 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_575
timestamp 1698431365
transform 1 0 65744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_579
timestamp 1698431365
transform 1 0 66192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_158
timestamp 1698431365
transform 1 0 19040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_176
timestamp 1698431365
transform 1 0 21056 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_184
timestamp 1698431365
transform 1 0 21952 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_201
timestamp 1698431365
transform 1 0 23856 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698431365
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_256
timestamp 1698431365
transform 1 0 30016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_260
timestamp 1698431365
transform 1 0 30464 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_267
timestamp 1698431365
transform 1 0 31248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_275
timestamp 1698431365
transform 1 0 32144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_277
timestamp 1698431365
transform 1 0 32368 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_314
timestamp 1698431365
transform 1 0 36512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_358
timestamp 1698431365
transform 1 0 41440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_456
timestamp 1698431365
transform 1 0 52416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_460
timestamp 1698431365
transform 1 0 52864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_464
timestamp 1698431365
transform 1 0 53312 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_487
timestamp 1698431365
transform 1 0 55888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_489
timestamp 1698431365
transform 1 0 56112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_500
timestamp 1698431365
transform 1 0 57344 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_517
timestamp 1698431365
transform 1 0 59248 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_549
timestamp 1698431365
transform 1 0 62832 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_557
timestamp 1698431365
transform 1 0 63728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_559
timestamp 1698431365
transform 1 0 63952 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_562
timestamp 1698431365
transform 1 0 64288 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_578
timestamp 1698431365
transform 1 0 66080 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_580
timestamp 1698431365
transform 1 0 66304 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_139
timestamp 1698431365
transform 1 0 16912 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_147
timestamp 1698431365
transform 1 0 17808 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_149
timestamp 1698431365
transform 1 0 18032 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_166
timestamp 1698431365
transform 1 0 19936 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698431365
transform 1 0 20832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_194
timestamp 1698431365
transform 1 0 23072 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_202
timestamp 1698431365
transform 1 0 23968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_260
timestamp 1698431365
transform 1 0 30464 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_268
timestamp 1698431365
transform 1 0 31360 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_303
timestamp 1698431365
transform 1 0 35280 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_307
timestamp 1698431365
transform 1 0 35728 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_325
timestamp 1698431365
transform 1 0 37744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_379
timestamp 1698431365
transform 1 0 43792 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_383
timestamp 1698431365
transform 1 0 44240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_423
timestamp 1698431365
transform 1 0 48720 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_431
timestamp 1698431365
transform 1 0 49616 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_454
timestamp 1698431365
transform 1 0 52192 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_461
timestamp 1698431365
transform 1 0 52976 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_465
timestamp 1698431365
transform 1 0 53424 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_482
timestamp 1698431365
transform 1 0 55328 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_486
timestamp 1698431365
transform 1 0 55776 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_490
timestamp 1698431365
transform 1 0 56224 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_507
timestamp 1698431365
transform 1 0 58128 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_523
timestamp 1698431365
transform 1 0 59920 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_527
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_559
timestamp 1698431365
transform 1 0 63952 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_575
timestamp 1698431365
transform 1 0 65744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_579
timestamp 1698431365
transform 1 0 66192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_174
timestamp 1698431365
transform 1 0 20832 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_182
timestamp 1698431365
transform 1 0 21728 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_186
timestamp 1698431365
transform 1 0 22176 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_204
timestamp 1698431365
transform 1 0 24192 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_208
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_218
timestamp 1698431365
transform 1 0 25760 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_222
timestamp 1698431365
transform 1 0 26208 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_230
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_234
timestamp 1698431365
transform 1 0 27552 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_238
timestamp 1698431365
transform 1 0 28000 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_255
timestamp 1698431365
transform 1 0 29904 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_263
timestamp 1698431365
transform 1 0 30800 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_290
timestamp 1698431365
transform 1 0 33824 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_307
timestamp 1698431365
transform 1 0 35728 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_315
timestamp 1698431365
transform 1 0 36624 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_332
timestamp 1698431365
transform 1 0 38528 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_348
timestamp 1698431365
transform 1 0 40320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_360
timestamp 1698431365
transform 1 0 41664 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_364
timestamp 1698431365
transform 1 0 42112 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_417
timestamp 1698431365
transform 1 0 48048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1698431365
transform 1 0 48272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_426
timestamp 1698431365
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_476
timestamp 1698431365
transform 1 0 54656 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_480
timestamp 1698431365
transform 1 0 55104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_484
timestamp 1698431365
transform 1 0 55552 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_488
timestamp 1698431365
transform 1 0 56000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_500
timestamp 1698431365
transform 1 0 57344 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_517
timestamp 1698431365
transform 1 0 59248 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_549
timestamp 1698431365
transform 1 0 62832 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_557
timestamp 1698431365
transform 1 0 63728 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_559
timestamp 1698431365
transform 1 0 63952 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_562
timestamp 1698431365
transform 1 0 64288 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_578
timestamp 1698431365
transform 1 0 66080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_580
timestamp 1698431365
transform 1 0 66304 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_193
timestamp 1698431365
transform 1 0 22960 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_201
timestamp 1698431365
transform 1 0 23856 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_203
timestamp 1698431365
transform 1 0 24080 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_236
timestamp 1698431365
transform 1 0 27776 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_263
timestamp 1698431365
transform 1 0 30800 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_271
timestamp 1698431365
transform 1 0 31696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_275
timestamp 1698431365
transform 1 0 32144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_277
timestamp 1698431365
transform 1 0 32368 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_294
timestamp 1698431365
transform 1 0 34272 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_310
timestamp 1698431365
transform 1 0 36064 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_349
timestamp 1698431365
transform 1 0 40432 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_365
timestamp 1698431365
transform 1 0 42224 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_383
timestamp 1698431365
transform 1 0 44240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_395
timestamp 1698431365
transform 1 0 45584 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_412
timestamp 1698431365
transform 1 0 47488 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_420
timestamp 1698431365
transform 1 0 48384 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_437
timestamp 1698431365
transform 1 0 50288 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_453
timestamp 1698431365
transform 1 0 52080 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_465
timestamp 1698431365
transform 1 0 53424 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_485
timestamp 1698431365
transform 1 0 55664 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_493
timestamp 1698431365
transform 1 0 56560 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_510
timestamp 1698431365
transform 1 0 58464 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_518
timestamp 1698431365
transform 1 0 59360 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_522
timestamp 1698431365
transform 1 0 59808 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_524
timestamp 1698431365
transform 1 0 60032 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_559
timestamp 1698431365
transform 1 0 63952 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_575
timestamp 1698431365
transform 1 0 65744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_579
timestamp 1698431365
transform 1 0 66192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_174
timestamp 1698431365
transform 1 0 20832 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_182
timestamp 1698431365
transform 1 0 21728 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_202
timestamp 1698431365
transform 1 0 23968 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_228
timestamp 1698431365
transform 1 0 26880 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_261
timestamp 1698431365
transform 1 0 30576 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_277
timestamp 1698431365
transform 1 0 32368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1698431365
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_314
timestamp 1698431365
transform 1 0 36512 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_331
timestamp 1698431365
transform 1 0 38416 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_360
timestamp 1698431365
transform 1 0 41664 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_377
timestamp 1698431365
transform 1 0 43568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_385
timestamp 1698431365
transform 1 0 44464 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_402
timestamp 1698431365
transform 1 0 46368 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_418
timestamp 1698431365
transform 1 0 48160 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_430
timestamp 1698431365
transform 1 0 49504 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_447
timestamp 1698431365
transform 1 0 51408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_455
timestamp 1698431365
transform 1 0 52304 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_472
timestamp 1698431365
transform 1 0 54208 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_488
timestamp 1698431365
transform 1 0 56000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698431365
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_562
timestamp 1698431365
transform 1 0 64288 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_578
timestamp 1698431365
transform 1 0 66080 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_580
timestamp 1698431365
transform 1 0 66304 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_209
timestamp 1698431365
transform 1 0 24752 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_225
timestamp 1698431365
transform 1 0 26544 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_259
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_276
timestamp 1698431365
transform 1 0 32256 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_292
timestamp 1698431365
transform 1 0 34048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_310
timestamp 1698431365
transform 1 0 36064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_342
timestamp 1698431365
transform 1 0 39648 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_350
timestamp 1698431365
transform 1 0 40544 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_367
timestamp 1698431365
transform 1 0 42448 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_383
timestamp 1698431365
transform 1 0 44240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_395
timestamp 1698431365
transform 1 0 45584 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_412
timestamp 1698431365
transform 1 0 47488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_420
timestamp 1698431365
transform 1 0 48384 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_437
timestamp 1698431365
transform 1 0 50288 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_453
timestamp 1698431365
transform 1 0 52080 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_559
timestamp 1698431365
transform 1 0 63952 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_575
timestamp 1698431365
transform 1 0 65744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_579
timestamp 1698431365
transform 1 0 66192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_244
timestamp 1698431365
transform 1 0 28672 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_260
timestamp 1698431365
transform 1 0 30464 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_314
timestamp 1698431365
transform 1 0 36512 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_322
timestamp 1698431365
transform 1 0 37408 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_339
timestamp 1698431365
transform 1 0 39312 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_347
timestamp 1698431365
transform 1 0 40208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_370
timestamp 1698431365
transform 1 0 42784 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_386
timestamp 1698431365
transform 1 0 44576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_404
timestamp 1698431365
transform 1 0 46592 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_430
timestamp 1698431365
transform 1 0 49504 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_450
timestamp 1698431365
transform 1 0 51744 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_482
timestamp 1698431365
transform 1 0 55328 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698431365
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_562
timestamp 1698431365
transform 1 0 64288 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_578
timestamp 1698431365
transform 1 0 66080 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_580
timestamp 1698431365
transform 1 0 66304 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_255
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_257
timestamp 1698431365
transform 1 0 30128 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_274
timestamp 1698431365
transform 1 0 32032 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_282
timestamp 1698431365
transform 1 0 32928 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_286
timestamp 1698431365
transform 1 0 33376 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_303
timestamp 1698431365
transform 1 0 35280 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_347
timestamp 1698431365
transform 1 0 40208 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_355
timestamp 1698431365
transform 1 0 41104 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_372
timestamp 1698431365
transform 1 0 43008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_380
timestamp 1698431365
transform 1 0 43904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698431365
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_395
timestamp 1698431365
transform 1 0 45584 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_412
timestamp 1698431365
transform 1 0 47488 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_444
timestamp 1698431365
transform 1 0 51072 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_452
timestamp 1698431365
transform 1 0 51968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698431365
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_559
timestamp 1698431365
transform 1 0 63952 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_575
timestamp 1698431365
transform 1 0 65744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_579
timestamp 1698431365
transform 1 0 66192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_384
timestamp 1698431365
transform 1 0 44352 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698431365
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_562
timestamp 1698431365
transform 1 0 64288 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_578
timestamp 1698431365
transform 1 0 66080 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_580
timestamp 1698431365
transform 1 0 66304 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698431365
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_521
timestamp 1698431365
transform 1 0 59696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_527
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_559
timestamp 1698431365
transform 1 0 63952 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_575
timestamp 1698431365
transform 1 0 65744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_579
timestamp 1698431365
transform 1 0 66192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_66
timestamp 1698431365
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_136
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_276
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_416
timestamp 1698431365
transform 1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_422
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_556
timestamp 1698431365
transform 1 0 63616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_562
timestamp 1698431365
transform 1 0 64288 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_578
timestamp 1698431365
transform 1 0 66080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_580
timestamp 1698431365
transform 1 0 66304 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_171
timestamp 1698431365
transform 1 0 20496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_241
timestamp 1698431365
transform 1 0 28336 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_311
timestamp 1698431365
transform 1 0 36176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_381
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_451
timestamp 1698431365
transform 1 0 51856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_521
timestamp 1698431365
transform 1 0 59696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_527
timestamp 1698431365
transform 1 0 60368 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_559
timestamp 1698431365
transform 1 0 63952 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_575
timestamp 1698431365
transform 1 0 65744 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_579
timestamp 1698431365
transform 1 0 66192 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1698431365
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_136
timestamp 1698431365
transform 1 0 16576 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_206
timestamp 1698431365
transform 1 0 24416 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_276
timestamp 1698431365
transform 1 0 32256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_416
timestamp 1698431365
transform 1 0 47936 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_486
timestamp 1698431365
transform 1 0 55776 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_556
timestamp 1698431365
transform 1 0 63616 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_562
timestamp 1698431365
transform 1 0 64288 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_578
timestamp 1698431365
transform 1 0 66080 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_580
timestamp 1698431365
transform 1 0 66304 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1698431365
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_311
timestamp 1698431365
transform 1 0 36176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_451
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_521
timestamp 1698431365
transform 1 0 59696 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_527
timestamp 1698431365
transform 1 0 60368 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_559
timestamp 1698431365
transform 1 0 63952 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_575
timestamp 1698431365
transform 1 0 65744 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_579
timestamp 1698431365
transform 1 0 66192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_66
timestamp 1698431365
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_206
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_276
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_346
timestamp 1698431365
transform 1 0 40096 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_422
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_486
timestamp 1698431365
transform 1 0 55776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_556
timestamp 1698431365
transform 1 0 63616 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_562
timestamp 1698431365
transform 1 0 64288 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_578
timestamp 1698431365
transform 1 0 66080 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_580
timestamp 1698431365
transform 1 0 66304 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_171
timestamp 1698431365
transform 1 0 20496 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_241
timestamp 1698431365
transform 1 0 28336 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_311
timestamp 1698431365
transform 1 0 36176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_381
timestamp 1698431365
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_451
timestamp 1698431365
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_521
timestamp 1698431365
transform 1 0 59696 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_527
timestamp 1698431365
transform 1 0 60368 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_559
timestamp 1698431365
transform 1 0 63952 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_575
timestamp 1698431365
transform 1 0 65744 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_579
timestamp 1698431365
transform 1 0 66192 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_66
timestamp 1698431365
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_206
timestamp 1698431365
transform 1 0 24416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_276
timestamp 1698431365
transform 1 0 32256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_282
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_346
timestamp 1698431365
transform 1 0 40096 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_416
timestamp 1698431365
transform 1 0 47936 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_422
timestamp 1698431365
transform 1 0 48608 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_486
timestamp 1698431365
transform 1 0 55776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_492
timestamp 1698431365
transform 1 0 56448 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_556
timestamp 1698431365
transform 1 0 63616 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_562
timestamp 1698431365
transform 1 0 64288 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_578
timestamp 1698431365
transform 1 0 66080 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_580
timestamp 1698431365
transform 1 0 66304 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_171
timestamp 1698431365
transform 1 0 20496 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_241
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_381
timestamp 1698431365
transform 1 0 44016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_451
timestamp 1698431365
transform 1 0 51856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_457
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_521
timestamp 1698431365
transform 1 0 59696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_527
timestamp 1698431365
transform 1 0 60368 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_559
timestamp 1698431365
transform 1 0 63952 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_575
timestamp 1698431365
transform 1 0 65744 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_579
timestamp 1698431365
transform 1 0 66192 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_66
timestamp 1698431365
transform 1 0 8736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_276
timestamp 1698431365
transform 1 0 32256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_346
timestamp 1698431365
transform 1 0 40096 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_416
timestamp 1698431365
transform 1 0 47936 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_422
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_486
timestamp 1698431365
transform 1 0 55776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_492
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_556
timestamp 1698431365
transform 1 0 63616 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_562
timestamp 1698431365
transform 1 0 64288 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_578
timestamp 1698431365
transform 1 0 66080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_580
timestamp 1698431365
transform 1 0 66304 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_101
timestamp 1698431365
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698431365
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_381
timestamp 1698431365
transform 1 0 44016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_451
timestamp 1698431365
transform 1 0 51856 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_521
timestamp 1698431365
transform 1 0 59696 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_527
timestamp 1698431365
transform 1 0 60368 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_559
timestamp 1698431365
transform 1 0 63952 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_575
timestamp 1698431365
transform 1 0 65744 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_36
timestamp 1698431365
transform 1 0 5376 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_70
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_104
timestamp 1698431365
transform 1 0 12992 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_138
timestamp 1698431365
transform 1 0 16800 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_172
timestamp 1698431365
transform 1 0 20608 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_206
timestamp 1698431365
transform 1 0 24416 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_240
timestamp 1698431365
transform 1 0 28224 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_274
timestamp 1698431365
transform 1 0 32032 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_308
timestamp 1698431365
transform 1 0 35840 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_342
timestamp 1698431365
transform 1 0 39648 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_376
timestamp 1698431365
transform 1 0 43456 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_410
timestamp 1698431365
transform 1 0 47264 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_444
timestamp 1698431365
transform 1 0 51072 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_478
timestamp 1698431365
transform 1 0 54880 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_486
timestamp 1698431365
transform 1 0 55776 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_490
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_492
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_497
timestamp 1698431365
transform 1 0 57008 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_505
timestamp 1698431365
transform 1 0 57904 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_509
timestamp 1698431365
transform 1 0 58352 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_512
timestamp 1698431365
transform 1 0 58688 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_546
timestamp 1698431365
transform 1 0 62496 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_580
timestamp 1698431365
transform 1 0 66304 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_4 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 65968 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_5
timestamp 1698431365
transform -1 0 40880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_6
timestamp 1698431365
transform -1 0 48944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_7
timestamp 1698431365
transform -1 0 41552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_8
timestamp 1698431365
transform -1 0 55328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_9
timestamp 1698431365
transform -1 0 44240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_10
timestamp 1698431365
transform -1 0 57008 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  grid_clb_11
timestamp 1698431365
transform -1 0 44912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 43456 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 43568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 35168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 29568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 35728 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform 1 0 29232 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform 1 0 33712 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 32704 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 35280 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform 1 0 30464 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 55328 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform 1 0 6384 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 54208 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 51744 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform 1 0 10416 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 59136 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform 1 0 14224 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform 1 0 6384 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 62048 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 59136 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 58128 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform -1 0 54208 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform 1 0 21504 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 25984 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 55216 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform -1 0 39536 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 51408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 16464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 62048 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 44240 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform 1 0 6384 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform 1 0 22064 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 48160 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 51520 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform -1 0 10304 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform -1 0 59248 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform -1 0 59136 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 59136 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 39648 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform -1 0 63168 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform -1 0 50288 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold50
timestamp 1698431365
transform 1 0 18256 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform -1 0 47488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform -1 0 62048 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform -1 0 46368 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform -1 0 62048 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 50288 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 39312 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform -1 0 62048 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform -1 0 63168 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform -1 0 46592 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform -1 0 51296 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform 1 0 10304 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform -1 0 51408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 62048 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform -1 0 62048 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform -1 0 55440 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold69
timestamp 1698431365
transform 1 0 40992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold70
timestamp 1698431365
transform -1 0 41776 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold71
timestamp 1698431365
transform -1 0 43568 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold72
timestamp 1698431365
transform -1 0 63168 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold73
timestamp 1698431365
transform -1 0 59360 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold74
timestamp 1698431365
transform -1 0 63056 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold75
timestamp 1698431365
transform -1 0 62048 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold76
timestamp 1698431365
transform -1 0 35728 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold77
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold78
timestamp 1698431365
transform 1 0 38640 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold79
timestamp 1698431365
transform -1 0 51408 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold80
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold81
timestamp 1698431365
transform 1 0 15344 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold82
timestamp 1698431365
transform -1 0 59584 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold83
timestamp 1698431365
transform -1 0 62048 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold84
timestamp 1698431365
transform -1 0 39984 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold85
timestamp 1698431365
transform -1 0 51744 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold86
timestamp 1698431365
transform -1 0 31808 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold87
timestamp 1698431365
transform -1 0 46368 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold88
timestamp 1698431365
transform -1 0 62048 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold89
timestamp 1698431365
transform -1 0 59136 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold90
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold91
timestamp 1698431365
transform -1 0 59136 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold92
timestamp 1698431365
transform 1 0 21952 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold93
timestamp 1698431365
transform -1 0 59136 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold94
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold95
timestamp 1698431365
transform 1 0 3584 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold96
timestamp 1698431365
transform -1 0 63168 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold97
timestamp 1698431365
transform -1 0 9968 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold98
timestamp 1698431365
transform 1 0 18144 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold99
timestamp 1698431365
transform -1 0 63168 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold100
timestamp 1698431365
transform -1 0 37296 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold101
timestamp 1698431365
transform -1 0 59248 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold102
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold103
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold104
timestamp 1698431365
transform -1 0 44240 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold105
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold106
timestamp 1698431365
transform 1 0 1680 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold107
timestamp 1698431365
transform -1 0 59248 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold108
timestamp 1698431365
transform 1 0 18144 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold109
timestamp 1698431365
transform 1 0 18144 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold110
timestamp 1698431365
transform -1 0 51856 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold111
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold112
timestamp 1698431365
transform -1 0 36064 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold113
timestamp 1698431365
transform -1 0 11536 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold114
timestamp 1698431365
transform -1 0 63168 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold115
timestamp 1698431365
transform -1 0 63168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold116
timestamp 1698431365
transform -1 0 20384 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold117
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold118
timestamp 1698431365
transform -1 0 59248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold119
timestamp 1698431365
transform 1 0 29344 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold120
timestamp 1698431365
transform -1 0 55664 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold121
timestamp 1698431365
transform -1 0 47824 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold122
timestamp 1698431365
transform -1 0 24304 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold123
timestamp 1698431365
transform -1 0 27888 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold124
timestamp 1698431365
transform -1 0 63168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold125
timestamp 1698431365
transform -1 0 59248 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold126
timestamp 1698431365
transform -1 0 59248 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold127
timestamp 1698431365
transform -1 0 62048 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold128
timestamp 1698431365
transform -1 0 16464 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold129
timestamp 1698431365
transform -1 0 59136 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold130
timestamp 1698431365
transform -1 0 43232 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold131
timestamp 1698431365
transform 1 0 25984 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold132
timestamp 1698431365
transform 1 0 2576 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold133
timestamp 1698431365
transform 1 0 17920 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold134
timestamp 1698431365
transform 1 0 21280 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold135
timestamp 1698431365
transform -1 0 18144 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold136
timestamp 1698431365
transform -1 0 40096 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold137
timestamp 1698431365
transform -1 0 55328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold138
timestamp 1698431365
transform 1 0 17472 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold139
timestamp 1698431365
transform 1 0 9520 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold140
timestamp 1698431365
transform -1 0 59248 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold141
timestamp 1698431365
transform -1 0 63168 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold142
timestamp 1698431365
transform -1 0 65968 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold143
timestamp 1698431365
transform 1 0 29232 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold144
timestamp 1698431365
transform -1 0 38976 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold145
timestamp 1698431365
transform -1 0 62048 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold146
timestamp 1698431365
transform -1 0 43008 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold147
timestamp 1698431365
transform 1 0 6496 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold148
timestamp 1698431365
transform -1 0 43792 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold149
timestamp 1698431365
transform -1 0 59248 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold150
timestamp 1698431365
transform 1 0 3584 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold151
timestamp 1698431365
transform -1 0 47488 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold152
timestamp 1698431365
transform 1 0 3584 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold153
timestamp 1698431365
transform 1 0 12880 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold154
timestamp 1698431365
transform -1 0 63168 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold155
timestamp 1698431365
transform -1 0 55664 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold156
timestamp 1698431365
transform -1 0 35728 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold157
timestamp 1698431365
transform 1 0 6384 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold158
timestamp 1698431365
transform -1 0 54208 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold159
timestamp 1698431365
transform -1 0 43568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold160
timestamp 1698431365
transform -1 0 43568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold161
timestamp 1698431365
transform -1 0 47488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold162
timestamp 1698431365
transform 1 0 11424 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold163
timestamp 1698431365
transform 1 0 36736 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold164
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold165
timestamp 1698431365
transform -1 0 38416 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold166
timestamp 1698431365
transform -1 0 63168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold167
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold168
timestamp 1698431365
transform -1 0 35728 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold169
timestamp 1698431365
transform -1 0 40208 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold170
timestamp 1698431365
transform 1 0 28784 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold171
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold172
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold173
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold174
timestamp 1698431365
transform -1 0 32704 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold175
timestamp 1698431365
transform -1 0 50288 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold176
timestamp 1698431365
transform -1 0 44352 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold177
timestamp 1698431365
transform -1 0 24976 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold178
timestamp 1698431365
transform -1 0 47488 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold179
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold180
timestamp 1698431365
transform -1 0 55216 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold181
timestamp 1698431365
transform -1 0 32032 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold182
timestamp 1698431365
transform -1 0 40544 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold183
timestamp 1698431365
transform 1 0 10416 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold184
timestamp 1698431365
transform 1 0 6496 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold185
timestamp 1698431365
transform -1 0 29904 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold186
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold187
timestamp 1698431365
transform -1 0 59248 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold188
timestamp 1698431365
transform 1 0 15344 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold189
timestamp 1698431365
transform -1 0 29904 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold190
timestamp 1698431365
transform 1 0 6384 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold191
timestamp 1698431365
transform -1 0 58464 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold192
timestamp 1698431365
transform -1 0 59248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold193
timestamp 1698431365
transform -1 0 59248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold194
timestamp 1698431365
transform 1 0 18144 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold195
timestamp 1698431365
transform 1 0 2576 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold196
timestamp 1698431365
transform -1 0 59248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold197
timestamp 1698431365
transform -1 0 59248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold198
timestamp 1698431365
transform -1 0 25984 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold199
timestamp 1698431365
transform 1 0 7504 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold200
timestamp 1698431365
transform 1 0 6496 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold201
timestamp 1698431365
transform -1 0 59248 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold202
timestamp 1698431365
transform 1 0 23184 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold203
timestamp 1698431365
transform 1 0 19264 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold204
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold205
timestamp 1698431365
transform -1 0 36512 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold206
timestamp 1698431365
transform 1 0 18144 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold207
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold208
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold209
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold210
timestamp 1698431365
transform -1 0 50288 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold211
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold212
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold213
timestamp 1698431365
transform -1 0 24976 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold214
timestamp 1698431365
transform -1 0 51296 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold215
timestamp 1698431365
transform 1 0 3584 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold216
timestamp 1698431365
transform -1 0 59248 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold217
timestamp 1698431365
transform -1 0 56112 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold218
timestamp 1698431365
transform -1 0 21952 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold219
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold220
timestamp 1698431365
transform -1 0 28784 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold221
timestamp 1698431365
transform 1 0 26096 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold222
timestamp 1698431365
transform 1 0 3584 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold223
timestamp 1698431365
transform 1 0 10304 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold224
timestamp 1698431365
transform -1 0 62048 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold225
timestamp 1698431365
transform -1 0 51296 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold226
timestamp 1698431365
transform -1 0 28784 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold227
timestamp 1698431365
transform -1 0 38528 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold228
timestamp 1698431365
transform -1 0 59248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold229
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold230
timestamp 1698431365
transform -1 0 63168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold231
timestamp 1698431365
transform -1 0 29120 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold232
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold233
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold234
timestamp 1698431365
transform -1 0 55328 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold235
timestamp 1698431365
transform 1 0 2576 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold236
timestamp 1698431365
transform -1 0 42448 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold237
timestamp 1698431365
transform 1 0 10304 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold238
timestamp 1698431365
transform -1 0 59248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold239
timestamp 1698431365
transform -1 0 59248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold240
timestamp 1698431365
transform -1 0 47488 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold241
timestamp 1698431365
transform -1 0 35616 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold242
timestamp 1698431365
transform 1 0 33824 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold243
timestamp 1698431365
transform 1 0 6272 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold244
timestamp 1698431365
transform -1 0 10304 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold245
timestamp 1698431365
transform -1 0 23520 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold246
timestamp 1698431365
transform 1 0 6384 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold247
timestamp 1698431365
transform 1 0 5712 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold248
timestamp 1698431365
transform -1 0 46368 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold249
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold250
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold251
timestamp 1698431365
transform -1 0 23968 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold252
timestamp 1698431365
transform -1 0 29232 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold253
timestamp 1698431365
transform -1 0 44352 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold254
timestamp 1698431365
transform -1 0 33600 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold255
timestamp 1698431365
transform -1 0 24192 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold256
timestamp 1698431365
transform -1 0 19712 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold257
timestamp 1698431365
transform -1 0 19824 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold258
timestamp 1698431365
transform -1 0 47488 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold259
timestamp 1698431365
transform -1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold260
timestamp 1698431365
transform -1 0 59248 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold261
timestamp 1698431365
transform 1 0 2464 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold262
timestamp 1698431365
transform -1 0 34272 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold263
timestamp 1698431365
transform -1 0 58128 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output3 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 64848 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_78 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 66640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 66640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 66640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 66640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 66640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 66640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 66640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 66640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 66640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 66640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 66640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 66640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 66640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 66640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 66640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 66640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 66640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 66640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 66640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 66640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 66640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 66640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 66640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 66640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 66640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 66640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 66640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 66640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 66640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 66640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 66640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 66640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 66640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 66640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 66640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 66640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 66640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 66640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 66640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 66640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 66640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 66640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 66640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 66640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 66640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 66640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 66640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 66640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 66640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 66640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 66640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 66640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 66640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 66640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 66640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 66640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 66640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 66640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 66640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 66640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 66640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 66640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 66640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 66640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 66640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 66640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 66640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 66640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 66640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 66640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 66640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 66640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 66640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 66640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 66640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 66640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 66640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 66640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_156 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_157
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_158
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_159
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_160
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_161
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_162
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_163
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_164
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_165
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_166
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_167
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_168
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_169
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_170
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_171
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_172
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_173
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_174
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_175
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_176
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_177
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_178
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_179
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_180
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_181
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_182
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_183
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_184
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_185
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_186
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_187
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_188
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_189
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_190
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_191
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_192
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_193
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_194
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_195
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_196
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_197
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_198
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_199
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_200
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_201
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_202
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_203
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_204
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_205
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_206
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_207
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_208
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_209
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_210
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_211
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_212
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_213
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_214
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_215
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_216
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_217
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_218
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_219
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_220
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_221
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_222
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_223
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_224
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_225
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_226
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_227
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_228
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_229
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_230
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_231
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_232
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_233
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_234
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_235
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_236
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_237
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_238
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_239
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_240
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_241
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_242
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_243
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_244
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_245
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_246
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_247
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_248
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_249
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_250
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_251
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_252
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_253
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_254
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_255
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_256
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_257
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_258
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_259
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_260
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_261
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_262
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_263
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_264
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_265
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_266
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_267
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_268
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_269
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_270
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_271
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_272
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_273
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_274
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_275
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_276
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_277
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_278
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_279
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_280
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_281
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_282
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_283
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_284
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_285
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_286
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_287
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_288
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_289
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_290
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_291
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_292
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_293
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_294
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_295
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_296
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_297
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_298
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_299
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_300
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_301
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_302
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_303
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_304
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_305
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_306
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_307
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_308
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_309
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_310
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_311
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_312
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_313
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_314
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_315
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_316
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_317
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_318
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_319
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_320
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_321
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_322
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_323
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_324
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_325
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_326
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_327
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_328
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_329
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_330
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_331
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_332
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_333
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_334
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_335
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_336
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_337
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_338
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_339
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_340
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_341
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_342
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_343
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_344
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_345
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_346
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_347
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_348
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_349
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_350
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_351
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_352
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_353
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_354
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_355
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_356
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_357
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_358
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_359
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_360
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_361
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_362
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_363
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_364
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_365
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_366
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_367
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_368
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_369
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_370
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_371
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_372
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_373
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_374
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_375
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_376
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_377
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_378
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_379
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_380
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_381
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_382
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_383
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_384
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_385
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_386
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_387
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_388
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_389
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_390
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_391
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_392
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_393
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_394
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_395
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_396
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_397
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_398
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_399
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_400
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_401
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_402
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_403
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_404
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_405
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_406
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_407
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_408
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_409
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_410
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_411
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_412
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_413
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_414
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_415
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_416
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_417
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_418
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_419
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_420
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_421
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_422
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_423
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_424
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_425
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_426
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_427
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_428
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_429
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_430
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_431
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_432
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_433
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_434
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_435
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_436
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_437
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_438
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_439
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_440
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_441
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_442
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_443
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_444
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_445
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_446
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_447
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_448
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_449
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_450
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_451
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_452
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_453
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_454
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_455
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_456
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_457
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_458
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_459
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_460
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_461
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_462
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_463
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_464
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_465
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_466
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_467
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_468
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_469
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_470
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_471
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_472
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_473
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_474
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_475
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_476
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_477
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_478
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_479
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_480
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_481
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_482
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_483
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_484
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_485
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_486
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_487
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_488
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_489
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_490
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_491
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_492
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_493
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_494
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_495
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_496
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_497
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_498
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_499
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_500
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_501
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_502
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_503
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_504
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_505
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_506
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_507
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_508
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_509
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_510
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_511
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_512
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_513
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_514
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_515
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_516
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_517
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_518
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_519
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_520
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_521
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_522
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_523
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_524
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_525
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_526
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_527
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_528
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_529
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_530
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_531
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_532
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_533
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_534
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_535
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_536
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_537
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_538
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_539
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_540
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_541
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_542
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_543
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_544
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_545
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_546
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_547
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_548
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_549
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_550
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_551
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_552
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_553
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_554
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_555
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_556
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_557
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_558
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_559
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_560
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_561
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_562
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_563
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_564
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_565
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_566
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_567
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_568
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_569
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_570
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_571
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_572
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_573
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_574
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_575
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_576
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_577
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_578
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_579
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_580
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_581
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_582
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_583
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_584
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_585
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_586
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_587
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_588
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_589
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_590
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_591
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_592
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_593
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_594
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_595
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_596
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_597
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_598
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_599
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_600
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_601
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_602
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_603
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_604
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_605
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_606
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_607
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_608
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_609
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_610
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_611
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_612
timestamp 1698431365
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_613
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_614
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_615
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_616
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_617
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_618
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_619
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_620
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_621
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_622
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_623
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_624
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_625
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_626
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_627
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_628
timestamp 1698431365
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_629
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_630
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_631
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_632
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_633
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_634
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_635
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_636
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_637
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_638
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_639
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_640
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_641
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_642
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_643
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_644
timestamp 1698431365
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_645
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_646
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_647
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_648
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_649
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_650
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_651
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_652
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_653
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_654
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_655
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_656
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_657
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_658
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_659
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_660
timestamp 1698431365
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_661
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_662
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_663
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_664
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_665
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_666
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_667
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_668
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_669
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_670
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_671
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_672
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_673
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_674
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_675
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_676
timestamp 1698431365
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_677
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_678
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_679
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_680
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_681
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_682
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_683
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_684
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_685
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_686
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_687
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_688
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_689
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_690
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_691
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_692
timestamp 1698431365
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_693
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_694
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_695
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_696
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_697
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_698
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_699
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_700
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_701
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_702
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_703
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_704
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_705
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_706
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_707
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_708
timestamp 1698431365
transform 1 0 64064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_709
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_710
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_711
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_712
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_713
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_714
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_715
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_716
timestamp 1698431365
transform 1 0 60144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_717
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_718
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_719
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_720
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_721
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_722
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_723
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_724
timestamp 1698431365
transform 1 0 64064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_725
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_726
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_727
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_728
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_729
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_730
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_731
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_732
timestamp 1698431365
transform 1 0 60144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_733
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_734
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_735
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_736
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_737
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_738
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_739
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_740
timestamp 1698431365
transform 1 0 64064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_741
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_742
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_743
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_744
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_745
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_746
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_747
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_748
timestamp 1698431365
transform 1 0 60144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_749
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_750
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_751
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_752
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_753
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_754
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_755
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_756
timestamp 1698431365
transform 1 0 64064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_757
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_758
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_759
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_760
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_761
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_762
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_763
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_764
timestamp 1698431365
transform 1 0 60144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_765
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_766
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_767
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_768
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_769
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_770
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_771
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_772
timestamp 1698431365
transform 1 0 64064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_773
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_774
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_775
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_776
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_777
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_778
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_779
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_780
timestamp 1698431365
transform 1 0 60144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_781
timestamp 1698431365
transform 1 0 5152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_782
timestamp 1698431365
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_783
timestamp 1698431365
transform 1 0 12768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_784
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_785
timestamp 1698431365
transform 1 0 20384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_786
timestamp 1698431365
transform 1 0 24192 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_787
timestamp 1698431365
transform 1 0 28000 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_788
timestamp 1698431365
transform 1 0 31808 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_789
timestamp 1698431365
transform 1 0 35616 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_790
timestamp 1698431365
transform 1 0 39424 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_791
timestamp 1698431365
transform 1 0 43232 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_792
timestamp 1698431365
transform 1 0 47040 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_793
timestamp 1698431365
transform 1 0 50848 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_794
timestamp 1698431365
transform 1 0 54656 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_795
timestamp 1698431365
transform 1 0 58464 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_796
timestamp 1698431365
transform 1 0 62272 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_797
timestamp 1698431365
transform 1 0 66080 0 -1 64288
box -86 -86 310 870
<< labels >>
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 bottom_width_0_height_0_subtile_0__pin_I_10_
port 0 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 bottom_width_0_height_0_subtile_0__pin_I_2_
port 1 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 bottom_width_0_height_0_subtile_0__pin_I_6_
port 2 nsew signal input
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 bottom_width_0_height_0_subtile_0__pin_O_2_
port 3 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 bottom_width_0_height_0_subtile_0__pin_O_6_
port 4 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 ccff_head
port 5 nsew signal input
flabel metal3 s 67200 30912 68000 31024 0 FreeSans 448 0 0 0 ccff_tail
port 6 nsew signal tristate
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 clk
port 7 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 left_width_0_height_0_subtile_0__pin_I_11_
port 8 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 left_width_0_height_0_subtile_0__pin_I_3_
port 9 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 left_width_0_height_0_subtile_0__pin_I_7_
port 10 nsew signal input
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 left_width_0_height_0_subtile_0__pin_O_3_
port 11 nsew signal tristate
flabel metal3 s 67200 62496 68000 62608 0 FreeSans 448 0 0 0 left_width_0_height_0_subtile_0__pin_O_7_
port 12 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 pReset
port 13 nsew signal input
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 prog_clk
port 14 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 reset
port 15 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 right_width_0_height_0_subtile_0__pin_I_1_
port 16 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 right_width_0_height_0_subtile_0__pin_I_5_
port 17 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 right_width_0_height_0_subtile_0__pin_I_9_
port 18 nsew signal input
flabel metal2 s 54432 0 54544 800 0 FreeSans 448 90 0 0 right_width_0_height_0_subtile_0__pin_O_1_
port 19 nsew signal tristate
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 right_width_0_height_0_subtile_0__pin_O_5_
port 20 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 set
port 21 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 top_width_0_height_0_subtile_0__pin_I_0_
port 22 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 top_width_0_height_0_subtile_0__pin_I_4_
port 23 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 top_width_0_height_0_subtile_0__pin_I_8_
port 24 nsew signal input
flabel metal2 s 56448 67200 56560 68000 0 FreeSans 448 90 0 0 top_width_0_height_0_subtile_0__pin_O_0_
port 25 nsew signal tristate
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 top_width_0_height_0_subtile_0__pin_O_4_
port 26 nsew signal tristate
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 top_width_0_height_0_subtile_0__pin_clk_0_
port 27 nsew signal input
flabel metal4 s 4448 3076 4768 64348 0 FreeSans 1280 90 0 0 vdd
port 28 nsew power bidirectional
flabel metal4 s 35168 3076 35488 64348 0 FreeSans 1280 90 0 0 vdd
port 28 nsew power bidirectional
flabel metal4 s 65888 3076 66208 64348 0 FreeSans 1280 90 0 0 vdd
port 28 nsew power bidirectional
flabel metal4 s 19808 3076 20128 64348 0 FreeSans 1280 90 0 0 vss
port 29 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 64348 0 FreeSans 1280 90 0 0 vss
port 29 nsew ground bidirectional
rlabel metal1 33992 63504 33992 63504 0 vdd
rlabel metal1 33992 64288 33992 64288 0 vss
rlabel metal2 53144 28000 53144 28000 0 _000_
rlabel metal2 47768 28392 47768 28392 0 _001_
rlabel metal2 48216 26124 48216 26124 0 _002_
rlabel metal3 48552 27720 48552 27720 0 _003_
rlabel metal2 51688 29848 51688 29848 0 _004_
rlabel metal2 51576 29120 51576 29120 0 _005_
rlabel metal2 53144 29848 53144 29848 0 _006_
rlabel metal2 54600 29512 54600 29512 0 _007_
rlabel metal2 55720 29736 55720 29736 0 _008_
rlabel metal2 59528 29960 59528 29960 0 _009_
rlabel metal2 51688 22120 51688 22120 0 _010_
rlabel metal2 51184 22120 51184 22120 0 _011_
rlabel metal2 51800 22792 51800 22792 0 _012_
rlabel metal2 55160 23240 55160 23240 0 _013_
rlabel metal2 55720 22176 55720 22176 0 _014_
rlabel metal2 54376 23744 54376 23744 0 _015_
rlabel metal3 57792 25256 57792 25256 0 _016_
rlabel metal2 55160 24976 55160 24976 0 _017_
rlabel metal2 55496 26656 55496 26656 0 _018_
rlabel metal2 59304 27384 59304 27384 0 _019_
rlabel metal2 47880 25088 47880 25088 0 _020_
rlabel metal3 49000 24920 49000 24920 0 _021_
rlabel metal2 46312 21224 46312 21224 0 _022_
rlabel metal2 42392 23184 42392 23184 0 _023_
rlabel metal2 43624 20552 43624 20552 0 _024_
rlabel metal2 43904 20888 43904 20888 0 _025_
rlabel metal3 45920 20104 45920 20104 0 _026_
rlabel metal2 47208 20272 47208 20272 0 _027_
rlabel metal2 47768 20328 47768 20328 0 _028_
rlabel metal2 48104 21000 48104 21000 0 _029_
rlabel metal2 40936 29736 40936 29736 0 _030_
rlabel metal2 41552 28504 41552 28504 0 _031_
rlabel metal2 43400 26236 43400 26236 0 _032_
rlabel metal2 41664 28056 41664 28056 0 _033_
rlabel metal2 39928 28168 39928 28168 0 _034_
rlabel metal2 39816 27496 39816 27496 0 _035_
rlabel metal2 39704 25648 39704 25648 0 _036_
rlabel metal2 41608 25312 41608 25312 0 _037_
rlabel metal2 43848 26208 43848 26208 0 _038_
rlabel metal2 49112 25648 49112 25648 0 _039_
rlabel metal2 34328 33824 34328 33824 0 _040_
rlabel metal2 35896 32368 35896 32368 0 _041_
rlabel metal3 35392 31864 35392 31864 0 _042_
rlabel metal2 29512 32984 29512 32984 0 _043_
rlabel metal2 33768 29568 33768 29568 0 _044_
rlabel metal2 30520 29120 30520 29120 0 _045_
rlabel metal2 33096 29736 33096 29736 0 _046_
rlabel metal3 38024 31192 38024 31192 0 _047_
rlabel metal2 36064 28728 36064 28728 0 _048_
rlabel metal2 37352 28000 37352 28000 0 _049_
rlabel metal3 41440 33432 41440 33432 0 _050_
rlabel metal2 42952 32368 42952 32368 0 _051_
rlabel metal2 44408 33040 44408 33040 0 _052_
rlabel metal2 46312 33992 46312 33992 0 _053_
rlabel metal2 39928 32928 39928 32928 0 _054_
rlabel metal2 41160 31584 41160 31584 0 _055_
rlabel metal2 43736 31360 43736 31360 0 _056_
rlabel metal2 45304 30576 45304 30576 0 _057_
rlabel metal3 49728 31528 49728 31528 0 _058_
rlabel metal2 47768 30632 47768 30632 0 _059_
rlabel metal2 55888 39368 55888 39368 0 _060_
rlabel metal2 51464 37184 51464 37184 0 _061_
rlabel metal2 53144 37408 53144 37408 0 _062_
rlabel metal2 55160 36008 55160 36008 0 _063_
rlabel metal2 55720 35112 55720 35112 0 _064_
rlabel metal2 50008 35112 50008 35112 0 _065_
rlabel metal2 51576 34552 51576 34552 0 _066_
rlabel metal2 51744 33096 51744 33096 0 _067_
rlabel metal2 54488 34160 54488 34160 0 _068_
rlabel metal2 55384 34496 55384 34496 0 _069_
rlabel metal2 49168 44072 49168 44072 0 _070_
rlabel metal2 51576 42784 51576 42784 0 _071_
rlabel metal2 51688 41888 51688 41888 0 _072_
rlabel metal3 56896 44184 56896 44184 0 _073_
rlabel metal3 60816 41832 60816 41832 0 _074_
rlabel metal2 59304 41720 59304 41720 0 _075_
rlabel metal2 55720 42168 55720 42168 0 _076_
rlabel metal2 51464 39928 51464 39928 0 _077_
rlabel metal2 52416 39032 52416 39032 0 _078_
rlabel metal2 55160 40488 55160 40488 0 _079_
rlabel metal2 39928 45248 39928 45248 0 _080_
rlabel metal2 43736 43904 43736 43904 0 _081_
rlabel metal2 45192 44800 45192 44800 0 _082_
rlabel metal3 37464 41272 37464 41272 0 _083_
rlabel metal3 41720 41272 41720 41272 0 _084_
rlabel metal2 39928 42952 39928 42952 0 _085_
rlabel metal2 43848 40936 43848 40936 0 _086_
rlabel metal3 44744 41272 44744 41272 0 _087_
rlabel metal2 46536 41888 46536 41888 0 _088_
rlabel metal2 47208 41664 47208 41664 0 _089_
rlabel metal2 49504 48440 49504 48440 0 _090_
rlabel metal2 51576 48048 51576 48048 0 _091_
rlabel metal2 53368 49952 53368 49952 0 _092_
rlabel metal2 55608 47656 55608 47656 0 _093_
rlabel metal3 54348 46760 54348 46760 0 _094_
rlabel metal2 55720 45752 55720 45752 0 _095_
rlabel metal2 58968 44800 58968 44800 0 _096_
rlabel metal2 50232 44800 50232 44800 0 _097_
rlabel metal2 51576 44520 51576 44520 0 _098_
rlabel metal3 53368 43624 53368 43624 0 _099_
rlabel metal2 38920 47488 38920 47488 0 _100_
rlabel metal2 42168 47992 42168 47992 0 _101_
rlabel metal2 39984 46760 39984 46760 0 _102_
rlabel metal3 42000 48776 42000 48776 0 _103_
rlabel metal2 43736 46956 43736 46956 0 _104_
rlabel metal2 45416 49952 45416 49952 0 _105_
rlabel metal3 46368 45304 46368 45304 0 _106_
rlabel metal2 44856 49056 44856 49056 0 _107_
rlabel metal2 46872 46032 46872 46032 0 _108_
rlabel metal2 47880 49280 47880 49280 0 _109_
rlabel metal2 29512 45640 29512 45640 0 _110_
rlabel metal3 30800 45752 30800 45752 0 _111_
rlabel metal2 27944 46480 27944 46480 0 _112_
rlabel metal2 29288 48664 29288 48664 0 _113_
rlabel metal2 30968 47488 30968 47488 0 _114_
rlabel metal2 32200 45640 32200 45640 0 _115_
rlabel metal2 34216 46200 34216 46200 0 _116_
rlabel metal2 35896 47824 35896 47824 0 _117_
rlabel metal3 33152 45304 33152 45304 0 _118_
rlabel metal2 35784 47208 35784 47208 0 _119_
rlabel metal2 21560 42784 21560 42784 0 _120_
rlabel metal3 23240 41272 23240 41272 0 _121_
rlabel metal2 27496 43008 27496 43008 0 _122_
rlabel metal2 25816 43344 25816 43344 0 _123_
rlabel metal2 17752 43848 17752 43848 0 _124_
rlabel metal2 23688 45752 23688 45752 0 _125_
rlabel metal2 17752 45416 17752 45416 0 _126_
rlabel metal2 23912 47488 23912 47488 0 _127_
rlabel metal2 24248 47096 24248 47096 0 _128_
rlabel metal3 27832 48776 27832 48776 0 _129_
rlabel metal3 30408 38920 30408 38920 0 _130_
rlabel metal2 31864 41216 31864 41216 0 _131_
rlabel metal3 36176 40936 36176 40936 0 _132_
rlabel metal2 36456 40824 36456 40824 0 _133_
rlabel metal2 25928 41664 25928 41664 0 _134_
rlabel metal2 28504 40040 28504 40040 0 _135_
rlabel metal3 30912 43624 30912 43624 0 _136_
rlabel metal2 32200 42952 32200 42952 0 _137_
rlabel metal2 34776 41888 34776 41888 0 _138_
rlabel metal2 36008 44128 36008 44128 0 _139_
rlabel metal2 40152 36736 40152 36736 0 _140_
rlabel metal2 42168 37856 42168 37856 0 _141_
rlabel metal2 43736 36120 43736 36120 0 _142_
rlabel metal2 47768 37296 47768 37296 0 _143_
rlabel metal2 47656 37576 47656 37576 0 _144_
rlabel metal2 49000 37296 49000 37296 0 _145_
rlabel metal3 48216 38696 48216 38696 0 _146_
rlabel metal2 42728 40712 42728 40712 0 _147_
rlabel metal2 41720 40264 41720 40264 0 _148_
rlabel metal2 43960 40040 43960 40040 0 _149_
rlabel metal3 31612 34328 31612 34328 0 _150_
rlabel metal2 33544 33600 33544 33600 0 _151_
rlabel metal2 29176 36904 29176 36904 0 _152_
rlabel metal2 32592 36232 32592 36232 0 _153_
rlabel metal2 31864 36624 31864 36624 0 _154_
rlabel metal2 34328 37632 34328 37632 0 _155_
rlabel metal2 36008 36288 36008 36288 0 _156_
rlabel metal2 37744 35896 37744 35896 0 _157_
rlabel metal2 37128 36008 37128 36008 0 _158_
rlabel metal2 38528 37464 38528 37464 0 _159_
rlabel metal2 12712 35952 12712 35952 0 _160_
rlabel metal2 16520 35000 16520 35000 0 _161_
rlabel metal2 16520 36008 16520 36008 0 _162_
rlabel metal2 11928 34384 11928 34384 0 _163_
rlabel metal2 12488 36288 12488 36288 0 _164_
rlabel metal2 15848 36232 15848 36232 0 _165_
rlabel metal2 10024 39536 10024 39536 0 _166_
rlabel metal2 16408 39032 16408 39032 0 _167_
rlabel metal2 17416 36512 17416 36512 0 _168_
rlabel metal2 16296 39928 16296 39928 0 _169_
rlabel metal2 20328 37688 20328 37688 0 _170_
rlabel metal2 20216 39424 20216 39424 0 _171_
rlabel metal2 23128 40936 23128 40936 0 _172_
rlabel metal2 22232 40096 22232 40096 0 _173_
rlabel metal2 26712 40096 26712 40096 0 _174_
rlabel metal2 21896 39256 21896 39256 0 _175_
rlabel metal2 26824 40712 26824 40712 0 _176_
rlabel metal2 20216 37688 20216 37688 0 _177_
rlabel metal2 19656 36904 19656 36904 0 _178_
rlabel metal2 24248 37408 24248 37408 0 _179_
rlabel metal3 20944 33432 20944 33432 0 _180_
rlabel metal3 26768 33320 26768 33320 0 _181_
rlabel metal2 27048 35616 27048 35616 0 _182_
rlabel metal2 24304 32648 24304 32648 0 _183_
rlabel metal2 21448 30632 21448 30632 0 _184_
rlabel metal2 22568 30744 22568 30744 0 _185_
rlabel metal2 23016 32200 23016 32200 0 _186_
rlabel metal2 23968 29624 23968 29624 0 _187_
rlabel metal2 24360 30240 24360 30240 0 _188_
rlabel metal2 25144 29176 25144 29176 0 _189_
rlabel metal3 9464 27944 9464 27944 0 _190_
rlabel metal2 12712 29176 12712 29176 0 _191_
rlabel metal2 13720 27552 13720 27552 0 _192_
rlabel metal2 15064 27440 15064 27440 0 _193_
rlabel metal2 8456 27216 8456 27216 0 _194_
rlabel metal2 7560 24752 7560 24752 0 _195_
rlabel metal2 12040 25872 12040 25872 0 _196_
rlabel metal2 7448 27440 7448 27440 0 _197_
rlabel metal3 6048 28728 6048 28728 0 _198_
rlabel metal2 7896 29120 7896 29120 0 _199_
rlabel metal3 9632 30296 9632 30296 0 _200_
rlabel metal2 12488 30744 12488 30744 0 _201_
rlabel metal3 13048 30184 13048 30184 0 _202_
rlabel metal2 15400 31416 15400 31416 0 _203_
rlabel metal2 16464 33992 16464 33992 0 _204_
rlabel metal2 17864 31024 17864 31024 0 _205_
rlabel metal2 16520 31976 16520 31976 0 _206_
rlabel metal2 11480 35728 11480 35728 0 _207_
rlabel metal2 13496 34048 13496 34048 0 _208_
rlabel metal2 8904 30576 8904 30576 0 _209_
rlabel metal2 28224 27160 28224 27160 0 _210_
rlabel metal2 28280 28336 28280 28336 0 _211_
rlabel metal2 29400 25872 29400 25872 0 _212_
rlabel metal2 31864 27328 31864 27328 0 _213_
rlabel metal2 33656 28168 33656 28168 0 _214_
rlabel metal3 28560 24024 28560 24024 0 _215_
rlabel metal2 28168 24528 28168 24528 0 _216_
rlabel metal2 32144 27720 32144 27720 0 _217_
rlabel metal3 35336 26936 35336 26936 0 _218_
rlabel metal2 34832 26488 34832 26488 0 _219_
rlabel metal2 37520 23352 37520 23352 0 _220_
rlabel metal2 39256 23464 39256 23464 0 _221_
rlabel metal2 37688 22624 37688 22624 0 _222_
rlabel metal2 35560 22960 35560 22960 0 _223_
rlabel metal3 36512 20888 36512 20888 0 _224_
rlabel metal2 36568 21840 36568 21840 0 _225_
rlabel metal2 28280 22904 28280 22904 0 _226_
rlabel metal2 30744 22736 30744 22736 0 _227_
rlabel metal2 32088 23296 32088 23296 0 _228_
rlabel metal2 33768 23296 33768 23296 0 _229_
rlabel metal2 21896 25088 21896 25088 0 _230_
rlabel metal2 24136 24136 24136 24136 0 _231_
rlabel metal2 25928 27272 25928 27272 0 _232_
rlabel metal2 20776 28112 20776 28112 0 _233_
rlabel metal2 20328 27832 20328 27832 0 _234_
rlabel metal3 16016 28056 16016 28056 0 _235_
rlabel metal2 18424 24920 18424 24920 0 _236_
rlabel metal2 18088 26040 18088 26040 0 _237_
rlabel metal3 24640 19096 24640 19096 0 _238_
rlabel metal2 24808 21056 24808 21056 0 _239_
rlabel metal2 10248 23520 10248 23520 0 _240_
rlabel metal2 6216 24472 6216 24472 0 _241_
rlabel metal2 8344 25144 8344 25144 0 _242_
rlabel metal2 8344 23968 8344 23968 0 _243_
rlabel metal2 12264 24416 12264 24416 0 _244_
rlabel metal2 5880 25088 5880 25088 0 _245_
rlabel metal2 8344 20888 8344 20888 0 _246_
rlabel metal2 8736 22120 8736 22120 0 _247_
rlabel metal2 10304 21784 10304 21784 0 _248_
rlabel metal2 13832 21336 13832 21336 0 _249_
rlabel metal2 14056 23800 14056 23800 0 _250_
rlabel metal2 16520 21112 16520 21112 0 _251_
rlabel metal2 15624 21056 15624 21056 0 _252_
rlabel metal2 18200 20328 18200 20328 0 _253_
rlabel metal2 18536 20160 18536 20160 0 _254_
rlabel metal2 20104 21336 20104 21336 0 _255_
rlabel metal2 22008 19544 22008 19544 0 _256_
rlabel metal2 20664 21336 20664 21336 0 _257_
rlabel metal3 17752 24024 17752 24024 0 _258_
rlabel metal2 21784 25984 21784 25984 0 _259_
rlabel metal2 20664 25088 20664 25088 0 _260_
rlabel metal2 23912 27328 23912 27328 0 _261_
rlabel metal3 21392 34104 21392 34104 0 _262_
rlabel metal2 20216 34496 20216 34496 0 _263_
rlabel metal2 26040 36456 26040 36456 0 _264_
rlabel metal2 26656 28056 26656 28056 0 _265_
rlabel metal2 48216 29120 48216 29120 0 _266_
rlabel metal2 55384 25480 55384 25480 0 _267_
rlabel metal2 49952 24808 49952 24808 0 _268_
rlabel metal2 46984 26096 46984 26096 0 _269_
rlabel metal2 33432 29008 33432 29008 0 _270_
rlabel metal2 47992 33824 47992 33824 0 _271_
rlabel metal2 44296 47880 44296 47880 0 _272_
rlabel metal2 50344 36176 50344 36176 0 _273_
rlabel metal2 50792 44072 50792 44072 0 _274_
rlabel metal2 45416 44240 45416 44240 0 _275_
rlabel metal3 48720 49672 48720 49672 0 _276_
rlabel metal2 46424 49336 46424 49336 0 _277_
rlabel metal2 36176 48216 36176 48216 0 _278_
rlabel metal2 21672 46088 21672 46088 0 _279_
rlabel metal2 32312 39704 32312 39704 0 _280_
rlabel metal2 48720 38696 48720 38696 0 _281_
rlabel metal2 38080 38136 38080 38136 0 _282_
rlabel metal2 26040 29624 26040 29624 0 _283_
rlabel metal2 14056 36680 14056 36680 0 _284_
rlabel metal2 20664 37912 20664 37912 0 _285_
rlabel metal3 22008 30184 22008 30184 0 _286_
rlabel metal3 7448 28616 7448 28616 0 _287_
rlabel metal2 9128 31080 9128 31080 0 _288_
rlabel metal2 28616 27944 28616 27944 0 _289_
rlabel metal3 39256 23128 39256 23128 0 _290_
rlabel metal3 22008 27048 22008 27048 0 _291_
rlabel metal2 5992 25928 5992 25928 0 _292_
rlabel metal2 15288 23128 15288 23128 0 _293_
rlabel metal2 1736 25144 1736 25144 0 ccff_head
rlabel metal3 66682 30968 66682 30968 0 ccff_tail
rlabel metal2 28504 34048 28504 34048 0 clknet_0_prog_clk
rlabel metal2 26096 30856 26096 30856 0 clknet_1_0__leaf_prog_clk
rlabel metal2 53032 22344 53032 22344 0 clknet_1_1__leaf_prog_clk
rlabel via2 1848 26264 1848 26264 0 clknet_leaf_0_prog_clk
rlabel metal3 46872 39704 46872 39704 0 clknet_leaf_10_prog_clk
rlabel metal2 48832 39368 48832 39368 0 clknet_leaf_11_prog_clk
rlabel metal2 31864 33488 31864 33488 0 clknet_leaf_12_prog_clk
rlabel metal2 53088 26488 53088 26488 0 clknet_leaf_13_prog_clk
rlabel metal2 52752 26488 52752 26488 0 clknet_leaf_14_prog_clk
rlabel metal2 52472 23912 52472 23912 0 clknet_leaf_15_prog_clk
rlabel metal3 48552 20104 48552 20104 0 clknet_leaf_16_prog_clk
rlabel metal3 30352 25480 30352 25480 0 clknet_leaf_17_prog_clk
rlabel metal2 31192 28616 31192 28616 0 clknet_leaf_18_prog_clk
rlabel metal2 29288 30968 29288 30968 0 clknet_leaf_19_prog_clk
rlabel metal2 24024 31472 24024 31472 0 clknet_leaf_1_prog_clk
rlabel metal2 27720 26936 27720 26936 0 clknet_leaf_20_prog_clk
rlabel metal2 15848 21560 15848 21560 0 clknet_leaf_21_prog_clk
rlabel metal3 5656 21616 5656 21616 0 clknet_leaf_22_prog_clk
rlabel metal2 28616 31472 28616 31472 0 clknet_leaf_2_prog_clk
rlabel metal2 9352 36400 9352 36400 0 clknet_leaf_3_prog_clk
rlabel metal2 26488 47432 26488 47432 0 clknet_leaf_4_prog_clk
rlabel metal3 22680 38024 22680 38024 0 clknet_leaf_5_prog_clk
rlabel metal3 40208 41944 40208 41944 0 clknet_leaf_6_prog_clk
rlabel metal2 42000 48216 42000 48216 0 clknet_leaf_7_prog_clk
rlabel metal2 45976 44072 45976 44072 0 clknet_leaf_8_prog_clk
rlabel metal2 53312 48216 53312 48216 0 clknet_leaf_9_prog_clk
rlabel metal2 24584 18816 24584 18816 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
rlabel metal3 10024 21784 10024 21784 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
rlabel metal3 22400 16744 22400 16744 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
rlabel metal2 3080 22120 3080 22120 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in
rlabel metal2 16184 18480 16184 18480 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in
rlabel metal2 16744 18032 16744 18032 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in
rlabel metal2 18424 17864 18424 17864 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in
rlabel metal2 19768 16184 19768 16184 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in
rlabel metal2 21336 18760 21336 18760 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in
rlabel metal2 22680 15400 22680 15400 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in
rlabel metal2 3192 21560 3192 21560 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in
rlabel metal2 9744 20216 9744 20216 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in
rlabel metal2 12992 24472 12992 24472 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in
rlabel metal2 4088 19152 4088 19152 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in
rlabel metal2 9408 17528 9408 17528 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in
rlabel metal3 10024 22120 10024 22120 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in
rlabel metal2 9632 18088 9632 18088 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in
rlabel metal3 11480 21112 11480 21112 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in
rlabel metal2 10920 21784 10920 21784 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in
rlabel metal2 26320 18984 26320 18984 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q
rlabel metal2 19152 14392 19152 14392 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q
rlabel metal2 17416 17528 17416 17528 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q
rlabel metal2 18872 17528 18872 17528 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q
rlabel metal2 15624 19880 15624 19880 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q
rlabel metal2 20888 26656 20888 26656 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q
rlabel metal2 18760 19712 18760 19712 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q
rlabel metal3 20776 26824 20776 26824 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
rlabel metal3 30576 28392 30576 28392 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
rlabel metal2 24080 17528 24080 17528 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
rlabel metal2 28728 19712 28728 19712 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in
rlabel metal2 33376 15960 33376 15960 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in
rlabel metal3 30072 20328 30072 20328 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in
rlabel metal2 32088 16968 32088 16968 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in
rlabel metal2 33992 17696 33992 17696 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in
rlabel metal2 29624 17472 29624 17472 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in
rlabel metal2 23688 17192 23688 17192 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in
rlabel metal2 29344 16968 29344 16968 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in
rlabel metal3 34048 16968 34048 16968 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in
rlabel metal2 38472 20160 38472 20160 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in
rlabel metal2 34440 20552 34440 20552 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in
rlabel metal2 38920 18816 38920 18816 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in
rlabel metal2 43064 19768 43064 19768 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in
rlabel metal2 36792 18760 36792 18760 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in
rlabel metal2 31528 19040 31528 19040 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in
rlabel metal2 38024 18088 38024 18088 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in
rlabel metal2 29456 18536 29456 18536 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q
rlabel metal3 33208 26824 33208 26824 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q
rlabel metal2 28392 22176 28392 22176 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q
rlabel metal3 29512 24584 29512 24584 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q
rlabel metal3 25312 27608 25312 27608 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q
rlabel metal2 3192 29624 3192 29624 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q
rlabel metal2 20776 28392 20776 28392 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q
rlabel metal2 4200 34160 4200 34160 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
rlabel metal2 6104 29568 6104 29568 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
rlabel metal3 4200 31640 4200 31640 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
rlabel metal2 4536 28784 4536 28784 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in
rlabel metal2 2072 27496 2072 27496 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in
rlabel metal2 3080 27272 3080 27272 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in
rlabel metal2 3080 36008 3080 36008 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in
rlabel metal2 13048 31892 13048 31892 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in
rlabel metal2 3080 33152 3080 33152 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in
rlabel metal3 9576 31080 9576 31080 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in
rlabel metal2 2968 25704 2968 25704 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in
rlabel metal2 13328 23352 13328 23352 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in
rlabel metal2 6664 26432 6664 26432 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in
rlabel metal2 9632 23128 9632 23128 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in
rlabel metal3 5376 20216 5376 20216 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in
rlabel metal3 4928 23800 4928 23800 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in
rlabel metal2 2744 23520 2744 23520 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in
rlabel metal2 8232 23744 8232 23744 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in
rlabel metal2 2856 26992 2856 26992 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in
rlabel metal3 14000 31640 14000 31640 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q
rlabel metal2 25200 26936 25200 26936 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q
rlabel metal2 4200 32816 4200 32816 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q
rlabel metal2 20888 32872 20888 32872 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q
rlabel metal2 4816 30184 4816 30184 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q
rlabel metal2 4256 37352 4256 37352 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q
rlabel metal2 3080 34832 3080 34832 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q
rlabel metal2 18872 30520 18872 30520 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
rlabel metal2 7000 35616 7000 35616 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
rlabel metal2 24808 38696 24808 38696 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
rlabel metal2 7112 37296 7112 37296 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in
rlabel metal2 21112 40824 21112 40824 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in
rlabel metal2 27496 40712 27496 40712 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in
rlabel metal2 21112 39592 21112 39592 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in
rlabel metal2 27720 38304 27720 38304 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in
rlabel metal2 20944 37464 20944 37464 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in
rlabel metal2 19208 36680 19208 36680 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in
rlabel metal2 7000 38528 7000 38528 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in
rlabel metal2 8120 38640 8120 38640 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in
rlabel metal3 11256 40600 11256 40600 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in
rlabel metal2 16968 37968 16968 37968 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in
rlabel metal2 16968 40544 16968 40544 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in
rlabel metal2 17528 46760 17528 46760 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in
rlabel metal2 21000 39200 21000 39200 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in
rlabel metal2 20888 41720 20888 41720 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in
rlabel metal2 23800 42280 23800 42280 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in
rlabel metal2 11928 36624 11928 36624 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q
rlabel metal2 7112 36232 7112 36232 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q
rlabel metal2 21000 34496 21000 34496 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q
rlabel metal2 20888 34440 20888 34440 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q
rlabel metal2 6664 32984 6664 32984 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q
rlabel metal2 24864 34328 24864 34328 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q
rlabel metal2 25704 45976 25704 45976 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q
rlabel metal2 31864 34776 31864 34776 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_0_.Q
rlabel metal2 35000 29428 35000 29428 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_1_.Q
rlabel metal2 28392 37072 28392 37072 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_2_.Q
rlabel metal2 26488 38472 26488 38472 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_3_.Q
rlabel metal2 29960 40432 29960 40432 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_4_.Q
rlabel metal3 39032 38248 39032 38248 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_5_.Q
rlabel metal3 47096 38808 47096 38808 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_6_.Q
rlabel metal2 38528 35896 38528 35896 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_7_.Q
rlabel metal2 42840 44072 42840 44072 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_8_.Q
rlabel metal2 47208 32816 47208 32816 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_9_.Q
rlabel metal3 46312 36680 46312 36680 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_0_.Q
rlabel metal2 55496 39704 55496 39704 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_1_.Q
rlabel metal3 47460 35896 47460 35896 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_2_.Q
rlabel metal2 48384 35896 48384 35896 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_3_.Q
rlabel metal3 49420 37800 49420 37800 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_4_.Q
rlabel metal2 48440 39872 48440 39872 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_5_.Q
rlabel metal3 57064 40544 57064 40544 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_6_.Q
rlabel metal2 38640 50456 38640 50456 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_7_.Q
rlabel metal3 47880 41104 47880 41104 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_8_.Q
rlabel metal2 44632 39256 44632 39256 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_9_.Q
rlabel metal2 18760 41328 18760 41328 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_0_.Q
rlabel metal2 25704 42728 25704 42728 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_1_.Q
rlabel metal2 35840 41384 35840 41384 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_2_.Q
rlabel metal2 33992 50428 33992 50428 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_3_.Q
rlabel metal2 25032 41832 25032 41832 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_4_.Q
rlabel metal2 31416 42224 31416 42224 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_5_.Q
rlabel metal2 27888 51464 27888 51464 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_6_.Q
rlabel metal2 32760 43176 32760 43176 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_7_.Q
rlabel metal3 36400 51464 36400 51464 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_8_.Q
rlabel metal2 32760 42728 32760 42728 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_9_.Q
rlabel metal2 20888 44072 20888 44072 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_0_.Q
rlabel metal2 18424 44072 18424 44072 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_1_.Q
rlabel metal2 26600 49672 26600 49672 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_2_.Q
rlabel metal2 23968 49896 23968 49896 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_3_.Q
rlabel metal2 17192 45080 17192 45080 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_4_.Q
rlabel metal2 24528 45304 24528 45304 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_5_.Q
rlabel metal2 17192 46648 17192 46648 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_6_.Q
rlabel metal2 19544 48048 19544 48048 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_7_.Q
rlabel metal2 24920 47208 24920 47208 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_8_.Q
rlabel metal2 28112 52024 28112 52024 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_9_.Q
rlabel metal2 28728 48272 28728 48272 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_0_.Q
rlabel metal2 22680 47208 22680 47208 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_1_.Q
rlabel metal2 28784 46088 28784 46088 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_2_.Q
rlabel metal2 29960 48832 29960 48832 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_3_.Q
rlabel metal2 31808 53032 31808 53032 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_4_.Q
rlabel metal2 32760 48272 32760 48272 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_5_.Q
rlabel metal3 35560 50792 35560 50792 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_6_.Q
rlabel metal2 39144 50792 39144 50792 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_7_.Q
rlabel metal3 34216 52024 34216 52024 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_8_.Q
rlabel metal3 37688 53032 37688 53032 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_9_.Q
rlabel metal2 39480 49560 39480 49560 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_0_.Q
rlabel metal3 38472 53592 38472 53592 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_1_.Q
rlabel metal2 40488 49448 40488 49448 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_2_.Q
rlabel metal2 43736 53368 43736 53368 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_3_.Q
rlabel metal2 44520 50232 44520 50232 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_4_.Q
rlabel metal2 45976 50736 45976 50736 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_5_.Q
rlabel metal2 44632 49952 44632 49952 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_6_.Q
rlabel metal2 45416 49000 45416 49000 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_7_.Q
rlabel metal2 48440 48272 48440 48272 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_8_.Q
rlabel metal2 48664 49840 48664 49840 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_9_.Q
rlabel metal2 48608 48440 48608 48440 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_0_.Q
rlabel metal2 52248 48216 52248 48216 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_1_.Q
rlabel metal2 53928 50232 53928 50232 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_2_.Q
rlabel metal2 56280 48776 56280 48776 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_3_.Q
rlabel metal2 52472 47376 52472 47376 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_4_.Q
rlabel metal2 56280 46592 56280 46592 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_5_.Q
rlabel metal2 56112 45304 56112 45304 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_6_.Q
rlabel metal2 52360 45528 52360 45528 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_7_.Q
rlabel metal2 61432 45808 61432 45808 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_8_.Q
rlabel metal2 47320 52024 47320 52024 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_9_.Q
rlabel metal2 40544 45304 40544 45304 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_0_.Q
rlabel metal2 44464 46648 44464 46648 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_1_.Q
rlabel metal2 42392 46648 42392 46648 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_2_.Q
rlabel metal2 35896 43400 35896 43400 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_3_.Q
rlabel metal2 40544 45080 40544 45080 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_4_.Q
rlabel metal2 45752 50792 45752 50792 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_5_.Q
rlabel metal2 43960 47068 43960 47068 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_6_.Q
rlabel metal3 47824 46760 47824 46760 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_7_.Q
rlabel metal3 51940 42616 51940 42616 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_8_.Q
rlabel metal2 48328 42560 48328 42560 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_9_.Q
rlabel metal2 49672 45360 49672 45360 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_0_.Q
rlabel metal2 52360 43400 52360 43400 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_1_.Q
rlabel metal2 52248 44744 52248 44744 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_2_.Q
rlabel metal3 59416 42616 59416 42616 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_3_.Q
rlabel metal3 61320 44184 61320 44184 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_4_.Q
rlabel metal2 56168 42784 56168 42784 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_5_.Q
rlabel metal2 56280 41720 56280 41720 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_6_.Q
rlabel metal2 61432 40712 61432 40712 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_7_.Q
rlabel metal2 62552 39200 62552 39200 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_8_.Q
rlabel metal2 56168 40656 56168 40656 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_9_.Q
rlabel metal2 61432 39144 61432 39144 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_0_.Q
rlabel metal2 61432 37576 61432 37576 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_1_.Q
rlabel metal2 53704 36680 53704 36680 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_2_.Q
rlabel metal2 62552 37296 62552 37296 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_3_.Q
rlabel metal3 58912 35112 58912 35112 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_4_.Q
rlabel metal3 62552 34720 62552 34720 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_5_.Q
rlabel metal3 56896 34328 56896 34328 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_6_.Q
rlabel metal2 61432 32872 61432 32872 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_7_.Q
rlabel metal3 62552 33096 62552 33096 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_8_.Q
rlabel metal2 56168 34552 56168 34552 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_9_.Q
rlabel metal3 48776 33544 48776 33544 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_0_.Q
rlabel metal3 52696 34104 52696 34104 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_1_.Q
rlabel metal3 45696 32760 45696 32760 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_2_.Q
rlabel metal2 48440 32928 48440 32928 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_3_.Q
rlabel metal2 40488 32144 40488 32144 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_4_.Q
rlabel metal3 43176 31584 43176 31584 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_5_.Q
rlabel metal3 48608 23800 48608 23800 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_6_.Q
rlabel metal3 48188 29176 48188 29176 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_7_.Q
rlabel metal2 48440 29736 48440 29736 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_8_.Q
rlabel metal2 48328 31528 48328 31528 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_9_.Q
rlabel metal2 21784 35112 21784 35112 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_0_.Q
rlabel metal2 47096 32032 47096 32032 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_1_.Q
rlabel metal3 34384 30296 34384 30296 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_2_.Q
rlabel metal3 29232 24248 29232 24248 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_3_.Q
rlabel metal2 32536 31528 32536 31528 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_4_.Q
rlabel metal3 25760 29176 25760 29176 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_5_.Q
rlabel metal2 32816 29960 32816 29960 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_6_.Q
rlabel metal3 37660 30744 37660 30744 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_7_.Q
rlabel metal2 37016 27272 37016 27272 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_8_.Q
rlabel metal2 38192 27608 38192 27608 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_9_.Q
rlabel metal3 46648 25256 46648 25256 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_0_.Q
rlabel metal3 42056 25032 42056 25032 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_1_.Q
rlabel metal3 52472 26376 52472 26376 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_2_.Q
rlabel metal2 40880 24024 40880 24024 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_3_.Q
rlabel metal2 37184 27384 37184 27384 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_4_.Q
rlabel metal2 40600 25592 40600 25592 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_5_.Q
rlabel metal2 42952 19376 42952 19376 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_6_.Q
rlabel metal2 45752 20048 45752 20048 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_7_.Q
rlabel metal2 44352 26824 44352 26824 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_8_.Q
rlabel metal2 45080 26656 45080 26656 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_9_.Q
rlabel metal2 58800 25592 58800 25592 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_0_.Q
rlabel metal2 50680 21224 50680 21224 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_1_.Q
rlabel metal2 49672 19432 49672 19432 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_2_.Q
rlabel metal3 42728 15960 42728 15960 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_3_.Q
rlabel metal2 47096 17976 47096 17976 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_4_.Q
rlabel metal2 46144 16968 46144 16968 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_5_.Q
rlabel metal3 47824 17528 47824 17528 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_6_.Q
rlabel metal2 53928 21168 53928 21168 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_7_.Q
rlabel metal2 54824 21336 54824 21336 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_8_.Q
rlabel metal2 51744 18536 51744 18536 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_9_.Q
rlabel metal2 58520 22568 58520 22568 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_0_.Q
rlabel metal3 53480 20664 53480 20664 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_1_.Q
rlabel metal2 52584 20748 52584 20748 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_2_.Q
rlabel metal3 57512 21672 57512 21672 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_3_.Q
rlabel metal2 56280 22904 56280 22904 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_4_.Q
rlabel metal2 61432 24640 61432 24640 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_5_.Q
rlabel metal3 57680 24808 57680 24808 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_6_.Q
rlabel metal2 62552 26488 62552 26488 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_7_.Q
rlabel metal2 56280 27608 56280 27608 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_8_.Q
rlabel metal2 61432 26544 61432 26544 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_9_.Q
rlabel metal3 54572 26488 54572 26488 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_0_.Q
rlabel metal2 48440 24696 48440 24696 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_1_.Q
rlabel metal3 57848 25424 57848 25424 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_2_.Q
rlabel metal2 61432 29176 61432 29176 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_3_.Q
rlabel metal2 62552 29512 62552 29512 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_4_.Q
rlabel metal2 62440 30912 62440 30912 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_5_.Q
rlabel metal3 62552 28448 62552 28448 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_6_.Q
rlabel metal2 62552 31472 62552 31472 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_7_.Q
rlabel metal2 65576 31584 65576 31584 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_8_.Q
rlabel metal2 2072 24976 2072 24976 0 net1
rlabel metal2 56616 64120 56616 64120 0 net10
rlabel metal2 49336 46312 49336 46312 0 net100
rlabel metal2 12208 21560 12208 21560 0 net101
rlabel metal3 41496 31080 41496 31080 0 net102
rlabel metal3 26712 27944 26712 27944 0 net103
rlabel metal2 49448 46256 49448 46256 0 net104
rlabel metal2 4088 21560 4088 21560 0 net105
rlabel metal2 5208 35448 5208 35448 0 net106
rlabel metal2 57064 42784 57064 42784 0 net107
rlabel metal3 5320 19320 5320 19320 0 net108
rlabel metal3 21112 37968 21112 37968 0 net109
rlabel metal2 44408 2030 44408 2030 0 net11
rlabel metal2 53704 39872 53704 39872 0 net110
rlabel metal2 34664 19656 34664 19656 0 net111
rlabel metal2 53144 44016 53144 44016 0 net112
rlabel metal2 26712 42336 26712 42336 0 net113
rlabel metal2 22344 18704 22344 18704 0 net114
rlabel metal2 41384 20384 41384 20384 0 net115
rlabel metal2 3976 34048 3976 34048 0 net116
rlabel metal2 3360 26152 3360 26152 0 net117
rlabel metal3 49448 43848 49448 43848 0 net118
rlabel metal2 21336 47376 21336 47376 0 net119
rlabel metal2 33824 27608 33824 27608 0 net12
rlabel metal2 21336 45584 21336 45584 0 net120
rlabel metal3 49784 23128 49784 23128 0 net121
rlabel metal3 17304 19320 17304 19320 0 net122
rlabel metal3 33936 52248 33936 52248 0 net123
rlabel metal2 10024 19264 10024 19264 0 net124
rlabel metal2 53032 43176 53032 43176 0 net125
rlabel metal2 53256 36512 53256 36512 0 net126
rlabel metal2 17864 21336 17864 21336 0 net127
rlabel metal2 9912 30464 9912 30464 0 net128
rlabel metal2 53256 21896 53256 21896 0 net129
rlabel metal2 41832 43232 41832 43232 0 net13
rlabel metal2 32032 38024 32032 38024 0 net130
rlabel metal2 53144 46536 53144 46536 0 net131
rlabel metal2 38696 34384 38696 34384 0 net132
rlabel metal2 21784 23520 21784 23520 0 net133
rlabel metal2 25368 23968 25368 23968 0 net134
rlabel metal2 53256 31808 53256 31808 0 net135
rlabel metal2 52920 46312 52920 46312 0 net136
rlabel metal2 55664 46648 55664 46648 0 net137
rlabel metal2 53256 42224 53256 42224 0 net138
rlabel metal2 14448 44408 14448 44408 0 net139
rlabel metal3 26824 38136 26824 38136 0 net14
rlabel metal2 45192 30800 45192 30800 0 net140
rlabel metal2 41552 19320 41552 19320 0 net141
rlabel metal2 27664 50680 27664 50680 0 net142
rlabel metal2 4200 29232 4200 29232 0 net143
rlabel metal2 24920 44632 24920 44632 0 net144
rlabel metal2 22904 48104 22904 48104 0 net145
rlabel metal2 16408 25480 16408 25480 0 net146
rlabel metal2 34552 39536 34552 39536 0 net147
rlabel metal2 53704 21056 53704 21056 0 net148
rlabel metal3 18368 46536 18368 46536 0 net149
rlabel metal3 26936 36568 26936 36568 0 net15
rlabel metal2 11032 20776 11032 20776 0 net150
rlabel metal3 46648 44184 46648 44184 0 net151
rlabel metal2 61544 40040 61544 40040 0 net152
rlabel metal2 64344 31640 64344 31640 0 net153
rlabel metal2 30016 31752 30016 31752 0 net154
rlabel metal2 36120 24920 36120 24920 0 net155
rlabel metal2 53480 25200 53480 25200 0 net156
rlabel metal2 40488 46592 40488 46592 0 net157
rlabel metal2 7896 37296 7896 37296 0 net158
rlabel metal3 41664 24920 41664 24920 0 net159
rlabel metal2 33544 36512 33544 36512 0 net16
rlabel metal2 57624 39144 57624 39144 0 net160
rlabel metal2 5208 33936 5208 33936 0 net161
rlabel metal2 35560 35840 35560 35840 0 net162
rlabel metal2 5208 32312 5208 32312 0 net163
rlabel metal2 15008 25592 15008 25592 0 net164
rlabel metal2 53368 36512 53368 36512 0 net165
rlabel metal3 53480 21672 53480 21672 0 net166
rlabel metal2 32088 44968 32088 44968 0 net167
rlabel metal2 8008 38528 8008 38528 0 net168
rlabel metal2 45416 20328 45416 20328 0 net169
rlabel metal2 33432 27944 33432 27944 0 net17
rlabel metal2 40040 21336 40040 21336 0 net170
rlabel metal2 38976 25480 38976 25480 0 net171
rlabel metal2 41272 21448 41272 21448 0 net172
rlabel metal2 13048 40320 13048 40320 0 net173
rlabel metal2 37408 42728 37408 42728 0 net174
rlabel metal2 22680 24752 22680 24752 0 net175
rlabel metal2 36848 51240 36848 51240 0 net176
rlabel metal2 53200 30968 53200 30968 0 net177
rlabel metal3 12768 20664 12768 20664 0 net178
rlabel metal2 34272 40376 34272 40376 0 net179
rlabel metal2 30856 27832 30856 27832 0 net18
rlabel metal2 38024 53816 38024 53816 0 net180
rlabel metal2 30128 51240 30128 51240 0 net181
rlabel metal2 4088 26376 4088 26376 0 net182
rlabel metal2 26992 26936 26992 26936 0 net183
rlabel metal3 26656 32984 26656 32984 0 net184
rlabel metal3 30408 49896 30408 49896 0 net185
rlabel metal2 45528 45584 45528 45584 0 net186
rlabel metal2 41496 50512 41496 50512 0 net187
rlabel metal2 23464 46592 23464 46592 0 net188
rlabel metal2 39032 49840 39032 49840 0 net189
rlabel metal2 32088 24584 32088 24584 0 net19
rlabel metal2 19544 18760 19544 18760 0 net190
rlabel metal2 43960 27552 43960 27552 0 net191
rlabel metal3 29512 53816 29512 53816 0 net192
rlabel metal2 37576 29176 37576 29176 0 net193
rlabel metal2 22232 37352 22232 37352 0 net194
rlabel metal3 18200 36512 18200 36512 0 net195
rlabel metal2 23800 44912 23800 44912 0 net196
rlabel metal3 6244 31864 6244 31864 0 net197
rlabel metal2 45416 30632 45416 30632 0 net198
rlabel metal3 22260 39592 22260 39592 0 net199
rlabel metal2 2072 36064 2072 36064 0 net2
rlabel metal3 30296 25592 30296 25592 0 net20
rlabel metal2 24136 20440 24136 20440 0 net200
rlabel metal2 20216 30744 20216 30744 0 net201
rlabel metal2 53032 48216 53032 48216 0 net202
rlabel metal2 51912 23856 51912 23856 0 net203
rlabel metal2 45416 38136 45416 38136 0 net204
rlabel metal3 21784 41160 21784 41160 0 net205
rlabel metal2 3976 24752 3976 24752 0 net206
rlabel metal3 47880 28560 47880 28560 0 net207
rlabel metal2 45304 36232 45304 36232 0 net208
rlabel metal2 24696 50680 24696 50680 0 net209
rlabel metal2 34664 22904 34664 22904 0 net21
rlabel metal3 11928 39704 11928 39704 0 net210
rlabel metal2 7896 31528 7896 31528 0 net211
rlabel metal2 47096 33712 47096 33712 0 net212
rlabel metal2 24864 17752 24864 17752 0 net213
rlabel metal2 20888 47544 20888 47544 0 net214
rlabel metal2 3864 24640 3864 24640 0 net215
rlabel metal3 34216 48776 34216 48776 0 net216
rlabel metal2 19768 19768 19768 19768 0 net217
rlabel metal2 19432 19936 19432 19936 0 net218
rlabel metal2 29624 24920 29624 24920 0 net219
rlabel metal2 31080 46592 31080 46592 0 net22
rlabel metal2 32424 19656 32424 19656 0 net220
rlabel metal2 44744 20776 44744 20776 0 net221
rlabel metal2 24416 29064 24416 29064 0 net222
rlabel metal2 23576 16856 23576 16856 0 net223
rlabel metal2 23296 14616 23296 14616 0 net224
rlabel metal3 44688 38472 44688 38472 0 net225
rlabel metal2 5992 20860 5992 20860 0 net226
rlabel metal3 50372 41944 50372 41944 0 net227
rlabel metal2 54432 38696 54432 38696 0 net228
rlabel metal2 19656 18312 19656 18312 0 net229
rlabel metal2 33600 53816 33600 53816 0 net23
rlabel metal2 13776 30968 13776 30968 0 net230
rlabel metal2 25592 48440 25592 48440 0 net231
rlabel metal3 28672 37240 28672 37240 0 net232
rlabel metal2 5208 37184 5208 37184 0 net233
rlabel metal2 11928 39648 11928 39648 0 net234
rlabel metal2 60368 26152 60368 26152 0 net235
rlabel metal3 33544 30128 33544 30128 0 net236
rlabel metal2 27048 51240 27048 51240 0 net237
rlabel metal3 35840 26712 35840 26712 0 net238
rlabel metal2 57624 24976 57624 24976 0 net239
rlabel metal2 32144 52248 32144 52248 0 net24
rlabel metal2 4088 28280 4088 28280 0 net240
rlabel metal3 57400 27048 57400 27048 0 net241
rlabel metal2 25816 22960 25816 22960 0 net242
rlabel metal2 18928 41832 18928 41832 0 net243
rlabel metal2 4088 23744 4088 23744 0 net244
rlabel metal2 45640 49056 45640 49056 0 net245
rlabel metal2 4200 22288 4200 22288 0 net246
rlabel metal3 39536 50568 39536 50568 0 net247
rlabel metal2 11928 40600 11928 40600 0 net248
rlabel metal3 37464 32592 37464 32592 0 net249
rlabel metal3 41496 34160 41496 34160 0 net25
rlabel metal3 51576 26152 51576 26152 0 net250
rlabel metal2 43064 51800 43064 51800 0 net251
rlabel metal2 31416 31416 31416 31416 0 net252
rlabel metal2 35056 23128 35056 23128 0 net253
rlabel metal2 7896 33600 7896 33600 0 net254
rlabel metal2 7672 23912 7672 23912 0 net255
rlabel metal2 16520 29400 16520 29400 0 net256
rlabel metal2 7896 20160 7896 20160 0 net257
rlabel metal3 17752 34944 17752 34944 0 net258
rlabel metal2 42840 19040 42840 19040 0 net259
rlabel metal3 21672 31696 21672 31696 0 net26
rlabel metal2 15064 36736 15064 36736 0 net260
rlabel metal3 28784 31864 28784 31864 0 net261
rlabel metal2 20328 47208 20328 47208 0 net262
rlabel metal3 25872 27048 25872 27048 0 net263
rlabel metal3 42728 38752 42728 38752 0 net264
rlabel metal2 26152 19376 26152 19376 0 net265
rlabel metal2 20216 44968 20216 44968 0 net266
rlabel metal2 18032 37240 18032 37240 0 net267
rlabel metal2 12600 22568 12600 22568 0 net268
rlabel metal2 46200 46368 46200 46368 0 net269
rlabel metal2 38696 31304 38696 31304 0 net27
rlabel metal2 7224 19208 7224 19208 0 net270
rlabel metal2 41160 33936 41160 33936 0 net271
rlabel metal2 4088 30240 4088 30240 0 net272
rlabel metal3 31920 48328 31920 48328 0 net273
rlabel metal2 36568 34552 36568 34552 0 net274
rlabel metal3 46536 24024 46536 24024 0 net28
rlabel metal3 20916 37240 20916 37240 0 net29
rlabel metal3 62608 30968 62608 30968 0 net3
rlabel metal3 45416 33208 45416 33208 0 net30
rlabel metal2 15848 42672 15848 42672 0 net31
rlabel metal2 8008 34944 8008 34944 0 net32
rlabel metal2 60424 33656 60424 33656 0 net33
rlabel metal2 3864 34160 3864 34160 0 net34
rlabel metal3 45416 27104 45416 27104 0 net35
rlabel metal2 50904 49616 50904 49616 0 net36
rlabel metal2 51800 48944 51800 48944 0 net37
rlabel metal2 23128 43624 23128 43624 0 net38
rlabel metal2 27216 14616 27216 14616 0 net39
rlabel metal2 66248 62720 66248 62720 0 net4
rlabel metal2 49448 44856 49448 44856 0 net40
rlabel metal2 37408 23912 37408 23912 0 net41
rlabel metal2 45976 23520 45976 23520 0 net42
rlabel metal2 14392 16184 14392 16184 0 net43
rlabel metal2 54152 44128 54152 44128 0 net44
rlabel metal3 42056 42840 42056 42840 0 net45
rlabel metal3 8204 37128 8204 37128 0 net46
rlabel metal2 29624 21672 29624 21672 0 net47
rlabel metal2 3976 27720 3976 27720 0 net48
rlabel metal2 23688 47544 23688 47544 0 net49
rlabel metal2 40376 2030 40376 2030 0 net5
rlabel metal2 19768 18088 19768 18088 0 net50
rlabel metal3 45136 24136 45136 24136 0 net51
rlabel metal3 45920 43960 45920 43960 0 net52
rlabel metal2 6216 20048 6216 20048 0 net53
rlabel metal3 40936 39704 40936 39704 0 net54
rlabel metal2 38976 21560 38976 21560 0 net55
rlabel metal3 53956 22456 53956 22456 0 net56
rlabel metal2 41608 38920 41608 38920 0 net57
rlabel metal2 35728 52248 35728 52248 0 net58
rlabel metal3 55944 30912 55944 30912 0 net59
rlabel metal2 48440 2030 48440 2030 0 net6
rlabel metal2 45472 47432 45472 47432 0 net60
rlabel metal2 25368 38584 25368 38584 0 net61
rlabel metal2 42280 26264 42280 26264 0 net62
rlabel metal2 47656 35224 47656 35224 0 net63
rlabel metal2 44464 18312 44464 18312 0 net64
rlabel metal2 49224 38192 49224 38192 0 net65
rlabel metal2 45416 22176 45416 22176 0 net66
rlabel metal2 34384 27160 34384 27160 0 net67
rlabel metal3 37072 52808 37072 52808 0 net68
rlabel metal2 53256 28168 53256 28168 0 net69
rlabel metal2 41048 2030 41048 2030 0 net7
rlabel metal2 53144 33880 53144 33880 0 net70
rlabel metal2 44968 51576 44968 51576 0 net71
rlabel metal2 41384 23744 41384 23744 0 net72
rlabel metal2 7112 30464 7112 30464 0 net73
rlabel metal2 15680 16744 15680 16744 0 net74
rlabel metal2 11816 21392 11816 21392 0 net75
rlabel metal3 36120 32648 36120 32648 0 net76
rlabel metal2 60424 41496 60424 41496 0 net77
rlabel metal3 49868 29400 49868 29400 0 net78
rlabel metal2 53704 22064 53704 22064 0 net79
rlabel metal2 54488 2030 54488 2030 0 net8
rlabel metal3 42112 44968 42112 44968 0 net80
rlabel metal2 40152 21000 40152 21000 0 net81
rlabel metal3 40544 49000 40544 49000 0 net82
rlabel metal2 49336 34216 49336 34216 0 net83
rlabel metal2 57736 24920 57736 24920 0 net84
rlabel metal2 55608 29736 55608 29736 0 net85
rlabel metal2 50680 37184 50680 37184 0 net86
rlabel metal2 31864 30296 31864 30296 0 net87
rlabel metal2 12712 25928 12712 25928 0 net88
rlabel metal2 39872 48664 39872 48664 0 net89
rlabel metal2 43736 2030 43736 2030 0 net9
rlabel metal2 47768 47656 47768 47656 0 net90
rlabel metal2 11032 23352 11032 23352 0 net91
rlabel metal2 16856 42224 16856 42224 0 net92
rlabel metal4 54040 39984 54040 39984 0 net93
rlabel metal2 51128 34216 51128 34216 0 net94
rlabel metal2 37632 27048 37632 27048 0 net95
rlabel metal2 49224 50120 49224 50120 0 net96
rlabel metal3 29344 18536 29344 18536 0 net97
rlabel metal2 44744 50232 44744 50232 0 net98
rlabel metal2 50232 39424 50232 39424 0 net99
rlabel metal3 1246 36344 1246 36344 0 pReset
rlabel metal3 2478 47768 2478 47768 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 68000 68000
<< end >>
