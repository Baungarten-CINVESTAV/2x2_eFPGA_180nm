// This is the unpowered netlist.
module sb_0__2_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
 input [19:0] chanx_right_in;
 output [19:0] chanx_right_out;
 input [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;

 wire net59;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net47;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire clknet_0_prog_clk;
 wire clknet_2_0__leaf_prog_clk;
 wire clknet_2_1__leaf_prog_clk;
 wire clknet_2_2__leaf_prog_clk;
 wire clknet_2_3__leaf_prog_clk;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_11.DFFR_0_.D ;
 wire \mem_bottom_track_11.DFFR_0_.Q ;
 wire \mem_bottom_track_11.DFFR_1_.Q ;
 wire \mem_bottom_track_21.DFFR_0_.Q ;
 wire \mem_bottom_track_21.DFFR_1_.Q ;
 wire \mem_bottom_track_23.DFFR_0_.Q ;
 wire \mem_bottom_track_23.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_27.DFFR_0_.Q ;
 wire \mem_bottom_track_27.DFFR_1_.Q ;
 wire \mem_bottom_track_29.DFFR_0_.Q ;
 wire \mem_bottom_track_29.DFFR_1_.Q ;
 wire \mem_bottom_track_3.DFFR_0_.Q ;
 wire \mem_bottom_track_3.DFFR_1_.Q ;
 wire \mem_bottom_track_31.DFFR_0_.Q ;
 wire \mem_bottom_track_5.DFFR_0_.Q ;
 wire \mem_bottom_track_5.DFFR_1_.Q ;
 wire \mem_bottom_track_7.DFFR_0_.Q ;
 wire \mem_bottom_track_7.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_10.DFFR_0_.D ;
 wire \mem_right_track_10.DFFR_0_.Q ;
 wire \mem_right_track_10.DFFR_1_.Q ;
 wire \mem_right_track_2.DFFR_0_.Q ;
 wire \mem_right_track_2.DFFR_1_.Q ;
 wire \mem_right_track_20.DFFR_0_.Q ;
 wire \mem_right_track_20.DFFR_1_.Q ;
 wire \mem_right_track_22.DFFR_0_.Q ;
 wire \mem_right_track_22.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_26.DFFR_0_.Q ;
 wire \mem_right_track_26.DFFR_1_.Q ;
 wire \mem_right_track_28.DFFR_0_.Q ;
 wire \mem_right_track_28.DFFR_1_.Q ;
 wire \mem_right_track_30.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_1_.Q ;
 wire \mem_right_track_6.DFFR_0_.Q ;
 wire \mem_right_track_6.DFFR_1_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net4;
 wire net5;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__054__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__055__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__056__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__057__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__058__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__059__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__060__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__061__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__062__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__063__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__064__I (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__065__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__089__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__091__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__092__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__093__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__094__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__095__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__096__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__097__I (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__100__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__I (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__116__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__122__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__CLK (.I(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(chany_bottom_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(chany_bottom_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(chany_bottom_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(chany_bottom_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(chany_bottom_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(chany_bottom_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(chany_bottom_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(chany_bottom_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(chanx_right_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(chanx_right_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(chanx_right_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(chanx_right_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(chanx_right_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(chanx_right_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(chanx_right_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(chanx_right_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_93 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _053_ (.I(net18),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _054_ (.I(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _055_ (.I(_049_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _056_ (.I(_049_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _057_ (.I(_049_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _058_ (.I(_049_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _059_ (.I(_049_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _060_ (.I(_049_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _061_ (.I(_049_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _062_ (.I(_049_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _063_ (.I(_049_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _064_ (.I(_049_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _065_ (.I(_048_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _066_ (.I(_050_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _067_ (.I(_050_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _068_ (.I(_050_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _069_ (.I(_050_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _070_ (.I(_050_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _071_ (.I(_050_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _072_ (.I(_050_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _073_ (.I(_050_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _074_ (.I(_050_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _075_ (.I(_050_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _076_ (.I(net18),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _077_ (.I(_051_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _078_ (.I(_051_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _079_ (.I(_051_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _080_ (.I(_051_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _081_ (.I(_051_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _082_ (.I(_051_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _083_ (.I(_051_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _084_ (.I(_051_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _085_ (.I(_051_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _086_ (.I(_051_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _087_ (.I(net18),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _088_ (.I(_052_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _089_ (.I(_052_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _090_ (.I(_052_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _091_ (.I(_052_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _092_ (.I(_052_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _093_ (.I(_052_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _094_ (.I(_052_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _095_ (.I(_052_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _096_ (.I(_052_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _097_ (.I(_052_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _098_ (.I(_048_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _099_ (.I(_048_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _100_ (.I(_048_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _101_ (.I(_048_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _102_ (.I(_048_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _103_ (.I(_048_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _104_ (.I(_048_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _105_ (.I(_048_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _106_ (.D(net83),
    .RN(_000_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _107_ (.D(net1),
    .RN(_001_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _108_ (.D(net89),
    .RN(_002_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _109_ (.D(net100),
    .RN(_003_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _110_ (.D(net95),
    .RN(_004_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _111_ (.D(net70),
    .RN(_005_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _112_ (.D(net68),
    .RN(_006_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _113_ (.D(net78),
    .RN(_007_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _114_ (.D(net71),
    .RN(_008_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_10.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _115_ (.D(net102),
    .RN(_009_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _116_ (.D(net80),
    .RN(_010_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_10.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _117_ (.D(net63),
    .RN(_011_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_10.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _118_ (.D(net92),
    .RN(_012_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_20.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _119_ (.D(net84),
    .RN(_013_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_20.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _120_ (.D(net73),
    .RN(_014_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_22.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _121_ (.D(net93),
    .RN(_015_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_22.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _122_ (.D(net98),
    .RN(_016_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _123_ (.D(net105),
    .RN(_017_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _124_ (.D(net60),
    .RN(_018_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_track_26.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _125_ (.D(net106),
    .RN(_019_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_track_26.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _126_ (.D(net65),
    .RN(_020_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_right_track_28.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _127_ (.D(net97),
    .RN(_021_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_track_28.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _128_ (.D(net79),
    .RN(_022_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _129_ (.D(net61),
    .RN(_023_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_track_30.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _130_ (.D(net82),
    .RN(_024_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _131_ (.D(net87),
    .RN(_025_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _132_ (.D(net85),
    .RN(_026_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_3.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _133_ (.D(net94),
    .RN(_027_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_3.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _134_ (.D(net91),
    .RN(_028_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_5.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _135_ (.D(net81),
    .RN(_029_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_5.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _136_ (.D(net69),
    .RN(_030_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_7.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _137_ (.D(net76),
    .RN(_031_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_7.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _138_ (.D(net74),
    .RN(_032_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_11.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _139_ (.D(net64),
    .RN(_033_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _140_ (.D(net75),
    .RN(_034_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_11.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _141_ (.D(net90),
    .RN(_035_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_11.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _142_ (.D(net96),
    .RN(_036_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_21.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _143_ (.D(net88),
    .RN(_037_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_21.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _144_ (.D(net103),
    .RN(_038_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_23.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _145_ (.D(net101),
    .RN(_039_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_23.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _146_ (.D(net104),
    .RN(_040_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _147_ (.D(net86),
    .RN(_041_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _148_ (.D(net62),
    .RN(_042_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_27.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _149_ (.D(net67),
    .RN(_043_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_bottom_track_27.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _150_ (.D(net66),
    .RN(_044_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_bottom_track_29.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _151_ (.D(net77),
    .RN(_045_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_bottom_track_29.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _152_ (.D(net99),
    .RN(_046_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _153_ (.D(net72),
    .RN(_047_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_bottom_track_31.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _178_ (.I(net14),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _179_ (.I(net10),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _180_ (.I(net15),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _181_ (.I(net16),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _182_ (.I(net17),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _183_ (.I(net11),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _184_ (.I(net12),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _185_ (.I(net13),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _186_ (.I(net6),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _187_ (.I(net2),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _188_ (.I(net7),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _189_ (.I(net8),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _190_ (.I(net9),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _191_ (.I(net3),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _192_ (.I(net4),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _193_ (.I(net5),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\mem_right_track_26.DFFR_0_.Q ),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\mem_bottom_track_7.DFFR_0_.Q ),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\mem_right_track_2.DFFR_1_.Q ),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\mem_right_track_8.DFFR_0_.Q ),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\mem_bottom_track_29.DFFR_1_.Q ),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\mem_right_track_22.DFFR_0_.Q ),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\mem_bottom_track_9.DFFR_0_.Q ),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\mem_bottom_track_11.DFFR_0_.Q ),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\mem_bottom_track_5.DFFR_1_.Q ),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\mem_bottom_track_27.DFFR_1_.Q ),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\mem_right_track_4.DFFR_1_.Q ),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\mem_right_track_28.DFFR_1_.Q ),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\mem_right_track_30.DFFR_0_.Q ),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\mem_right_track_10.DFFR_0_.Q ),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\mem_bottom_track_3.DFFR_1_.Q ),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\mem_bottom_track_1.DFFR_0_.Q ),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\mem_right_track_0.DFFR_0_.Q ),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\mem_right_track_10.DFFR_1_.Q ),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\mem_bottom_track_3.DFFR_0_.Q ),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\mem_bottom_track_23.DFFR_1_.Q ),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\mem_bottom_track_1.DFFR_0_.D ),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\mem_bottom_track_11.DFFR_1_.Q ),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\mem_bottom_track_27.DFFR_0_.Q ),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\mem_right_track_2.DFFR_0_.Q ),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\mem_bottom_track_11.DFFR_0_.D ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\mem_bottom_track_5.DFFR_0_.Q ),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\mem_right_track_20.DFFR_0_.Q ),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\mem_right_track_20.DFFR_1_.Q ),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\mem_bottom_track_1.DFFR_1_.Q ),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\mem_right_track_4.DFFR_0_.Q ),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\mem_bottom_track_21.DFFR_0_.Q ),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\mem_right_track_26.DFFR_1_.Q ),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\mem_right_track_24.DFFR_0_.Q ),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\mem_right_track_10.DFFR_0_.D ),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\mem_bottom_track_31.DFFR_0_.Q ),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\mem_right_track_0.DFFR_1_.Q ),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\mem_bottom_track_21.DFFR_1_.Q ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\mem_right_track_6.DFFR_1_.Q ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\mem_bottom_track_23.DFFR_0_.Q ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\mem_bottom_track_25.DFFR_0_.Q ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\mem_right_track_22.DFFR_1_.Q ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\mem_right_track_24.DFFR_1_.Q ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\mem_bottom_track_7.DFFR_1_.Q ),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\mem_right_track_28.DFFR_0_.Q ),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\mem_bottom_track_29.DFFR_0_.Q ),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\mem_bottom_track_25.DFFR_1_.Q ),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\mem_right_track_6.DFFR_0_.Q ),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(chany_bottom_in[0]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(chany_bottom_in[10]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(chany_bottom_in[11]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(chany_bottom_in[12]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(chany_bottom_in[19]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(chany_bottom_in[1]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(chany_bottom_in[2]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(chany_bottom_in[9]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(pReset),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(chanx_right_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(chanx_right_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(chanx_right_in[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(chanx_right_in[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(chanx_right_in[19]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(chanx_right_in[1]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(chanx_right_in[2]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(chanx_right_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output19 (.I(net19),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output20 (.I(net20),
    .Z(chanx_right_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output21 (.I(net21),
    .Z(chanx_right_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output22 (.I(net22),
    .Z(chanx_right_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output23 (.I(net23),
    .Z(chanx_right_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output24 (.I(net24),
    .Z(chanx_right_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output25 (.I(net25),
    .Z(chanx_right_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(chanx_right_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output27 (.I(net27),
    .Z(chanx_right_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(chany_bottom_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output29 (.I(net29),
    .Z(chany_bottom_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output30 (.I(net30),
    .Z(chany_bottom_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output31 (.I(net31),
    .Z(chany_bottom_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output32 (.I(net32),
    .Z(chany_bottom_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output33 (.I(net33),
    .Z(chany_bottom_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output34 (.I(net34),
    .Z(chany_bottom_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output35 (.I(net35),
    .Z(chany_bottom_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__2__59 (.ZN(net59));
 assign chanx_right_out[0] = net59;
 assign chanx_right_out[10] = net53;
 assign chanx_right_out[11] = net52;
 assign chanx_right_out[12] = net51;
 assign chanx_right_out[13] = net50;
 assign chanx_right_out[14] = net49;
 assign chanx_right_out[15] = net48;
 assign chanx_right_out[1] = net58;
 assign chanx_right_out[2] = net57;
 assign chanx_right_out[3] = net56;
 assign chanx_right_out[4] = net55;
 assign chanx_right_out[5] = net54;
 assign chany_bottom_out[0] = net47;
 assign chany_bottom_out[10] = net41;
 assign chany_bottom_out[11] = net40;
 assign chany_bottom_out[12] = net39;
 assign chany_bottom_out[13] = net38;
 assign chany_bottom_out[14] = net37;
 assign chany_bottom_out[15] = net36;
 assign chany_bottom_out[1] = net46;
 assign chany_bottom_out[2] = net45;
 assign chany_bottom_out[3] = net44;
 assign chany_bottom_out[4] = net43;
 assign chany_bottom_out[5] = net42;
endmodule

