* NGSPICE file created from sb_2__0_.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

.subckt sb_2__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
+ pReset prog_clk top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ vdd vss chanx_left_out[14] chanx_left_out[15] chany_top_out[0] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13]
XFILLER_0_7_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__140__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_131_ net87 _025_ clknet_2_1__leaf_prog_clk mem_left_track_1.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_062_ _049_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_28_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_114_ net71 _008_ clknet_2_0__leaf_prog_clk mem_top_track_10.DFFR_0_.D vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold30 mem_top_track_2.DFFR_0_.Q net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold41 mem_top_track_0.DFFR_1_.Q net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput31 net31 chany_top_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput20 net20 chanx_left_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__090__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_130_ net82 _024_ clknet_2_1__leaf_prog_clk mem_left_track_1.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_061_ _049_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__153__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_113_ net78 _007_ clknet_2_0__leaf_prog_clk mem_top_track_6.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold42 mem_left_track_21.DFFR_1_.Q net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold31 mem_left_track_11.DFFR_0_.D net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_15_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold20 mem_top_track_30.DFFR_0_.Q net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I chany_top_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__093__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput32 net32 chany_top_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput21 net21 chanx_left_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__088__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I chanx_left_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_060_ _049_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_189_ net9 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__096__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_112_ net68 _006_ clknet_2_0__leaf_prog_clk mem_top_track_6.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__120__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__143__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold10 mem_left_track_7.DFFR_0_.Q net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold32 mem_left_track_5.DFFR_0_.Q net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold43 mem_top_track_6.DFFR_1_.Q net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold21 mem_top_track_10.DFFR_0_.Q net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net33 chany_top_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput22 net22 chanx_left_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__099__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_188_ net8 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_24_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_111_ net70 _005_ clknet_2_0__leaf_prog_clk mem_top_track_4.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_21_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold22 mem_left_track_3.DFFR_1_.Q net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold11 mem_top_track_2.DFFR_1_.Q net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 mem_top_track_20.DFFR_0_.Q net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold44 mem_left_track_23.DFFR_0_.Q net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_16_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput34 net34 chany_top_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput23 net23 chanx_left_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_11_Left_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_187_ net7 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_110_ net95 _004_ clknet_2_0__leaf_prog_clk mem_top_track_4.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold45 mem_left_track_25.DFFR_0_.Q net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold23 mem_left_track_1.DFFR_0_.Q net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 mem_top_track_20.DFFR_1_.Q net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold12 mem_top_track_8.DFFR_0_.Q net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_2_3__f_prog_clk clknet_0_prog_clk clknet_2_3__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput24 net24 chanx_left_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput35 net35 chany_top_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I ccff_head vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__123__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_186_ net6 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2__f_prog_clk clknet_0_prog_clk clknet_2_2__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold13 mem_left_track_29.DFFR_1_.Q net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold35 mem_left_track_1.DFFR_1_.Q net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 mem_top_track_22.DFFR_1_.Q net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold24 mem_top_track_0.DFFR_0_.Q net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__102__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 chanx_left_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_185_ net13 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_2_1__f_prog_clk clknet_0_prog_clk clknet_2_1__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__105__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_099_ _048_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold14 mem_top_track_22.DFFR_0_.Q net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 mem_top_track_10.DFFR_1_.Q net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold36 mem_top_track_4.DFFR_0_.Q net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold47 mem_top_track_24.DFFR_1_.Q net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_29_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput26 net26 chanx_left_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_0__f_prog_clk clknet_0_prog_clk clknet_2_0__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_184_ net12 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_098_ _048_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_3_Left_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold37 mem_left_track_21.DFFR_0_.Q net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold15 mem_left_track_9.DFFR_0_.Q net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold26 mem_left_track_3.DFFR_0_.Q net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_10_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput27 net27 chanx_left_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_183_ net11 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_097_ _052_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold16 mem_left_track_11.DFFR_0_.Q net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I pReset vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold27 mem_left_track_23.DFFR_1_.Q net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold38 mem_top_track_26.DFFR_1_.Q net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_10_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_149_ net67 _043_ clknet_2_1__leaf_prog_clk mem_left_track_27.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_16_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput28 net28 chany_top_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__116__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__139__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_182_ net10 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_096_ _052_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold17 mem_left_track_5.DFFR_1_.Q net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 mem_left_track_1.DFFR_0_.D net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold39 mem_top_track_24.DFFR_0_.Q net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_10_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_148_ net62 _042_ clknet_2_3__leaf_prog_clk mem_left_track_27.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput29 net29 chany_top_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_079_ _051_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_19_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_181_ net17 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__061__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_095_ _052_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold29 mem_left_track_11.DFFR_1_.Q net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold18 mem_left_track_27.DFFR_1_.Q net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__129__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__056__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_147_ net86 _041_ clknet_2_3__leaf_prog_clk mem_left_track_25.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_7_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_078_ _051_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput19 net19 ccff_tail vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__064__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__059__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_180_ net16 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_094_ _052_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_23_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold19 mem_top_track_4.DFFR_1_.Q net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_29_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_146_ net104 _040_ clknet_2_1__leaf_prog_clk mem_left_track_25.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_077_ _051_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input16_I chany_top_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__119__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I chanx_left_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_129_ net61 _023_ clknet_2_3__leaf_prog_clk mem_top_track_30.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_10_Left_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_2__0__50 chanx_left_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_093_ _052_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__152__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_prog_clk prog_clk clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput1 ccff_head net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_29_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_076_ net18 _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_145_ net101 _039_ clknet_2_3__leaf_prog_clk mem_left_track_23.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_17_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_128_ net79 _022_ clknet_2_1__leaf_prog_clk mem_left_track_1.DFFR_0_.D vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_059_ _049_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_22_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__091__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_2__0__51 chanx_left_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__40 chany_top_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_092_ _052_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput2 chanx_left_in[11] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_144_ net103 _038_ clknet_2_3__leaf_prog_clk mem_left_track_23.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_075_ _050_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__142__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_058_ _049_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_127_ net97 _021_ clknet_2_0__leaf_prog_clk mem_top_track_28.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_22_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__094__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__089__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsb_2__0__52 chanx_left_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__41 chany_top_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_091_ _052_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__097__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 chanx_left_in[12] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_143_ net88 _037_ clknet_2_3__leaf_prog_clk mem_left_track_21.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_074_ _050_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_27_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_126_ net65 _020_ clknet_2_1__leaf_prog_clk mem_top_track_28.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_057_ _049_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input14_I chany_top_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input6_I chanx_left_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_109_ net100 _003_ clknet_2_0__leaf_prog_clk mem_top_track_2.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_27_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xsb_2__0__53 chanx_left_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__42 chany_top_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_090_ _052_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput4 chanx_left_in[13] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_142_ net96 _036_ clknet_2_3__leaf_prog_clk mem_left_track_21.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_073_ _050_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_125_ net106 _019_ clknet_2_2__leaf_prog_clk mem_top_track_26.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_056_ _049_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_108_ net89 _002_ clknet_2_0__leaf_prog_clk mem_top_track_2.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsb_2__0__54 chanx_left_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__122__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_2__0__43 chany_top_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__145__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 chanx_left_in[14] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_141_ net90 _035_ clknet_2_3__leaf_prog_clk mem_left_track_11.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_072_ _050_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_124_ net60 _018_ clknet_2_3__leaf_prog_clk mem_top_track_26.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_055_ _049_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_107_ net1 _001_ clknet_2_0__leaf_prog_clk mem_top_track_0.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsb_2__0__55 chanx_left_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__100__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_2__0__44 chany_top_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput6 chanx_left_in[1] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_140_ net75 _034_ clknet_2_3__leaf_prog_clk mem_left_track_11.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_071_ _050_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_123_ net105 _017_ clknet_2_2__leaf_prog_clk mem_top_track_24.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_054_ _048_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__103__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_106_ net83 _000_ clknet_2_0__leaf_prog_clk mem_top_track_0.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_28_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I chany_top_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I chanx_left_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_2__0__45 chany_top_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__56 chanx_left_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 chanx_left_in[2] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_070_ _050_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_9_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_053_ net18 _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_122_ net98 _016_ clknet_2_2__leaf_prog_clk mem_top_track_24.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput10 chany_top_in[11] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_105_ _048_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__125__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__148__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsb_2__0__46 chany_top_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__57 chanx_left_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput8 chanx_left_in[3] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_121_ net93 _015_ clknet_2_2__leaf_prog_clk mem_top_track_22.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput11 chany_top_in[12] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_104_ _048_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_2__0__47 chany_top_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__36 chany_top_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__58 chanx_left_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__138__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 chanx_left_in[4] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_120_ net73 _014_ clknet_2_2__leaf_prog_clk mem_top_track_22.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_16_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput12 chany_top_in[13] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_103_ _048_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 mem_top_track_26.DFFR_0_.Q net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xsb_2__0__59 chanx_left_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input10_I chany_top_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_2__0__37 chany_top_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__48 chanx_left_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input2_I chanx_left_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 chany_top_in[14] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_179_ net15 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_102_ _048_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__054__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold2 mem_top_track_28.DFFR_1_.Q net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_4_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsb_2__0__38 chany_top_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__0__49 chanx_left_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__062__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__057__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput14 chany_top_in[1] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_178_ net14 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__118__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_101_ _048_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold3 mem_left_track_27.DFFR_0_.Q net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_4_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__065__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_2__0__39 chany_top_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_17_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__151__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput15 chany_top_in[2] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_100_ _048_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_21_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold4 mem_top_track_10.DFFR_0_.D net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_prog_clk_I prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_193_ net5 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__141__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 chany_top_in[3] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 mem_left_track_7.DFFR_1_.Q net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_20_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__092__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_192_ net4 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 chany_top_in[4] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__095__I _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_089_ _052_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold6 mem_top_track_28.DFFR_0_.Q net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_191_ net3 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__098__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 pReset net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_5_Left_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_088_ _052_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_12_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold7 mem_left_track_29.DFFR_0_.Q net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__121__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__144__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_190_ net2 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_087_ net18 _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input17_I chany_top_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold8 mem_left_track_25.DFFR_1_.Q net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input9_I chanx_left_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_139_ net64 _033_ clknet_2_3__leaf_prog_clk mem_left_track_9.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_28_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_086_ _051_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_12_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 mem_top_track_6.DFFR_0_.Q net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_138_ net74 _032_ clknet_2_3__leaf_prog_clk mem_left_track_11.DFFR_0_.D vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_069_ _050_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_28_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__101__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_085_ _051_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__124__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__147__CLK clknet_2_3__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__104__I _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Left_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_137_ net76 _031_ clknet_2_1__leaf_prog_clk mem_left_track_7.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_068_ _050_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_9_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_084_ _051_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_153_ net72 _047_ clknet_2_2__leaf_prog_clk mem_left_track_31.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_136_ net69 _030_ clknet_2_1__leaf_prog_clk mem_left_track_7.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_29_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_067_ _050_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input15_I chany_top_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I chanx_left_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_119_ net84 _013_ clknet_2_2__leaf_prog_clk mem_top_track_20.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_12_Left_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_083_ _051_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_0_Left_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_152_ net99 _046_ clknet_2_2__leaf_prog_clk net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_28_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_135_ net81 _029_ clknet_2_1__leaf_prog_clk mem_left_track_5.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_066_ _050_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_118_ net92 _012_ clknet_2_2__leaf_prog_clk mem_top_track_20.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_21_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_151_ net77 _045_ clknet_2_3__leaf_prog_clk mem_left_track_29.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_082_ _051_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_29_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_134_ net91 _028_ clknet_2_1__leaf_prog_clk mem_left_track_5.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_065_ _048_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_117_ net63 _011_ clknet_2_2__leaf_prog_clk mem_top_track_10.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_081_ _051_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_150_ net66 _044_ clknet_2_2__leaf_prog_clk mem_left_track_29.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__117__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__060__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_133_ net94 _027_ clknet_2_1__leaf_prog_clk mem_left_track_3.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_064_ _049_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__055__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_116_ net80 _010_ clknet_2_2__leaf_prog_clk mem_top_track_10.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input13_I chany_top_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__150__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I chanx_left_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__063__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__058__I _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_080_ _051_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_132_ net85 _026_ clknet_2_1__leaf_prog_clk mem_left_track_3.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_063_ _049_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_4_Left_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_115_ net102 _009_ clknet_2_0__leaf_prog_clk mem_top_track_8.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold40 mem_left_track_31.DFFR_0_.Q net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xoutput30 net30 chany_top_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_27_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

