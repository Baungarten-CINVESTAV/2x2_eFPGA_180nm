magic
tech gf180mcuD
magscale 1 10
timestamp 1702153875
<< metal1 >>
rect 2034 26798 2046 26850
rect 2098 26847 2110 26850
rect 2594 26847 2606 26850
rect 2098 26801 2606 26847
rect 2098 26798 2110 26801
rect 2594 26798 2606 26801
rect 2658 26798 2670 26850
rect 13458 26798 13470 26850
rect 13522 26847 13534 26850
rect 14130 26847 14142 26850
rect 13522 26801 14142 26847
rect 13522 26798 13534 26801
rect 14130 26798 14142 26801
rect 14194 26798 14206 26850
rect 18834 26798 18846 26850
rect 18898 26847 18910 26850
rect 20066 26847 20078 26850
rect 18898 26801 20078 26847
rect 18898 26798 18910 26801
rect 20066 26798 20078 26801
rect 20130 26798 20142 26850
rect 20290 26798 20302 26850
rect 20354 26847 20366 26850
rect 21186 26847 21198 26850
rect 20354 26801 21198 26847
rect 20354 26798 20366 26801
rect 21186 26798 21198 26801
rect 21250 26798 21262 26850
rect 22194 26798 22206 26850
rect 22258 26847 22270 26850
rect 22866 26847 22878 26850
rect 22258 26801 22878 26847
rect 22258 26798 22270 26801
rect 22866 26798 22878 26801
rect 22930 26798 22942 26850
rect 24210 26798 24222 26850
rect 24274 26847 24286 26850
rect 24770 26847 24782 26850
rect 24274 26801 24782 26847
rect 24274 26798 24286 26801
rect 24770 26798 24782 26801
rect 24834 26798 24846 26850
rect 1344 26682 28720 26716
rect 1344 26630 8018 26682
rect 8070 26630 8122 26682
rect 8174 26630 8226 26682
rect 8278 26630 14822 26682
rect 14874 26630 14926 26682
rect 14978 26630 15030 26682
rect 15082 26630 21626 26682
rect 21678 26630 21730 26682
rect 21782 26630 21834 26682
rect 21886 26630 28430 26682
rect 28482 26630 28534 26682
rect 28586 26630 28638 26682
rect 28690 26630 28720 26682
rect 1344 26596 28720 26630
rect 15486 26514 15538 26526
rect 15486 26450 15538 26462
rect 20078 26514 20130 26526
rect 20078 26450 20130 26462
rect 24110 26514 24162 26526
rect 24110 26450 24162 26462
rect 26126 26514 26178 26526
rect 26126 26450 26178 26462
rect 4286 26402 4338 26414
rect 2594 26350 2606 26402
rect 2658 26350 2670 26402
rect 4286 26338 4338 26350
rect 4958 26402 5010 26414
rect 15710 26402 15762 26414
rect 7858 26350 7870 26402
rect 7922 26350 7934 26402
rect 10658 26350 10670 26402
rect 10722 26350 10734 26402
rect 12226 26350 12238 26402
rect 12290 26350 12302 26402
rect 4958 26338 5010 26350
rect 15710 26338 15762 26350
rect 13694 26290 13746 26302
rect 16942 26290 16994 26302
rect 20750 26290 20802 26302
rect 24558 26290 24610 26302
rect 3378 26238 3390 26290
rect 3442 26238 3454 26290
rect 4050 26238 4062 26290
rect 4114 26238 4126 26290
rect 4722 26238 4734 26290
rect 4786 26238 4798 26290
rect 6850 26238 6862 26290
rect 6914 26238 6926 26290
rect 8530 26238 8542 26290
rect 8594 26238 8606 26290
rect 9986 26238 9998 26290
rect 10050 26238 10062 26290
rect 11330 26238 11342 26290
rect 11394 26238 11406 26290
rect 15922 26238 15934 26290
rect 15986 26238 15998 26290
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 22418 26238 22430 26290
rect 22482 26238 22494 26290
rect 26562 26238 26574 26290
rect 26626 26238 26638 26290
rect 13694 26226 13746 26238
rect 16942 26226 16994 26238
rect 20750 26226 20802 26238
rect 24558 26226 24610 26238
rect 5842 26126 5854 26178
rect 5906 26126 5918 26178
rect 14130 26126 14142 26178
rect 14194 26126 14206 26178
rect 17378 26126 17390 26178
rect 17442 26126 17454 26178
rect 18946 26126 18958 26178
rect 19010 26126 19022 26178
rect 21186 26126 21198 26178
rect 21250 26126 21262 26178
rect 22754 26126 22766 26178
rect 22818 26126 22830 26178
rect 24994 26126 25006 26178
rect 25058 26126 25070 26178
rect 27682 26126 27694 26178
rect 27746 26126 27758 26178
rect 1344 25898 28560 25932
rect 1344 25846 4616 25898
rect 4668 25846 4720 25898
rect 4772 25846 4824 25898
rect 4876 25846 11420 25898
rect 11472 25846 11524 25898
rect 11576 25846 11628 25898
rect 11680 25846 18224 25898
rect 18276 25846 18328 25898
rect 18380 25846 18432 25898
rect 18484 25846 25028 25898
rect 25080 25846 25132 25898
rect 25184 25846 25236 25898
rect 25288 25846 28560 25898
rect 1344 25812 28560 25846
rect 10558 25730 10610 25742
rect 10558 25666 10610 25678
rect 1822 25618 1874 25630
rect 1822 25554 1874 25566
rect 5070 25618 5122 25630
rect 5070 25554 5122 25566
rect 6078 25618 6130 25630
rect 6078 25554 6130 25566
rect 8766 25618 8818 25630
rect 14814 25618 14866 25630
rect 12114 25566 12126 25618
rect 12178 25566 12190 25618
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 8766 25554 8818 25566
rect 14814 25554 14866 25566
rect 16830 25618 16882 25630
rect 19630 25618 19682 25630
rect 18834 25566 18846 25618
rect 18898 25566 18910 25618
rect 16830 25554 16882 25566
rect 19630 25554 19682 25566
rect 20862 25618 20914 25630
rect 22866 25566 22878 25618
rect 22930 25566 22942 25618
rect 25890 25566 25902 25618
rect 25954 25566 25966 25618
rect 20862 25554 20914 25566
rect 3614 25506 3666 25518
rect 3614 25442 3666 25454
rect 6302 25506 6354 25518
rect 6302 25442 6354 25454
rect 6974 25506 7026 25518
rect 6974 25442 7026 25454
rect 7646 25506 7698 25518
rect 7646 25442 7698 25454
rect 8990 25506 9042 25518
rect 15038 25506 15090 25518
rect 21310 25506 21362 25518
rect 11778 25454 11790 25506
rect 11842 25454 11854 25506
rect 17266 25454 17278 25506
rect 17330 25454 17342 25506
rect 18498 25454 18510 25506
rect 18562 25454 18574 25506
rect 20178 25454 20190 25506
rect 20242 25454 20254 25506
rect 8990 25442 9042 25454
rect 15038 25442 15090 25454
rect 21310 25442 21362 25454
rect 23662 25506 23714 25518
rect 24210 25454 24222 25506
rect 24274 25454 24286 25506
rect 24882 25454 24894 25506
rect 24946 25454 24958 25506
rect 23662 25442 23714 25454
rect 3950 25394 4002 25406
rect 3950 25330 4002 25342
rect 4286 25394 4338 25406
rect 4286 25330 4338 25342
rect 6638 25394 6690 25406
rect 6638 25330 6690 25342
rect 7310 25394 7362 25406
rect 7310 25330 7362 25342
rect 7982 25394 8034 25406
rect 7982 25330 8034 25342
rect 2158 25282 2210 25294
rect 2158 25218 2210 25230
rect 2942 25282 2994 25294
rect 2942 25218 2994 25230
rect 4622 25282 4674 25294
rect 4622 25218 4674 25230
rect 9326 25282 9378 25294
rect 9326 25218 9378 25230
rect 11342 25282 11394 25294
rect 11342 25218 11394 25230
rect 13470 25282 13522 25294
rect 13470 25218 13522 25230
rect 15374 25282 15426 25294
rect 15374 25218 15426 25230
rect 17054 25282 17106 25294
rect 17054 25218 17106 25230
rect 19966 25282 20018 25294
rect 19966 25218 20018 25230
rect 21646 25282 21698 25294
rect 21646 25218 21698 25230
rect 22430 25282 22482 25294
rect 22430 25218 22482 25230
rect 23998 25282 24050 25294
rect 23998 25218 24050 25230
rect 24670 25282 24722 25294
rect 24670 25218 24722 25230
rect 25342 25282 25394 25294
rect 25342 25218 25394 25230
rect 26910 25282 26962 25294
rect 26910 25218 26962 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 1344 25114 28720 25148
rect 1344 25062 8018 25114
rect 8070 25062 8122 25114
rect 8174 25062 8226 25114
rect 8278 25062 14822 25114
rect 14874 25062 14926 25114
rect 14978 25062 15030 25114
rect 15082 25062 21626 25114
rect 21678 25062 21730 25114
rect 21782 25062 21834 25114
rect 21886 25062 28430 25114
rect 28482 25062 28534 25114
rect 28586 25062 28638 25114
rect 28690 25062 28720 25114
rect 1344 25028 28720 25062
rect 3278 24946 3330 24958
rect 3278 24882 3330 24894
rect 3502 24946 3554 24958
rect 3502 24882 3554 24894
rect 4286 24946 4338 24958
rect 4286 24882 4338 24894
rect 4734 24946 4786 24958
rect 4734 24882 4786 24894
rect 6078 24946 6130 24958
rect 6078 24882 6130 24894
rect 7422 24946 7474 24958
rect 7422 24882 7474 24894
rect 10446 24946 10498 24958
rect 10446 24882 10498 24894
rect 25454 24946 25506 24958
rect 25454 24882 25506 24894
rect 2046 24834 2098 24846
rect 2046 24770 2098 24782
rect 2382 24834 2434 24846
rect 2382 24770 2434 24782
rect 9662 24834 9714 24846
rect 9662 24770 9714 24782
rect 14366 24834 14418 24846
rect 14366 24770 14418 24782
rect 23326 24834 23378 24846
rect 23326 24770 23378 24782
rect 23998 24834 24050 24846
rect 23998 24770 24050 24782
rect 24334 24834 24386 24846
rect 24334 24770 24386 24782
rect 24670 24722 24722 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 3714 24670 3726 24722
rect 3778 24670 3790 24722
rect 14578 24670 14590 24722
rect 14642 24670 14654 24722
rect 23090 24670 23102 24722
rect 23154 24670 23166 24722
rect 23762 24670 23774 24722
rect 23826 24670 23838 24722
rect 24670 24658 24722 24670
rect 26574 24722 26626 24734
rect 26898 24670 26910 24722
rect 26962 24670 26974 24722
rect 26574 24658 26626 24670
rect 14142 24610 14194 24622
rect 14142 24546 14194 24558
rect 22766 24610 22818 24622
rect 26114 24558 26126 24610
rect 26178 24558 26190 24610
rect 28018 24558 28030 24610
rect 28082 24558 28094 24610
rect 22766 24546 22818 24558
rect 1344 24330 28560 24364
rect 1344 24278 4616 24330
rect 4668 24278 4720 24330
rect 4772 24278 4824 24330
rect 4876 24278 11420 24330
rect 11472 24278 11524 24330
rect 11576 24278 11628 24330
rect 11680 24278 18224 24330
rect 18276 24278 18328 24330
rect 18380 24278 18432 24330
rect 18484 24278 25028 24330
rect 25080 24278 25132 24330
rect 25184 24278 25236 24330
rect 25288 24278 28560 24330
rect 1344 24244 28560 24278
rect 27694 24162 27746 24174
rect 27694 24098 27746 24110
rect 23662 24050 23714 24062
rect 23662 23986 23714 23998
rect 9662 23938 9714 23950
rect 8418 23886 8430 23938
rect 8482 23886 8494 23938
rect 9202 23886 9214 23938
rect 9266 23886 9278 23938
rect 9662 23874 9714 23886
rect 10670 23938 10722 23950
rect 10670 23874 10722 23886
rect 11006 23938 11058 23950
rect 13806 23938 13858 23950
rect 15598 23938 15650 23950
rect 11890 23886 11902 23938
rect 11954 23886 11966 23938
rect 15026 23886 15038 23938
rect 15090 23886 15102 23938
rect 11006 23874 11058 23886
rect 13806 23874 13858 23886
rect 15598 23874 15650 23886
rect 16494 23938 16546 23950
rect 25230 23938 25282 23950
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 20514 23886 20526 23938
rect 20578 23886 20590 23938
rect 21410 23886 21422 23938
rect 21474 23886 21486 23938
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 16494 23874 16546 23886
rect 25230 23874 25282 23886
rect 25902 23938 25954 23950
rect 25902 23874 25954 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 2046 23762 2098 23774
rect 8654 23826 8706 23838
rect 8654 23762 8706 23774
rect 9998 23826 10050 23838
rect 9998 23762 10050 23774
rect 10334 23826 10386 23838
rect 10334 23762 10386 23774
rect 11342 23826 11394 23838
rect 11342 23762 11394 23774
rect 11678 23826 11730 23838
rect 11678 23762 11730 23774
rect 13470 23826 13522 23838
rect 13470 23762 13522 23774
rect 15262 23826 15314 23838
rect 15262 23762 15314 23774
rect 15934 23826 15986 23838
rect 15934 23762 15986 23774
rect 16830 23826 16882 23838
rect 16830 23762 16882 23774
rect 20078 23826 20130 23838
rect 20078 23762 20130 23774
rect 20750 23826 20802 23838
rect 20750 23762 20802 23774
rect 21646 23826 21698 23838
rect 21646 23762 21698 23774
rect 24222 23826 24274 23838
rect 24222 23762 24274 23774
rect 24558 23826 24610 23838
rect 24558 23762 24610 23774
rect 24894 23826 24946 23838
rect 24894 23762 24946 23774
rect 25566 23826 25618 23838
rect 25566 23762 25618 23774
rect 26238 23826 26290 23838
rect 26238 23762 26290 23774
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 8990 23714 9042 23726
rect 8990 23650 9042 23662
rect 26910 23714 26962 23726
rect 26910 23650 26962 23662
rect 1344 23546 28720 23580
rect 1344 23494 8018 23546
rect 8070 23494 8122 23546
rect 8174 23494 8226 23546
rect 8278 23494 14822 23546
rect 14874 23494 14926 23546
rect 14978 23494 15030 23546
rect 15082 23494 21626 23546
rect 21678 23494 21730 23546
rect 21782 23494 21834 23546
rect 21886 23494 28430 23546
rect 28482 23494 28534 23546
rect 28586 23494 28638 23546
rect 28690 23494 28720 23546
rect 1344 23460 28720 23494
rect 9550 23378 9602 23390
rect 9550 23314 9602 23326
rect 10558 23378 10610 23390
rect 10558 23314 10610 23326
rect 10894 23378 10946 23390
rect 10894 23314 10946 23326
rect 20862 23378 20914 23390
rect 20862 23314 20914 23326
rect 25566 23378 25618 23390
rect 25566 23314 25618 23326
rect 10222 23266 10274 23278
rect 10222 23202 10274 23214
rect 24670 23266 24722 23278
rect 24670 23202 24722 23214
rect 26238 23266 26290 23278
rect 26238 23202 26290 23214
rect 26910 23266 26962 23278
rect 26910 23202 26962 23214
rect 9762 23102 9774 23154
rect 9826 23102 9838 23154
rect 11106 23102 11118 23154
rect 11170 23102 11182 23154
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 24434 23102 24446 23154
rect 24498 23102 24510 23154
rect 25330 23102 25342 23154
rect 25394 23102 25406 23154
rect 26002 23102 26014 23154
rect 26066 23102 26078 23154
rect 28254 23042 28306 23054
rect 27458 22990 27470 23042
rect 27522 22990 27534 23042
rect 28254 22978 28306 22990
rect 1344 22762 28560 22796
rect 1344 22710 4616 22762
rect 4668 22710 4720 22762
rect 4772 22710 4824 22762
rect 4876 22710 11420 22762
rect 11472 22710 11524 22762
rect 11576 22710 11628 22762
rect 11680 22710 18224 22762
rect 18276 22710 18328 22762
rect 18380 22710 18432 22762
rect 18484 22710 25028 22762
rect 25080 22710 25132 22762
rect 25184 22710 25236 22762
rect 25288 22710 28560 22762
rect 1344 22676 28560 22710
rect 25666 22318 25678 22370
rect 25730 22318 25742 22370
rect 26898 22318 26910 22370
rect 26962 22318 26974 22370
rect 26238 22258 26290 22270
rect 26238 22194 26290 22206
rect 26574 22258 26626 22270
rect 28018 22206 28030 22258
rect 28082 22206 28094 22258
rect 26574 22194 26626 22206
rect 25902 22146 25954 22158
rect 25902 22082 25954 22094
rect 1344 21978 28720 22012
rect 1344 21926 8018 21978
rect 8070 21926 8122 21978
rect 8174 21926 8226 21978
rect 8278 21926 14822 21978
rect 14874 21926 14926 21978
rect 14978 21926 15030 21978
rect 15082 21926 21626 21978
rect 21678 21926 21730 21978
rect 21782 21926 21834 21978
rect 21886 21926 28430 21978
rect 28482 21926 28534 21978
rect 28586 21926 28638 21978
rect 28690 21926 28720 21978
rect 1344 21892 28720 21926
rect 26462 21810 26514 21822
rect 26462 21746 26514 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 26798 21698 26850 21710
rect 14802 21646 14814 21698
rect 14866 21646 14878 21698
rect 26798 21634 26850 21646
rect 27134 21698 27186 21710
rect 27134 21634 27186 21646
rect 27470 21586 27522 21598
rect 27470 21522 27522 21534
rect 28142 21586 28194 21598
rect 28142 21522 28194 21534
rect 26238 21474 26290 21486
rect 13794 21422 13806 21474
rect 13858 21422 13870 21474
rect 26238 21410 26290 21422
rect 1344 21194 28560 21228
rect 1344 21142 4616 21194
rect 4668 21142 4720 21194
rect 4772 21142 4824 21194
rect 4876 21142 11420 21194
rect 11472 21142 11524 21194
rect 11576 21142 11628 21194
rect 11680 21142 18224 21194
rect 18276 21142 18328 21194
rect 18380 21142 18432 21194
rect 18484 21142 25028 21194
rect 25080 21142 25132 21194
rect 25184 21142 25236 21194
rect 25288 21142 28560 21194
rect 1344 21108 28560 21142
rect 26686 20914 26738 20926
rect 16258 20862 16270 20914
rect 16322 20862 16334 20914
rect 24434 20862 24446 20914
rect 24498 20862 24510 20914
rect 26686 20850 26738 20862
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 17266 20638 17278 20690
rect 17330 20638 17342 20690
rect 25442 20638 25454 20690
rect 25506 20638 25518 20690
rect 28018 20638 28030 20690
rect 28082 20638 28094 20690
rect 23998 20578 24050 20590
rect 23998 20514 24050 20526
rect 1344 20410 28720 20444
rect 1344 20358 8018 20410
rect 8070 20358 8122 20410
rect 8174 20358 8226 20410
rect 8278 20358 14822 20410
rect 14874 20358 14926 20410
rect 14978 20358 15030 20410
rect 15082 20358 21626 20410
rect 21678 20358 21730 20410
rect 21782 20358 21834 20410
rect 21886 20358 28430 20410
rect 28482 20358 28534 20410
rect 28586 20358 28638 20410
rect 28690 20358 28720 20410
rect 1344 20324 28720 20358
rect 20514 20190 20526 20242
rect 20578 20190 20590 20242
rect 14590 20130 14642 20142
rect 14590 20066 14642 20078
rect 15374 20130 15426 20142
rect 27806 20130 27858 20142
rect 23538 20078 23550 20130
rect 23602 20078 23614 20130
rect 15374 20066 15426 20078
rect 27806 20066 27858 20078
rect 11902 20018 11954 20030
rect 17614 20018 17666 20030
rect 21086 20018 21138 20030
rect 28142 20018 28194 20030
rect 9874 19966 9886 20018
rect 9938 19966 9950 20018
rect 12338 19966 12350 20018
rect 12402 19966 12414 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 18050 19966 18062 20018
rect 18114 19966 18126 20018
rect 24434 19966 24446 20018
rect 24498 19966 24510 20018
rect 11902 19954 11954 19966
rect 17614 19954 17666 19966
rect 21086 19954 21138 19966
rect 28142 19954 28194 19966
rect 21534 19906 21586 19918
rect 21534 19842 21586 19854
rect 21870 19906 21922 19918
rect 25454 19906 25506 19918
rect 22306 19854 22318 19906
rect 22370 19854 22382 19906
rect 21870 19842 21922 19854
rect 25454 19842 25506 19854
rect 25902 19906 25954 19918
rect 25902 19842 25954 19854
rect 26238 19906 26290 19918
rect 26238 19842 26290 19854
rect 27582 19906 27634 19918
rect 27582 19842 27634 19854
rect 9538 19742 9550 19794
rect 9602 19742 9614 19794
rect 16370 19742 16382 19794
rect 16434 19742 16446 19794
rect 24098 19742 24110 19794
rect 24162 19742 24174 19794
rect 25442 19742 25454 19794
rect 25506 19791 25518 19794
rect 25890 19791 25902 19794
rect 25506 19745 25902 19791
rect 25506 19742 25518 19745
rect 25890 19742 25902 19745
rect 25954 19742 25966 19794
rect 1344 19626 28560 19660
rect 1344 19574 4616 19626
rect 4668 19574 4720 19626
rect 4772 19574 4824 19626
rect 4876 19574 11420 19626
rect 11472 19574 11524 19626
rect 11576 19574 11628 19626
rect 11680 19574 18224 19626
rect 18276 19574 18328 19626
rect 18380 19574 18432 19626
rect 18484 19574 25028 19626
rect 25080 19574 25132 19626
rect 25184 19574 25236 19626
rect 25288 19574 28560 19626
rect 1344 19540 28560 19574
rect 13022 19458 13074 19470
rect 14018 19406 14030 19458
rect 14082 19406 14094 19458
rect 21298 19406 21310 19458
rect 21362 19406 21374 19458
rect 13022 19394 13074 19406
rect 7634 19294 7646 19346
rect 7698 19294 7710 19346
rect 19170 19294 19182 19346
rect 19234 19294 19246 19346
rect 9550 19234 9602 19246
rect 14254 19234 14306 19246
rect 22430 19234 22482 19246
rect 9986 19182 9998 19234
rect 10050 19182 10062 19234
rect 13458 19182 13470 19234
rect 13522 19182 13534 19234
rect 14914 19182 14926 19234
rect 14978 19182 14990 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 26338 19182 26350 19234
rect 26402 19182 26414 19234
rect 9550 19170 9602 19182
rect 14254 19170 14306 19182
rect 22430 19170 22482 19182
rect 17166 19122 17218 19134
rect 8978 19070 8990 19122
rect 9042 19070 9054 19122
rect 17166 19058 17218 19070
rect 17950 19122 18002 19134
rect 27806 19122 27858 19134
rect 20178 19070 20190 19122
rect 20242 19070 20254 19122
rect 17950 19058 18002 19070
rect 27806 19058 27858 19070
rect 28142 19122 28194 19134
rect 28142 19058 28194 19070
rect 25902 19010 25954 19022
rect 27582 19010 27634 19022
rect 12226 18958 12238 19010
rect 12290 18958 12302 19010
rect 25106 18958 25118 19010
rect 25170 18958 25182 19010
rect 26114 18958 26126 19010
rect 26178 18958 26190 19010
rect 25902 18946 25954 18958
rect 27582 18946 27634 18958
rect 1344 18842 28720 18876
rect 1344 18790 8018 18842
rect 8070 18790 8122 18842
rect 8174 18790 8226 18842
rect 8278 18790 14822 18842
rect 14874 18790 14926 18842
rect 14978 18790 15030 18842
rect 15082 18790 21626 18842
rect 21678 18790 21730 18842
rect 21782 18790 21834 18842
rect 21886 18790 28430 18842
rect 28482 18790 28534 18842
rect 28586 18790 28638 18842
rect 28690 18790 28720 18842
rect 1344 18756 28720 18790
rect 8530 18622 8542 18674
rect 8594 18622 8606 18674
rect 23202 18622 23214 18674
rect 23266 18622 23278 18674
rect 24658 18622 24670 18674
rect 24722 18622 24734 18674
rect 16158 18562 16210 18574
rect 12562 18510 12574 18562
rect 12626 18510 12638 18562
rect 19394 18510 19406 18562
rect 19458 18510 19470 18562
rect 25890 18510 25902 18562
rect 25954 18510 25966 18562
rect 16158 18498 16210 18510
rect 13246 18450 13298 18462
rect 16942 18450 16994 18462
rect 23774 18450 23826 18462
rect 5506 18398 5518 18450
rect 5570 18398 5582 18450
rect 6066 18398 6078 18450
rect 6130 18398 6142 18450
rect 9874 18398 9886 18450
rect 9938 18398 9950 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 20178 18398 20190 18450
rect 20242 18398 20254 18450
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 24434 18398 24446 18450
rect 24498 18398 24510 18450
rect 13246 18386 13298 18398
rect 16942 18386 16994 18398
rect 23774 18386 23826 18398
rect 25342 18338 25394 18350
rect 27694 18338 27746 18350
rect 11554 18286 11566 18338
rect 11618 18286 11630 18338
rect 18386 18286 18398 18338
rect 18450 18286 18462 18338
rect 27122 18286 27134 18338
rect 27186 18286 27198 18338
rect 25342 18274 25394 18286
rect 27694 18274 27746 18286
rect 9102 18226 9154 18238
rect 10210 18174 10222 18226
rect 10274 18174 10286 18226
rect 9102 18162 9154 18174
rect 1344 18058 28560 18092
rect 1344 18006 4616 18058
rect 4668 18006 4720 18058
rect 4772 18006 4824 18058
rect 4876 18006 11420 18058
rect 11472 18006 11524 18058
rect 11576 18006 11628 18058
rect 11680 18006 18224 18058
rect 18276 18006 18328 18058
rect 18380 18006 18432 18058
rect 18484 18006 25028 18058
rect 25080 18006 25132 18058
rect 25184 18006 25236 18058
rect 25288 18006 28560 18058
rect 1344 17972 28560 18006
rect 11230 17890 11282 17902
rect 15822 17890 15874 17902
rect 12002 17838 12014 17890
rect 12066 17838 12078 17890
rect 11230 17826 11282 17838
rect 15822 17826 15874 17838
rect 21422 17778 21474 17790
rect 21422 17714 21474 17726
rect 23102 17778 23154 17790
rect 23102 17714 23154 17726
rect 7534 17666 7586 17678
rect 16158 17666 16210 17678
rect 27022 17666 27074 17678
rect 4498 17614 4510 17666
rect 4562 17614 4574 17666
rect 5618 17614 5630 17666
rect 5682 17614 5694 17666
rect 8194 17614 8206 17666
rect 8258 17614 8270 17666
rect 11666 17614 11678 17666
rect 11730 17614 11742 17666
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 15698 17614 15710 17666
rect 15762 17614 15774 17666
rect 16818 17614 16830 17666
rect 16882 17614 16894 17666
rect 20626 17614 20638 17666
rect 20690 17614 20702 17666
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 26338 17614 26350 17666
rect 26402 17614 26414 17666
rect 7534 17602 7586 17614
rect 16158 17602 16210 17614
rect 27022 17602 27074 17614
rect 28142 17666 28194 17678
rect 28142 17602 28194 17614
rect 10446 17554 10498 17566
rect 10446 17490 10498 17502
rect 27806 17554 27858 17566
rect 27806 17490 27858 17502
rect 4958 17442 5010 17454
rect 6638 17442 6690 17454
rect 3938 17390 3950 17442
rect 4002 17390 4014 17442
rect 6178 17390 6190 17442
rect 6242 17390 6254 17442
rect 4958 17378 5010 17390
rect 6638 17378 6690 17390
rect 13806 17442 13858 17454
rect 19854 17442 19906 17454
rect 22542 17442 22594 17454
rect 19282 17390 19294 17442
rect 19346 17390 19358 17442
rect 20066 17390 20078 17442
rect 20130 17390 20142 17442
rect 13806 17378 13858 17390
rect 19854 17378 19906 17390
rect 22542 17378 22594 17390
rect 23326 17442 23378 17454
rect 27358 17442 27410 17454
rect 23874 17390 23886 17442
rect 23938 17390 23950 17442
rect 23326 17378 23378 17390
rect 27358 17378 27410 17390
rect 1344 17274 28720 17308
rect 1344 17222 8018 17274
rect 8070 17222 8122 17274
rect 8174 17222 8226 17274
rect 8278 17222 14822 17274
rect 14874 17222 14926 17274
rect 14978 17222 15030 17274
rect 15082 17222 21626 17274
rect 21678 17222 21730 17274
rect 21782 17222 21834 17274
rect 21886 17222 28430 17274
rect 28482 17222 28534 17274
rect 28586 17222 28638 17274
rect 28690 17222 28720 17274
rect 1344 17188 28720 17222
rect 9102 17106 9154 17118
rect 2258 17054 2270 17106
rect 2322 17054 2334 17106
rect 9102 17042 9154 17054
rect 21646 17106 21698 17118
rect 21646 17042 21698 17054
rect 8318 16994 8370 17006
rect 20862 16994 20914 17006
rect 9762 16942 9774 16994
rect 9826 16942 9838 16994
rect 23986 16942 23998 16994
rect 24050 16942 24062 16994
rect 27682 16942 27694 16994
rect 27746 16942 27758 16994
rect 8318 16930 8370 16942
rect 20862 16930 20914 16942
rect 5070 16882 5122 16894
rect 17950 16882 18002 16894
rect 21982 16882 22034 16894
rect 4610 16830 4622 16882
rect 4674 16830 4686 16882
rect 5506 16830 5518 16882
rect 5570 16830 5582 16882
rect 6066 16830 6078 16882
rect 6130 16830 6142 16882
rect 14578 16830 14590 16882
rect 14642 16830 14654 16882
rect 18610 16830 18622 16882
rect 18674 16830 18686 16882
rect 5070 16818 5122 16830
rect 17950 16818 18002 16830
rect 21982 16818 22034 16830
rect 22430 16882 22482 16894
rect 22430 16818 22482 16830
rect 22866 16718 22878 16770
rect 22930 16718 22942 16770
rect 26674 16718 26686 16770
rect 26738 16718 26750 16770
rect 1598 16658 1650 16670
rect 1598 16594 1650 16606
rect 1344 16490 28560 16524
rect 1344 16438 4616 16490
rect 4668 16438 4720 16490
rect 4772 16438 4824 16490
rect 4876 16438 11420 16490
rect 11472 16438 11524 16490
rect 11576 16438 11628 16490
rect 11680 16438 18224 16490
rect 18276 16438 18328 16490
rect 18380 16438 18432 16490
rect 18484 16438 25028 16490
rect 25080 16438 25132 16490
rect 25184 16438 25236 16490
rect 25288 16438 28560 16490
rect 1344 16404 28560 16438
rect 3938 16158 3950 16210
rect 4002 16158 4014 16210
rect 6962 16158 6974 16210
rect 7026 16158 7038 16210
rect 9762 16158 9774 16210
rect 9826 16158 9838 16210
rect 14690 16158 14702 16210
rect 14754 16158 14766 16210
rect 19282 16158 19294 16210
rect 19346 16158 19358 16210
rect 21970 16046 21982 16098
rect 22034 16046 22046 16098
rect 2706 15934 2718 15986
rect 2770 15934 2782 15986
rect 7970 15934 7982 15986
rect 8034 15934 8046 15986
rect 10770 15934 10782 15986
rect 10834 15934 10846 15986
rect 13570 15934 13582 15986
rect 13634 15934 13646 15986
rect 20290 15934 20302 15986
rect 20354 15934 20366 15986
rect 25778 15934 25790 15986
rect 25842 15934 25854 15986
rect 1344 15706 28720 15740
rect 1344 15654 8018 15706
rect 8070 15654 8122 15706
rect 8174 15654 8226 15706
rect 8278 15654 14822 15706
rect 14874 15654 14926 15706
rect 14978 15654 15030 15706
rect 15082 15654 21626 15706
rect 21678 15654 21730 15706
rect 21782 15654 21834 15706
rect 21886 15654 28430 15706
rect 28482 15654 28534 15706
rect 28586 15654 28638 15706
rect 28690 15654 28720 15706
rect 1344 15620 28720 15654
rect 7086 15538 7138 15550
rect 12014 15538 12066 15550
rect 6290 15486 6302 15538
rect 6354 15486 6366 15538
rect 8418 15486 8430 15538
rect 8482 15486 8494 15538
rect 12786 15486 12798 15538
rect 12850 15486 12862 15538
rect 22754 15486 22766 15538
rect 22818 15486 22830 15538
rect 7086 15474 7138 15486
rect 12014 15474 12066 15486
rect 27234 15374 27246 15426
rect 27298 15374 27310 15426
rect 3614 15314 3666 15326
rect 15710 15314 15762 15326
rect 2706 15262 2718 15314
rect 2770 15262 2782 15314
rect 3938 15262 3950 15314
rect 4002 15262 4014 15314
rect 8978 15262 8990 15314
rect 9042 15262 9054 15314
rect 11442 15262 11454 15314
rect 11506 15262 11518 15314
rect 15026 15262 15038 15314
rect 15090 15262 15102 15314
rect 3614 15250 3666 15262
rect 15710 15250 15762 15262
rect 16046 15314 16098 15326
rect 16046 15250 16098 15262
rect 20078 15314 20130 15326
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 24546 15262 24558 15314
rect 24610 15262 24622 15314
rect 20078 15250 20130 15262
rect 2046 15202 2098 15214
rect 25342 15202 25394 15214
rect 2594 15150 2606 15202
rect 2658 15150 2670 15202
rect 2046 15138 2098 15150
rect 25342 15138 25394 15150
rect 25790 15202 25842 15214
rect 26226 15150 26238 15202
rect 26290 15150 26302 15202
rect 25790 15138 25842 15150
rect 23550 15090 23602 15102
rect 11218 15038 11230 15090
rect 11282 15038 11294 15090
rect 23550 15026 23602 15038
rect 24446 15090 24498 15102
rect 24446 15026 24498 15038
rect 1344 14922 28560 14956
rect 1344 14870 4616 14922
rect 4668 14870 4720 14922
rect 4772 14870 4824 14922
rect 4876 14870 11420 14922
rect 11472 14870 11524 14922
rect 11576 14870 11628 14922
rect 11680 14870 18224 14922
rect 18276 14870 18328 14922
rect 18380 14870 18432 14922
rect 18484 14870 25028 14922
rect 25080 14870 25132 14922
rect 25184 14870 25236 14922
rect 25288 14870 28560 14922
rect 1344 14836 28560 14870
rect 25566 14754 25618 14766
rect 2258 14702 2270 14754
rect 2322 14702 2334 14754
rect 20738 14702 20750 14754
rect 20802 14702 20814 14754
rect 25566 14690 25618 14702
rect 4050 14590 4062 14642
rect 4114 14590 4126 14642
rect 14466 14590 14478 14642
rect 14530 14590 14542 14642
rect 25890 14590 25902 14642
rect 25954 14590 25966 14642
rect 9214 14530 9266 14542
rect 2034 14478 2046 14530
rect 2098 14478 2110 14530
rect 8642 14478 8654 14530
rect 8706 14478 8718 14530
rect 9214 14466 9266 14478
rect 9550 14530 9602 14542
rect 22094 14530 22146 14542
rect 28142 14530 28194 14542
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 20514 14478 20526 14530
rect 20578 14478 20590 14530
rect 22530 14478 22542 14530
rect 22594 14478 22606 14530
rect 26338 14478 26350 14530
rect 26402 14478 26414 14530
rect 27122 14478 27134 14530
rect 27186 14478 27198 14530
rect 9550 14466 9602 14478
rect 22094 14466 22146 14478
rect 28142 14466 28194 14478
rect 5518 14418 5570 14430
rect 3042 14366 3054 14418
rect 3106 14366 3118 14418
rect 5518 14354 5570 14366
rect 13022 14418 13074 14430
rect 24782 14418 24834 14430
rect 15474 14366 15486 14418
rect 15538 14366 15550 14418
rect 13022 14354 13074 14366
rect 24782 14354 24834 14366
rect 4510 14306 4562 14318
rect 19854 14306 19906 14318
rect 27694 14306 27746 14318
rect 6066 14254 6078 14306
rect 6130 14254 6142 14306
rect 12450 14254 12462 14306
rect 12514 14254 12526 14306
rect 26674 14254 26686 14306
rect 26738 14254 26750 14306
rect 4510 14242 4562 14254
rect 19854 14242 19906 14254
rect 27694 14242 27746 14254
rect 1344 14138 28720 14172
rect 1344 14086 8018 14138
rect 8070 14086 8122 14138
rect 8174 14086 8226 14138
rect 8278 14086 14822 14138
rect 14874 14086 14926 14138
rect 14978 14086 15030 14138
rect 15082 14086 21626 14138
rect 21678 14086 21730 14138
rect 21782 14086 21834 14138
rect 21886 14086 28430 14138
rect 28482 14086 28534 14138
rect 28586 14086 28638 14138
rect 28690 14086 28720 14138
rect 1344 14052 28720 14086
rect 25454 13970 25506 13982
rect 2594 13918 2606 13970
rect 2658 13918 2670 13970
rect 24210 13918 24222 13970
rect 24274 13918 24286 13970
rect 25454 13906 25506 13918
rect 6962 13806 6974 13858
rect 7026 13806 7038 13858
rect 18834 13806 18846 13858
rect 18898 13806 18910 13858
rect 27234 13806 27246 13858
rect 27298 13806 27310 13858
rect 5742 13746 5794 13758
rect 10894 13746 10946 13758
rect 21310 13746 21362 13758
rect 5058 13694 5070 13746
rect 5122 13694 5134 13746
rect 10098 13694 10110 13746
rect 10162 13694 10174 13746
rect 14466 13694 14478 13746
rect 14530 13694 14542 13746
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 5742 13682 5794 13694
rect 10894 13682 10946 13694
rect 21310 13682 21362 13694
rect 26014 13634 26066 13646
rect 7970 13582 7982 13634
rect 8034 13582 8046 13634
rect 19842 13582 19854 13634
rect 19906 13582 19918 13634
rect 26226 13582 26238 13634
rect 26290 13582 26302 13634
rect 26014 13570 26066 13582
rect 2046 13522 2098 13534
rect 13918 13522 13970 13534
rect 10434 13470 10446 13522
rect 10498 13470 10510 13522
rect 2046 13458 2098 13470
rect 13918 13458 13970 13470
rect 24782 13522 24834 13534
rect 24782 13458 24834 13470
rect 1344 13354 28560 13388
rect 1344 13302 4616 13354
rect 4668 13302 4720 13354
rect 4772 13302 4824 13354
rect 4876 13302 11420 13354
rect 11472 13302 11524 13354
rect 11576 13302 11628 13354
rect 11680 13302 18224 13354
rect 18276 13302 18328 13354
rect 18380 13302 18432 13354
rect 18484 13302 25028 13354
rect 25080 13302 25132 13354
rect 25184 13302 25236 13354
rect 25288 13302 28560 13354
rect 1344 13268 28560 13302
rect 9102 13186 9154 13198
rect 13458 13134 13470 13186
rect 13522 13134 13534 13186
rect 9102 13122 9154 13134
rect 27134 13074 27186 13086
rect 4050 13022 4062 13074
rect 4114 13022 4126 13074
rect 7858 13022 7870 13074
rect 7922 13022 7934 13074
rect 16818 13022 16830 13074
rect 16882 13022 16894 13074
rect 27134 13010 27186 13022
rect 12574 12962 12626 12974
rect 23214 12962 23266 12974
rect 12226 12910 12238 12962
rect 12290 12910 12302 12962
rect 13906 12910 13918 12962
rect 13970 12910 13982 12962
rect 15138 12910 15150 12962
rect 15202 12910 15214 12962
rect 23650 12910 23662 12962
rect 23714 12910 23726 12962
rect 12574 12898 12626 12910
rect 23214 12898 23266 12910
rect 9886 12850 9938 12862
rect 2706 12798 2718 12850
rect 2770 12798 2782 12850
rect 6514 12798 6526 12850
rect 6578 12798 6590 12850
rect 9886 12786 9938 12798
rect 25902 12850 25954 12862
rect 25902 12786 25954 12798
rect 26686 12738 26738 12750
rect 26686 12674 26738 12686
rect 1344 12570 28720 12604
rect 1344 12518 8018 12570
rect 8070 12518 8122 12570
rect 8174 12518 8226 12570
rect 8278 12518 14822 12570
rect 14874 12518 14926 12570
rect 14978 12518 15030 12570
rect 15082 12518 21626 12570
rect 21678 12518 21730 12570
rect 21782 12518 21834 12570
rect 21886 12518 28430 12570
rect 28482 12518 28534 12570
rect 28586 12518 28638 12570
rect 28690 12518 28720 12570
rect 1344 12484 28720 12518
rect 5406 12402 5458 12414
rect 5406 12338 5458 12350
rect 15262 12402 15314 12414
rect 15262 12338 15314 12350
rect 19742 12402 19794 12414
rect 19742 12338 19794 12350
rect 2382 12290 2434 12302
rect 2382 12226 2434 12238
rect 6190 12290 6242 12302
rect 6190 12226 6242 12238
rect 20526 12290 20578 12302
rect 27346 12238 27358 12290
rect 27410 12238 27422 12290
rect 20526 12226 20578 12238
rect 5294 12178 5346 12190
rect 9102 12178 9154 12190
rect 23438 12178 23490 12190
rect 4610 12126 4622 12178
rect 4674 12126 4686 12178
rect 8418 12126 8430 12178
rect 8482 12126 8494 12178
rect 14578 12126 14590 12178
rect 14642 12126 14654 12178
rect 22866 12126 22878 12178
rect 22930 12126 22942 12178
rect 24546 12126 24558 12178
rect 24610 12126 24622 12178
rect 5294 12114 5346 12126
rect 9102 12114 9154 12126
rect 23438 12114 23490 12126
rect 25342 12066 25394 12078
rect 10770 12014 10782 12066
rect 10834 12014 10846 12066
rect 26450 12014 26462 12066
rect 26514 12014 26526 12066
rect 25342 12002 25394 12014
rect 1598 11954 1650 11966
rect 24098 11902 24110 11954
rect 24162 11902 24174 11954
rect 1598 11890 1650 11902
rect 1344 11786 28560 11820
rect 1344 11734 4616 11786
rect 4668 11734 4720 11786
rect 4772 11734 4824 11786
rect 4876 11734 11420 11786
rect 11472 11734 11524 11786
rect 11576 11734 11628 11786
rect 11680 11734 18224 11786
rect 18276 11734 18328 11786
rect 18380 11734 18432 11786
rect 18484 11734 25028 11786
rect 25080 11734 25132 11786
rect 25184 11734 25236 11786
rect 25288 11734 28560 11786
rect 1344 11700 28560 11734
rect 3826 11454 3838 11506
rect 3890 11454 3902 11506
rect 18050 11454 18062 11506
rect 18114 11454 18126 11506
rect 7310 11394 7362 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 6290 11342 6302 11394
rect 6354 11342 6366 11394
rect 7310 11330 7362 11342
rect 7758 11394 7810 11406
rect 14142 11394 14194 11406
rect 8082 11342 8094 11394
rect 8146 11342 8158 11394
rect 14466 11342 14478 11394
rect 14530 11342 14542 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 21970 11342 21982 11394
rect 22034 11342 22046 11394
rect 27346 11342 27358 11394
rect 27410 11342 27422 11394
rect 7758 11330 7810 11342
rect 14142 11330 14194 11342
rect 10446 11282 10498 11294
rect 2706 11230 2718 11282
rect 2770 11230 2782 11282
rect 13794 11230 13806 11282
rect 13858 11230 13870 11282
rect 24322 11230 24334 11282
rect 24386 11230 24398 11282
rect 10446 11218 10498 11230
rect 2046 11170 2098 11182
rect 11230 11170 11282 11182
rect 6850 11118 6862 11170
rect 6914 11118 6926 11170
rect 20738 11118 20750 11170
rect 20802 11118 20814 11170
rect 26898 11118 26910 11170
rect 26962 11118 26974 11170
rect 2046 11106 2098 11118
rect 11230 11106 11282 11118
rect 1344 11002 28720 11036
rect 1344 10950 8018 11002
rect 8070 10950 8122 11002
rect 8174 10950 8226 11002
rect 8278 10950 14822 11002
rect 14874 10950 14926 11002
rect 14978 10950 15030 11002
rect 15082 10950 21626 11002
rect 21678 10950 21730 11002
rect 21782 10950 21834 11002
rect 21886 10950 28430 11002
rect 28482 10950 28534 11002
rect 28586 10950 28638 11002
rect 28690 10950 28720 11002
rect 1344 10916 28720 10950
rect 1822 10834 1874 10846
rect 23774 10834 23826 10846
rect 6962 10782 6974 10834
rect 7026 10782 7038 10834
rect 8082 10782 8094 10834
rect 8146 10782 8158 10834
rect 22306 10782 22318 10834
rect 22370 10782 22382 10834
rect 1822 10770 1874 10782
rect 23774 10770 23826 10782
rect 23102 10722 23154 10734
rect 15810 10670 15822 10722
rect 15874 10670 15886 10722
rect 27234 10670 27246 10722
rect 27298 10670 27310 10722
rect 23102 10658 23154 10670
rect 2942 10610 2994 10622
rect 4286 10610 4338 10622
rect 19630 10610 19682 10622
rect 3266 10558 3278 10610
rect 3330 10558 3342 10610
rect 4722 10558 4734 10610
rect 4786 10558 4798 10610
rect 8530 10558 8542 10610
rect 8594 10558 8606 10610
rect 13458 10558 13470 10610
rect 13522 10558 13534 10610
rect 18274 10558 18286 10610
rect 18338 10558 18350 10610
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 23874 10558 23886 10610
rect 23938 10558 23950 10610
rect 2942 10546 2994 10558
rect 4286 10546 4338 10558
rect 19630 10546 19682 10558
rect 24334 10498 24386 10510
rect 3714 10446 3726 10498
rect 3778 10446 3790 10498
rect 9874 10446 9886 10498
rect 9938 10446 9950 10498
rect 14802 10446 14814 10498
rect 14866 10446 14878 10498
rect 26226 10446 26238 10498
rect 26290 10446 26302 10498
rect 24334 10434 24386 10446
rect 7758 10386 7810 10398
rect 18050 10334 18062 10386
rect 18114 10334 18126 10386
rect 7758 10322 7810 10334
rect 1344 10218 28560 10252
rect 1344 10166 4616 10218
rect 4668 10166 4720 10218
rect 4772 10166 4824 10218
rect 4876 10166 11420 10218
rect 11472 10166 11524 10218
rect 11576 10166 11628 10218
rect 11680 10166 18224 10218
rect 18276 10166 18328 10218
rect 18380 10166 18432 10218
rect 18484 10166 25028 10218
rect 25080 10166 25132 10218
rect 25184 10166 25236 10218
rect 25288 10166 28560 10218
rect 1344 10132 28560 10166
rect 12686 10050 12738 10062
rect 12686 9986 12738 9998
rect 17502 10050 17554 10062
rect 17502 9986 17554 9998
rect 6638 9938 6690 9950
rect 8990 9938 9042 9950
rect 3826 9886 3838 9938
rect 3890 9886 3902 9938
rect 8418 9886 8430 9938
rect 8482 9886 8494 9938
rect 19058 9886 19070 9938
rect 19122 9886 19134 9938
rect 27458 9886 27470 9938
rect 27522 9886 27534 9938
rect 6638 9874 6690 9886
rect 8990 9874 9042 9886
rect 21534 9826 21586 9838
rect 6178 9774 6190 9826
rect 6242 9774 6254 9826
rect 10322 9774 10334 9826
rect 10386 9774 10398 9826
rect 14130 9774 14142 9826
rect 14194 9774 14206 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 21534 9762 21586 9774
rect 4946 9662 4958 9714
rect 5010 9662 5022 9714
rect 7522 9662 7534 9714
rect 7586 9662 7598 9714
rect 20402 9662 20414 9714
rect 20466 9662 20478 9714
rect 26338 9662 26350 9714
rect 26402 9662 26414 9714
rect 25006 9602 25058 9614
rect 5618 9550 5630 9602
rect 5682 9550 5694 9602
rect 24434 9550 24446 9602
rect 24498 9550 24510 9602
rect 25006 9538 25058 9550
rect 25342 9602 25394 9614
rect 25342 9538 25394 9550
rect 1344 9434 28720 9468
rect 1344 9382 8018 9434
rect 8070 9382 8122 9434
rect 8174 9382 8226 9434
rect 8278 9382 14822 9434
rect 14874 9382 14926 9434
rect 14978 9382 15030 9434
rect 15082 9382 21626 9434
rect 21678 9382 21730 9434
rect 21782 9382 21834 9434
rect 21886 9382 28430 9434
rect 28482 9382 28534 9434
rect 28586 9382 28638 9434
rect 28690 9382 28720 9434
rect 1344 9348 28720 9382
rect 16270 9266 16322 9278
rect 5618 9214 5630 9266
rect 5682 9214 5694 9266
rect 15362 9214 15374 9266
rect 15426 9214 15438 9266
rect 16270 9202 16322 9214
rect 20190 9154 20242 9166
rect 20190 9090 20242 9102
rect 21870 9154 21922 9166
rect 27234 9102 27246 9154
rect 27298 9102 27310 9154
rect 21870 9090 21922 9102
rect 2718 9042 2770 9054
rect 12238 9042 12290 9054
rect 15934 9042 15986 9054
rect 3378 8990 3390 9042
rect 3442 8990 3454 9042
rect 12898 8990 12910 9042
rect 12962 8990 12974 9042
rect 2718 8978 2770 8990
rect 12238 8978 12290 8990
rect 15934 8978 15986 8990
rect 17278 9042 17330 9054
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 24658 8990 24670 9042
rect 24722 8990 24734 9042
rect 17278 8978 17330 8990
rect 16158 8930 16210 8942
rect 16158 8866 16210 8878
rect 25342 8930 25394 8942
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 25342 8866 25394 8878
rect 6414 8818 6466 8830
rect 6414 8754 6466 8766
rect 20974 8818 21026 8830
rect 20974 8754 21026 8766
rect 21086 8818 21138 8830
rect 21086 8754 21138 8766
rect 1344 8650 28560 8684
rect 1344 8598 4616 8650
rect 4668 8598 4720 8650
rect 4772 8598 4824 8650
rect 4876 8598 11420 8650
rect 11472 8598 11524 8650
rect 11576 8598 11628 8650
rect 11680 8598 18224 8650
rect 18276 8598 18328 8650
rect 18380 8598 18432 8650
rect 18484 8598 25028 8650
rect 25080 8598 25132 8650
rect 25184 8598 25236 8650
rect 25288 8598 28560 8650
rect 1344 8564 28560 8598
rect 4498 8430 4510 8482
rect 4562 8430 4574 8482
rect 22754 8430 22766 8482
rect 22818 8430 22830 8482
rect 5854 8370 5906 8382
rect 23550 8370 23602 8382
rect 6738 8318 6750 8370
rect 6802 8318 6814 8370
rect 19282 8318 19294 8370
rect 19346 8318 19358 8370
rect 5854 8306 5906 8318
rect 23550 8306 23602 8318
rect 14926 8258 14978 8270
rect 4834 8206 4846 8258
rect 4898 8206 4910 8258
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 19058 8206 19070 8258
rect 19122 8206 19134 8258
rect 21410 8206 21422 8258
rect 21474 8206 21486 8258
rect 22978 8206 22990 8258
rect 23042 8206 23054 8258
rect 26674 8206 26686 8258
rect 26738 8206 26750 8258
rect 27122 8206 27134 8258
rect 27186 8206 27198 8258
rect 27458 8206 27470 8258
rect 27522 8206 27534 8258
rect 14926 8194 14978 8206
rect 7746 8094 7758 8146
rect 7810 8094 7822 8146
rect 18398 8034 18450 8046
rect 17826 7982 17838 8034
rect 17890 7982 17902 8034
rect 18398 7970 18450 7982
rect 20750 8034 20802 8046
rect 27582 8034 27634 8046
rect 21970 7982 21982 8034
rect 22034 7982 22046 8034
rect 24210 7982 24222 8034
rect 24274 7982 24286 8034
rect 20750 7970 20802 7982
rect 27582 7970 27634 7982
rect 1344 7866 28720 7900
rect 1344 7814 8018 7866
rect 8070 7814 8122 7866
rect 8174 7814 8226 7866
rect 8278 7814 14822 7866
rect 14874 7814 14926 7866
rect 14978 7814 15030 7866
rect 15082 7814 21626 7866
rect 21678 7814 21730 7866
rect 21782 7814 21834 7866
rect 21886 7814 28430 7866
rect 28482 7814 28534 7866
rect 28586 7814 28638 7866
rect 28690 7814 28720 7866
rect 1344 7780 28720 7814
rect 5518 7698 5570 7710
rect 18510 7698 18562 7710
rect 4722 7646 4734 7698
rect 4786 7646 4798 7698
rect 13682 7646 13694 7698
rect 13746 7646 13758 7698
rect 22194 7646 22206 7698
rect 22258 7646 22270 7698
rect 5518 7634 5570 7646
rect 18510 7634 18562 7646
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 2046 7474 2098 7486
rect 10782 7474 10834 7486
rect 19294 7474 19346 7486
rect 2370 7422 2382 7474
rect 2434 7422 2446 7474
rect 11218 7422 11230 7474
rect 11282 7422 11294 7474
rect 19954 7422 19966 7474
rect 20018 7422 20030 7474
rect 24322 7422 24334 7474
rect 24386 7422 24398 7474
rect 2046 7410 2098 7422
rect 10782 7410 10834 7422
rect 19294 7410 19346 7422
rect 23326 7362 23378 7374
rect 28142 7362 28194 7374
rect 26226 7310 26238 7362
rect 26290 7310 26302 7362
rect 23326 7298 23378 7310
rect 28142 7298 28194 7310
rect 14254 7250 14306 7262
rect 14254 7186 14306 7198
rect 22990 7250 23042 7262
rect 22990 7186 23042 7198
rect 24558 7250 24610 7262
rect 24558 7186 24610 7198
rect 1344 7082 28560 7116
rect 1344 7030 4616 7082
rect 4668 7030 4720 7082
rect 4772 7030 4824 7082
rect 4876 7030 11420 7082
rect 11472 7030 11524 7082
rect 11576 7030 11628 7082
rect 11680 7030 18224 7082
rect 18276 7030 18328 7082
rect 18380 7030 18432 7082
rect 18484 7030 25028 7082
rect 25080 7030 25132 7082
rect 25184 7030 25236 7082
rect 25288 7030 28560 7082
rect 1344 6996 28560 7030
rect 14466 6750 14478 6802
rect 14530 6750 14542 6802
rect 17266 6750 17278 6802
rect 17330 6750 17342 6802
rect 22654 6690 22706 6702
rect 27694 6690 27746 6702
rect 23314 6638 23326 6690
rect 23378 6638 23390 6690
rect 22654 6626 22706 6638
rect 27694 6626 27746 6638
rect 15474 6526 15486 6578
rect 15538 6526 15550 6578
rect 18610 6526 18622 6578
rect 18674 6526 18686 6578
rect 1710 6466 1762 6478
rect 26350 6466 26402 6478
rect 25778 6414 25790 6466
rect 25842 6414 25854 6466
rect 1710 6402 1762 6414
rect 26350 6402 26402 6414
rect 26910 6466 26962 6478
rect 26910 6402 26962 6414
rect 28142 6466 28194 6478
rect 28142 6402 28194 6414
rect 1344 6298 28720 6332
rect 1344 6246 8018 6298
rect 8070 6246 8122 6298
rect 8174 6246 8226 6298
rect 8278 6246 14822 6298
rect 14874 6246 14926 6298
rect 14978 6246 15030 6298
rect 15082 6246 21626 6298
rect 21678 6246 21730 6298
rect 21782 6246 21834 6298
rect 21886 6246 28430 6298
rect 28482 6246 28534 6298
rect 28586 6246 28638 6298
rect 28690 6246 28720 6298
rect 1344 6212 28720 6246
rect 24670 6018 24722 6030
rect 20290 5966 20302 6018
rect 20354 5966 20366 6018
rect 23090 5966 23102 6018
rect 23154 5966 23166 6018
rect 27234 5966 27246 6018
rect 27298 5966 27310 6018
rect 24670 5954 24722 5966
rect 24334 5906 24386 5918
rect 24334 5842 24386 5854
rect 19506 5742 19518 5794
rect 19570 5742 19582 5794
rect 22082 5742 22094 5794
rect 22146 5742 22158 5794
rect 26226 5742 26238 5794
rect 26290 5742 26302 5794
rect 1344 5514 28560 5548
rect 1344 5462 4616 5514
rect 4668 5462 4720 5514
rect 4772 5462 4824 5514
rect 4876 5462 11420 5514
rect 11472 5462 11524 5514
rect 11576 5462 11628 5514
rect 11680 5462 18224 5514
rect 18276 5462 18328 5514
rect 18380 5462 18432 5514
rect 18484 5462 25028 5514
rect 25080 5462 25132 5514
rect 25184 5462 25236 5514
rect 25288 5462 28560 5514
rect 1344 5428 28560 5462
rect 26126 5346 26178 5358
rect 26126 5282 26178 5294
rect 27694 5346 27746 5358
rect 27694 5282 27746 5294
rect 28142 5234 28194 5246
rect 28142 5170 28194 5182
rect 21870 5122 21922 5134
rect 9986 5070 9998 5122
rect 10050 5070 10062 5122
rect 12002 5070 12014 5122
rect 12066 5070 12078 5122
rect 12674 5070 12686 5122
rect 12738 5070 12750 5122
rect 18274 5070 18286 5122
rect 18338 5070 18350 5122
rect 21870 5058 21922 5070
rect 22654 5122 22706 5134
rect 26910 5122 26962 5134
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 22654 5058 22706 5070
rect 26910 5058 26962 5070
rect 10558 5010 10610 5022
rect 10558 4946 10610 4958
rect 10894 5010 10946 5022
rect 10894 4946 10946 4958
rect 11230 5010 11282 5022
rect 11230 4946 11282 4958
rect 13470 5010 13522 5022
rect 13470 4946 13522 4958
rect 14478 5010 14530 5022
rect 14478 4946 14530 4958
rect 25342 5010 25394 5022
rect 25342 4946 25394 4958
rect 10222 4898 10274 4910
rect 10222 4834 10274 4846
rect 11566 4898 11618 4910
rect 11566 4834 11618 4846
rect 12238 4898 12290 4910
rect 12238 4834 12290 4846
rect 12910 4898 12962 4910
rect 12910 4834 12962 4846
rect 13806 4898 13858 4910
rect 13806 4834 13858 4846
rect 14814 4898 14866 4910
rect 14814 4834 14866 4846
rect 17838 4898 17890 4910
rect 17838 4834 17890 4846
rect 18510 4898 18562 4910
rect 18510 4834 18562 4846
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 22206 4898 22258 4910
rect 22206 4834 22258 4846
rect 26574 4898 26626 4910
rect 26574 4834 26626 4846
rect 1344 4730 28720 4764
rect 1344 4678 8018 4730
rect 8070 4678 8122 4730
rect 8174 4678 8226 4730
rect 8278 4678 14822 4730
rect 14874 4678 14926 4730
rect 14978 4678 15030 4730
rect 15082 4678 21626 4730
rect 21678 4678 21730 4730
rect 21782 4678 21834 4730
rect 21886 4678 28430 4730
rect 28482 4678 28534 4730
rect 28586 4678 28638 4730
rect 28690 4678 28720 4730
rect 1344 4644 28720 4678
rect 10334 4562 10386 4574
rect 10334 4498 10386 4510
rect 12126 4562 12178 4574
rect 12126 4498 12178 4510
rect 13694 4562 13746 4574
rect 13694 4498 13746 4510
rect 15262 4562 15314 4574
rect 15262 4498 15314 4510
rect 18062 4562 18114 4574
rect 18062 4498 18114 4510
rect 18734 4562 18786 4574
rect 18734 4498 18786 4510
rect 24222 4562 24274 4574
rect 24222 4498 24274 4510
rect 24782 4562 24834 4574
rect 24782 4498 24834 4510
rect 8654 4450 8706 4462
rect 8654 4386 8706 4398
rect 9662 4450 9714 4462
rect 17390 4450 17442 4462
rect 9986 4398 9998 4450
rect 10050 4398 10062 4450
rect 9662 4386 9714 4398
rect 17390 4386 17442 4398
rect 20414 4450 20466 4462
rect 20414 4386 20466 4398
rect 20750 4450 20802 4462
rect 20750 4386 20802 4398
rect 21086 4450 21138 4462
rect 21086 4386 21138 4398
rect 21758 4450 21810 4462
rect 21758 4386 21810 4398
rect 22430 4450 22482 4462
rect 22430 4386 22482 4398
rect 22766 4450 22818 4462
rect 22766 4386 22818 4398
rect 23102 4450 23154 4462
rect 23102 4386 23154 4398
rect 23438 4450 23490 4462
rect 27458 4398 27470 4450
rect 27522 4398 27534 4450
rect 23438 4386 23490 4398
rect 14926 4338 14978 4350
rect 10546 4286 10558 4338
rect 10610 4286 10622 4338
rect 14926 4274 14978 4286
rect 15598 4338 15650 4350
rect 19070 4338 19122 4350
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 18274 4286 18286 4338
rect 18338 4286 18350 4338
rect 20178 4286 20190 4338
rect 20242 4286 20254 4338
rect 21522 4286 21534 4338
rect 21586 4286 21598 4338
rect 22194 4286 22206 4338
rect 22258 4286 22270 4338
rect 15598 4274 15650 4286
rect 19070 4274 19122 4286
rect 9102 4226 9154 4238
rect 9102 4162 9154 4174
rect 11342 4226 11394 4238
rect 11342 4162 11394 4174
rect 11790 4226 11842 4238
rect 16830 4226 16882 4238
rect 12786 4174 12798 4226
rect 12850 4174 12862 4226
rect 14130 4174 14142 4226
rect 14194 4174 14206 4226
rect 26450 4174 26462 4226
rect 26514 4174 26526 4226
rect 11790 4162 11842 4174
rect 16830 4162 16882 4174
rect 1344 3946 28560 3980
rect 1344 3894 4616 3946
rect 4668 3894 4720 3946
rect 4772 3894 4824 3946
rect 4876 3894 11420 3946
rect 11472 3894 11524 3946
rect 11576 3894 11628 3946
rect 11680 3894 18224 3946
rect 18276 3894 18328 3946
rect 18380 3894 18432 3946
rect 18484 3894 25028 3946
rect 25080 3894 25132 3946
rect 25184 3894 25236 3946
rect 25288 3894 28560 3946
rect 1344 3860 28560 3894
rect 27358 3778 27410 3790
rect 27358 3714 27410 3726
rect 24670 3666 24722 3678
rect 15586 3614 15598 3666
rect 15650 3614 15662 3666
rect 17378 3614 17390 3666
rect 17442 3614 17454 3666
rect 19394 3614 19406 3666
rect 19458 3614 19470 3666
rect 23202 3614 23214 3666
rect 23266 3614 23278 3666
rect 25666 3614 25678 3666
rect 25730 3614 25742 3666
rect 24670 3602 24722 3614
rect 11230 3554 11282 3566
rect 13582 3554 13634 3566
rect 8642 3502 8654 3554
rect 8706 3502 8718 3554
rect 10434 3502 10446 3554
rect 10498 3502 10510 3554
rect 11778 3502 11790 3554
rect 11842 3502 11854 3554
rect 11230 3490 11282 3502
rect 13582 3490 13634 3502
rect 15150 3554 15202 3566
rect 15150 3490 15202 3502
rect 16942 3554 16994 3566
rect 16942 3490 16994 3502
rect 18958 3554 19010 3566
rect 22430 3554 22482 3566
rect 25006 3554 25058 3566
rect 20850 3502 20862 3554
rect 20914 3502 20926 3554
rect 21522 3502 21534 3554
rect 21586 3502 21598 3554
rect 22866 3502 22878 3554
rect 22930 3502 22942 3554
rect 18958 3490 19010 3502
rect 22430 3490 22482 3502
rect 25006 3490 25058 3502
rect 26574 3554 26626 3566
rect 26574 3490 26626 3502
rect 10894 3442 10946 3454
rect 10894 3378 10946 3390
rect 12238 3442 12290 3454
rect 12238 3378 12290 3390
rect 12574 3442 12626 3454
rect 12574 3378 12626 3390
rect 13246 3442 13298 3454
rect 13246 3378 13298 3390
rect 18398 3442 18450 3454
rect 18398 3378 18450 3390
rect 20302 3442 20354 3454
rect 20302 3378 20354 3390
rect 21086 3442 21138 3454
rect 21086 3378 21138 3390
rect 21758 3442 21810 3454
rect 21758 3378 21810 3390
rect 22094 3442 22146 3454
rect 22094 3378 22146 3390
rect 24110 3442 24162 3454
rect 24110 3378 24162 3390
rect 6750 3330 6802 3342
rect 6750 3266 6802 3278
rect 7198 3330 7250 3342
rect 7198 3266 7250 3278
rect 7982 3330 8034 3342
rect 7982 3266 8034 3278
rect 9774 3330 9826 3342
rect 9774 3266 9826 3278
rect 11566 3330 11618 3342
rect 11566 3266 11618 3278
rect 14366 3330 14418 3342
rect 14366 3266 14418 3278
rect 1344 3162 28720 3196
rect 1344 3110 8018 3162
rect 8070 3110 8122 3162
rect 8174 3110 8226 3162
rect 8278 3110 14822 3162
rect 14874 3110 14926 3162
rect 14978 3110 15030 3162
rect 15082 3110 21626 3162
rect 21678 3110 21730 3162
rect 21782 3110 21834 3162
rect 21886 3110 28430 3162
rect 28482 3110 28534 3162
rect 28586 3110 28638 3162
rect 28690 3110 28720 3162
rect 1344 3076 28720 3110
<< via1 >>
rect 2046 26798 2098 26850
rect 2606 26798 2658 26850
rect 13470 26798 13522 26850
rect 14142 26798 14194 26850
rect 18846 26798 18898 26850
rect 20078 26798 20130 26850
rect 20302 26798 20354 26850
rect 21198 26798 21250 26850
rect 22206 26798 22258 26850
rect 22878 26798 22930 26850
rect 24222 26798 24274 26850
rect 24782 26798 24834 26850
rect 8018 26630 8070 26682
rect 8122 26630 8174 26682
rect 8226 26630 8278 26682
rect 14822 26630 14874 26682
rect 14926 26630 14978 26682
rect 15030 26630 15082 26682
rect 21626 26630 21678 26682
rect 21730 26630 21782 26682
rect 21834 26630 21886 26682
rect 28430 26630 28482 26682
rect 28534 26630 28586 26682
rect 28638 26630 28690 26682
rect 15486 26462 15538 26514
rect 20078 26462 20130 26514
rect 24110 26462 24162 26514
rect 26126 26462 26178 26514
rect 2606 26350 2658 26402
rect 4286 26350 4338 26402
rect 4958 26350 5010 26402
rect 7870 26350 7922 26402
rect 10670 26350 10722 26402
rect 12238 26350 12290 26402
rect 15710 26350 15762 26402
rect 3390 26238 3442 26290
rect 4062 26238 4114 26290
rect 4734 26238 4786 26290
rect 6862 26238 6914 26290
rect 8542 26238 8594 26290
rect 9998 26238 10050 26290
rect 11342 26238 11394 26290
rect 13694 26238 13746 26290
rect 15934 26238 15986 26290
rect 16942 26238 16994 26290
rect 18622 26238 18674 26290
rect 20750 26238 20802 26290
rect 22430 26238 22482 26290
rect 24558 26238 24610 26290
rect 26574 26238 26626 26290
rect 5854 26126 5906 26178
rect 14142 26126 14194 26178
rect 17390 26126 17442 26178
rect 18958 26126 19010 26178
rect 21198 26126 21250 26178
rect 22766 26126 22818 26178
rect 25006 26126 25058 26178
rect 27694 26126 27746 26178
rect 4616 25846 4668 25898
rect 4720 25846 4772 25898
rect 4824 25846 4876 25898
rect 11420 25846 11472 25898
rect 11524 25846 11576 25898
rect 11628 25846 11680 25898
rect 18224 25846 18276 25898
rect 18328 25846 18380 25898
rect 18432 25846 18484 25898
rect 25028 25846 25080 25898
rect 25132 25846 25184 25898
rect 25236 25846 25288 25898
rect 10558 25678 10610 25730
rect 1822 25566 1874 25618
rect 5070 25566 5122 25618
rect 6078 25566 6130 25618
rect 8766 25566 8818 25618
rect 12126 25566 12178 25618
rect 13918 25566 13970 25618
rect 14814 25566 14866 25618
rect 16830 25566 16882 25618
rect 18846 25566 18898 25618
rect 19630 25566 19682 25618
rect 20862 25566 20914 25618
rect 22878 25566 22930 25618
rect 25902 25566 25954 25618
rect 3614 25454 3666 25506
rect 6302 25454 6354 25506
rect 6974 25454 7026 25506
rect 7646 25454 7698 25506
rect 8990 25454 9042 25506
rect 11790 25454 11842 25506
rect 15038 25454 15090 25506
rect 17278 25454 17330 25506
rect 18510 25454 18562 25506
rect 20190 25454 20242 25506
rect 21310 25454 21362 25506
rect 23662 25454 23714 25506
rect 24222 25454 24274 25506
rect 24894 25454 24946 25506
rect 3950 25342 4002 25394
rect 4286 25342 4338 25394
rect 6638 25342 6690 25394
rect 7310 25342 7362 25394
rect 7982 25342 8034 25394
rect 2158 25230 2210 25282
rect 2942 25230 2994 25282
rect 4622 25230 4674 25282
rect 9326 25230 9378 25282
rect 11342 25230 11394 25282
rect 13470 25230 13522 25282
rect 15374 25230 15426 25282
rect 17054 25230 17106 25282
rect 19966 25230 20018 25282
rect 21646 25230 21698 25282
rect 22430 25230 22482 25282
rect 23998 25230 24050 25282
rect 24670 25230 24722 25282
rect 25342 25230 25394 25282
rect 26910 25230 26962 25282
rect 27694 25230 27746 25282
rect 8018 25062 8070 25114
rect 8122 25062 8174 25114
rect 8226 25062 8278 25114
rect 14822 25062 14874 25114
rect 14926 25062 14978 25114
rect 15030 25062 15082 25114
rect 21626 25062 21678 25114
rect 21730 25062 21782 25114
rect 21834 25062 21886 25114
rect 28430 25062 28482 25114
rect 28534 25062 28586 25114
rect 28638 25062 28690 25114
rect 3278 24894 3330 24946
rect 3502 24894 3554 24946
rect 4286 24894 4338 24946
rect 4734 24894 4786 24946
rect 6078 24894 6130 24946
rect 7422 24894 7474 24946
rect 10446 24894 10498 24946
rect 25454 24894 25506 24946
rect 2046 24782 2098 24834
rect 2382 24782 2434 24834
rect 9662 24782 9714 24834
rect 14366 24782 14418 24834
rect 23326 24782 23378 24834
rect 23998 24782 24050 24834
rect 24334 24782 24386 24834
rect 1822 24670 1874 24722
rect 3726 24670 3778 24722
rect 14590 24670 14642 24722
rect 23102 24670 23154 24722
rect 23774 24670 23826 24722
rect 24670 24670 24722 24722
rect 26574 24670 26626 24722
rect 26910 24670 26962 24722
rect 14142 24558 14194 24610
rect 22766 24558 22818 24610
rect 26126 24558 26178 24610
rect 28030 24558 28082 24610
rect 4616 24278 4668 24330
rect 4720 24278 4772 24330
rect 4824 24278 4876 24330
rect 11420 24278 11472 24330
rect 11524 24278 11576 24330
rect 11628 24278 11680 24330
rect 18224 24278 18276 24330
rect 18328 24278 18380 24330
rect 18432 24278 18484 24330
rect 25028 24278 25080 24330
rect 25132 24278 25184 24330
rect 25236 24278 25288 24330
rect 27694 24110 27746 24162
rect 23662 23998 23714 24050
rect 8430 23886 8482 23938
rect 9214 23886 9266 23938
rect 9662 23886 9714 23938
rect 10670 23886 10722 23938
rect 11006 23886 11058 23938
rect 11902 23886 11954 23938
rect 13806 23886 13858 23938
rect 15038 23886 15090 23938
rect 15598 23886 15650 23938
rect 16494 23886 16546 23938
rect 19854 23886 19906 23938
rect 20526 23886 20578 23938
rect 21422 23886 21474 23938
rect 23998 23886 24050 23938
rect 25230 23886 25282 23938
rect 25902 23886 25954 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 8654 23774 8706 23826
rect 9998 23774 10050 23826
rect 10334 23774 10386 23826
rect 11342 23774 11394 23826
rect 11678 23774 11730 23826
rect 13470 23774 13522 23826
rect 15262 23774 15314 23826
rect 15934 23774 15986 23826
rect 16830 23774 16882 23826
rect 20078 23774 20130 23826
rect 20750 23774 20802 23826
rect 21646 23774 21698 23826
rect 24222 23774 24274 23826
rect 24558 23774 24610 23826
rect 24894 23774 24946 23826
rect 25566 23774 25618 23826
rect 26238 23774 26290 23826
rect 2494 23662 2546 23714
rect 8990 23662 9042 23714
rect 26910 23662 26962 23714
rect 8018 23494 8070 23546
rect 8122 23494 8174 23546
rect 8226 23494 8278 23546
rect 14822 23494 14874 23546
rect 14926 23494 14978 23546
rect 15030 23494 15082 23546
rect 21626 23494 21678 23546
rect 21730 23494 21782 23546
rect 21834 23494 21886 23546
rect 28430 23494 28482 23546
rect 28534 23494 28586 23546
rect 28638 23494 28690 23546
rect 9550 23326 9602 23378
rect 10558 23326 10610 23378
rect 10894 23326 10946 23378
rect 20862 23326 20914 23378
rect 25566 23326 25618 23378
rect 10222 23214 10274 23266
rect 24670 23214 24722 23266
rect 26238 23214 26290 23266
rect 26910 23214 26962 23266
rect 9774 23102 9826 23154
rect 11118 23102 11170 23154
rect 20638 23102 20690 23154
rect 24446 23102 24498 23154
rect 25342 23102 25394 23154
rect 26014 23102 26066 23154
rect 27470 22990 27522 23042
rect 28254 22990 28306 23042
rect 4616 22710 4668 22762
rect 4720 22710 4772 22762
rect 4824 22710 4876 22762
rect 11420 22710 11472 22762
rect 11524 22710 11576 22762
rect 11628 22710 11680 22762
rect 18224 22710 18276 22762
rect 18328 22710 18380 22762
rect 18432 22710 18484 22762
rect 25028 22710 25080 22762
rect 25132 22710 25184 22762
rect 25236 22710 25288 22762
rect 25678 22318 25730 22370
rect 26910 22318 26962 22370
rect 26238 22206 26290 22258
rect 26574 22206 26626 22258
rect 28030 22206 28082 22258
rect 25902 22094 25954 22146
rect 8018 21926 8070 21978
rect 8122 21926 8174 21978
rect 8226 21926 8278 21978
rect 14822 21926 14874 21978
rect 14926 21926 14978 21978
rect 15030 21926 15082 21978
rect 21626 21926 21678 21978
rect 21730 21926 21782 21978
rect 21834 21926 21886 21978
rect 28430 21926 28482 21978
rect 28534 21926 28586 21978
rect 28638 21926 28690 21978
rect 26462 21758 26514 21810
rect 27806 21758 27858 21810
rect 14814 21646 14866 21698
rect 26798 21646 26850 21698
rect 27134 21646 27186 21698
rect 27470 21534 27522 21586
rect 28142 21534 28194 21586
rect 13806 21422 13858 21474
rect 26238 21422 26290 21474
rect 4616 21142 4668 21194
rect 4720 21142 4772 21194
rect 4824 21142 4876 21194
rect 11420 21142 11472 21194
rect 11524 21142 11576 21194
rect 11628 21142 11680 21194
rect 18224 21142 18276 21194
rect 18328 21142 18380 21194
rect 18432 21142 18484 21194
rect 25028 21142 25080 21194
rect 25132 21142 25184 21194
rect 25236 21142 25288 21194
rect 16270 20862 16322 20914
rect 24446 20862 24498 20914
rect 26686 20862 26738 20914
rect 26910 20750 26962 20802
rect 17278 20638 17330 20690
rect 25454 20638 25506 20690
rect 28030 20638 28082 20690
rect 23998 20526 24050 20578
rect 8018 20358 8070 20410
rect 8122 20358 8174 20410
rect 8226 20358 8278 20410
rect 14822 20358 14874 20410
rect 14926 20358 14978 20410
rect 15030 20358 15082 20410
rect 21626 20358 21678 20410
rect 21730 20358 21782 20410
rect 21834 20358 21886 20410
rect 28430 20358 28482 20410
rect 28534 20358 28586 20410
rect 28638 20358 28690 20410
rect 20526 20190 20578 20242
rect 14590 20078 14642 20130
rect 15374 20078 15426 20130
rect 23550 20078 23602 20130
rect 27806 20078 27858 20130
rect 9886 19966 9938 20018
rect 11902 19966 11954 20018
rect 12350 19966 12402 20018
rect 15822 19966 15874 20018
rect 17614 19966 17666 20018
rect 18062 19966 18114 20018
rect 21086 19966 21138 20018
rect 24446 19966 24498 20018
rect 28142 19966 28194 20018
rect 21534 19854 21586 19906
rect 21870 19854 21922 19906
rect 22318 19854 22370 19906
rect 25454 19854 25506 19906
rect 25902 19854 25954 19906
rect 26238 19854 26290 19906
rect 27582 19854 27634 19906
rect 9550 19742 9602 19794
rect 16382 19742 16434 19794
rect 24110 19742 24162 19794
rect 25454 19742 25506 19794
rect 25902 19742 25954 19794
rect 4616 19574 4668 19626
rect 4720 19574 4772 19626
rect 4824 19574 4876 19626
rect 11420 19574 11472 19626
rect 11524 19574 11576 19626
rect 11628 19574 11680 19626
rect 18224 19574 18276 19626
rect 18328 19574 18380 19626
rect 18432 19574 18484 19626
rect 25028 19574 25080 19626
rect 25132 19574 25184 19626
rect 25236 19574 25288 19626
rect 13022 19406 13074 19458
rect 14030 19406 14082 19458
rect 21310 19406 21362 19458
rect 7646 19294 7698 19346
rect 19182 19294 19234 19346
rect 9550 19182 9602 19234
rect 9998 19182 10050 19234
rect 13470 19182 13522 19234
rect 14254 19182 14306 19234
rect 14926 19182 14978 19234
rect 21534 19182 21586 19234
rect 22430 19182 22482 19234
rect 22878 19182 22930 19234
rect 26350 19182 26402 19234
rect 8990 19070 9042 19122
rect 17166 19070 17218 19122
rect 17950 19070 18002 19122
rect 20190 19070 20242 19122
rect 27806 19070 27858 19122
rect 28142 19070 28194 19122
rect 12238 18958 12290 19010
rect 25118 18958 25170 19010
rect 25902 18958 25954 19010
rect 26126 18958 26178 19010
rect 27582 18958 27634 19010
rect 8018 18790 8070 18842
rect 8122 18790 8174 18842
rect 8226 18790 8278 18842
rect 14822 18790 14874 18842
rect 14926 18790 14978 18842
rect 15030 18790 15082 18842
rect 21626 18790 21678 18842
rect 21730 18790 21782 18842
rect 21834 18790 21886 18842
rect 28430 18790 28482 18842
rect 28534 18790 28586 18842
rect 28638 18790 28690 18842
rect 8542 18622 8594 18674
rect 23214 18622 23266 18674
rect 24670 18622 24722 18674
rect 12574 18510 12626 18562
rect 16158 18510 16210 18562
rect 19406 18510 19458 18562
rect 25902 18510 25954 18562
rect 5518 18398 5570 18450
rect 6078 18398 6130 18450
rect 9886 18398 9938 18450
rect 13246 18398 13298 18450
rect 13918 18398 13970 18450
rect 16942 18398 16994 18450
rect 20190 18398 20242 18450
rect 20750 18398 20802 18450
rect 23774 18398 23826 18450
rect 24446 18398 24498 18450
rect 11566 18286 11618 18338
rect 18398 18286 18450 18338
rect 25342 18286 25394 18338
rect 27134 18286 27186 18338
rect 27694 18286 27746 18338
rect 9102 18174 9154 18226
rect 10222 18174 10274 18226
rect 4616 18006 4668 18058
rect 4720 18006 4772 18058
rect 4824 18006 4876 18058
rect 11420 18006 11472 18058
rect 11524 18006 11576 18058
rect 11628 18006 11680 18058
rect 18224 18006 18276 18058
rect 18328 18006 18380 18058
rect 18432 18006 18484 18058
rect 25028 18006 25080 18058
rect 25132 18006 25184 18058
rect 25236 18006 25288 18058
rect 11230 17838 11282 17890
rect 12014 17838 12066 17890
rect 15822 17838 15874 17890
rect 21422 17726 21474 17778
rect 23102 17726 23154 17778
rect 4510 17614 4562 17666
rect 5630 17614 5682 17666
rect 7534 17614 7586 17666
rect 8206 17614 8258 17666
rect 11678 17614 11730 17666
rect 13694 17614 13746 17666
rect 15710 17614 15762 17666
rect 16158 17614 16210 17666
rect 16830 17614 16882 17666
rect 20638 17614 20690 17666
rect 22654 17614 22706 17666
rect 26350 17614 26402 17666
rect 27022 17614 27074 17666
rect 28142 17614 28194 17666
rect 10446 17502 10498 17554
rect 27806 17502 27858 17554
rect 3950 17390 4002 17442
rect 4958 17390 5010 17442
rect 6190 17390 6242 17442
rect 6638 17390 6690 17442
rect 13806 17390 13858 17442
rect 19294 17390 19346 17442
rect 19854 17390 19906 17442
rect 20078 17390 20130 17442
rect 22542 17390 22594 17442
rect 23326 17390 23378 17442
rect 23886 17390 23938 17442
rect 27358 17390 27410 17442
rect 8018 17222 8070 17274
rect 8122 17222 8174 17274
rect 8226 17222 8278 17274
rect 14822 17222 14874 17274
rect 14926 17222 14978 17274
rect 15030 17222 15082 17274
rect 21626 17222 21678 17274
rect 21730 17222 21782 17274
rect 21834 17222 21886 17274
rect 28430 17222 28482 17274
rect 28534 17222 28586 17274
rect 28638 17222 28690 17274
rect 2270 17054 2322 17106
rect 9102 17054 9154 17106
rect 21646 17054 21698 17106
rect 8318 16942 8370 16994
rect 9774 16942 9826 16994
rect 20862 16942 20914 16994
rect 23998 16942 24050 16994
rect 27694 16942 27746 16994
rect 4622 16830 4674 16882
rect 5070 16830 5122 16882
rect 5518 16830 5570 16882
rect 6078 16830 6130 16882
rect 14590 16830 14642 16882
rect 17950 16830 18002 16882
rect 18622 16830 18674 16882
rect 21982 16830 22034 16882
rect 22430 16830 22482 16882
rect 22878 16718 22930 16770
rect 26686 16718 26738 16770
rect 1598 16606 1650 16658
rect 4616 16438 4668 16490
rect 4720 16438 4772 16490
rect 4824 16438 4876 16490
rect 11420 16438 11472 16490
rect 11524 16438 11576 16490
rect 11628 16438 11680 16490
rect 18224 16438 18276 16490
rect 18328 16438 18380 16490
rect 18432 16438 18484 16490
rect 25028 16438 25080 16490
rect 25132 16438 25184 16490
rect 25236 16438 25288 16490
rect 3950 16158 4002 16210
rect 6974 16158 7026 16210
rect 9774 16158 9826 16210
rect 14702 16158 14754 16210
rect 19294 16158 19346 16210
rect 21982 16046 22034 16098
rect 2718 15934 2770 15986
rect 7982 15934 8034 15986
rect 10782 15934 10834 15986
rect 13582 15934 13634 15986
rect 20302 15934 20354 15986
rect 25790 15934 25842 15986
rect 8018 15654 8070 15706
rect 8122 15654 8174 15706
rect 8226 15654 8278 15706
rect 14822 15654 14874 15706
rect 14926 15654 14978 15706
rect 15030 15654 15082 15706
rect 21626 15654 21678 15706
rect 21730 15654 21782 15706
rect 21834 15654 21886 15706
rect 28430 15654 28482 15706
rect 28534 15654 28586 15706
rect 28638 15654 28690 15706
rect 6302 15486 6354 15538
rect 7086 15486 7138 15538
rect 8430 15486 8482 15538
rect 12014 15486 12066 15538
rect 12798 15486 12850 15538
rect 22766 15486 22818 15538
rect 27246 15374 27298 15426
rect 2718 15262 2770 15314
rect 3614 15262 3666 15314
rect 3950 15262 4002 15314
rect 8990 15262 9042 15314
rect 11454 15262 11506 15314
rect 15038 15262 15090 15314
rect 15710 15262 15762 15314
rect 16046 15262 16098 15314
rect 20078 15262 20130 15314
rect 20526 15262 20578 15314
rect 24558 15262 24610 15314
rect 2046 15150 2098 15202
rect 2606 15150 2658 15202
rect 25342 15150 25394 15202
rect 25790 15150 25842 15202
rect 26238 15150 26290 15202
rect 11230 15038 11282 15090
rect 23550 15038 23602 15090
rect 24446 15038 24498 15090
rect 4616 14870 4668 14922
rect 4720 14870 4772 14922
rect 4824 14870 4876 14922
rect 11420 14870 11472 14922
rect 11524 14870 11576 14922
rect 11628 14870 11680 14922
rect 18224 14870 18276 14922
rect 18328 14870 18380 14922
rect 18432 14870 18484 14922
rect 25028 14870 25080 14922
rect 25132 14870 25184 14922
rect 25236 14870 25288 14922
rect 2270 14702 2322 14754
rect 20750 14702 20802 14754
rect 25566 14702 25618 14754
rect 4062 14590 4114 14642
rect 14478 14590 14530 14642
rect 25902 14590 25954 14642
rect 2046 14478 2098 14530
rect 8654 14478 8706 14530
rect 9214 14478 9266 14530
rect 9550 14478 9602 14530
rect 9886 14478 9938 14530
rect 20526 14478 20578 14530
rect 22094 14478 22146 14530
rect 22542 14478 22594 14530
rect 26350 14478 26402 14530
rect 27134 14478 27186 14530
rect 28142 14478 28194 14530
rect 3054 14366 3106 14418
rect 5518 14366 5570 14418
rect 13022 14366 13074 14418
rect 15486 14366 15538 14418
rect 24782 14366 24834 14418
rect 4510 14254 4562 14306
rect 6078 14254 6130 14306
rect 12462 14254 12514 14306
rect 19854 14254 19906 14306
rect 26686 14254 26738 14306
rect 27694 14254 27746 14306
rect 8018 14086 8070 14138
rect 8122 14086 8174 14138
rect 8226 14086 8278 14138
rect 14822 14086 14874 14138
rect 14926 14086 14978 14138
rect 15030 14086 15082 14138
rect 21626 14086 21678 14138
rect 21730 14086 21782 14138
rect 21834 14086 21886 14138
rect 28430 14086 28482 14138
rect 28534 14086 28586 14138
rect 28638 14086 28690 14138
rect 2606 13918 2658 13970
rect 24222 13918 24274 13970
rect 25454 13918 25506 13970
rect 6974 13806 7026 13858
rect 18846 13806 18898 13858
rect 27246 13806 27298 13858
rect 5070 13694 5122 13746
rect 5742 13694 5794 13746
rect 10110 13694 10162 13746
rect 10894 13694 10946 13746
rect 14478 13694 14530 13746
rect 21310 13694 21362 13746
rect 21758 13694 21810 13746
rect 7982 13582 8034 13634
rect 19854 13582 19906 13634
rect 26014 13582 26066 13634
rect 26238 13582 26290 13634
rect 2046 13470 2098 13522
rect 10446 13470 10498 13522
rect 13918 13470 13970 13522
rect 24782 13470 24834 13522
rect 4616 13302 4668 13354
rect 4720 13302 4772 13354
rect 4824 13302 4876 13354
rect 11420 13302 11472 13354
rect 11524 13302 11576 13354
rect 11628 13302 11680 13354
rect 18224 13302 18276 13354
rect 18328 13302 18380 13354
rect 18432 13302 18484 13354
rect 25028 13302 25080 13354
rect 25132 13302 25184 13354
rect 25236 13302 25288 13354
rect 9102 13134 9154 13186
rect 13470 13134 13522 13186
rect 4062 13022 4114 13074
rect 7870 13022 7922 13074
rect 16830 13022 16882 13074
rect 27134 13022 27186 13074
rect 12238 12910 12290 12962
rect 12574 12910 12626 12962
rect 13918 12910 13970 12962
rect 15150 12910 15202 12962
rect 23214 12910 23266 12962
rect 23662 12910 23714 12962
rect 2718 12798 2770 12850
rect 6526 12798 6578 12850
rect 9886 12798 9938 12850
rect 25902 12798 25954 12850
rect 26686 12686 26738 12738
rect 8018 12518 8070 12570
rect 8122 12518 8174 12570
rect 8226 12518 8278 12570
rect 14822 12518 14874 12570
rect 14926 12518 14978 12570
rect 15030 12518 15082 12570
rect 21626 12518 21678 12570
rect 21730 12518 21782 12570
rect 21834 12518 21886 12570
rect 28430 12518 28482 12570
rect 28534 12518 28586 12570
rect 28638 12518 28690 12570
rect 5406 12350 5458 12402
rect 15262 12350 15314 12402
rect 19742 12350 19794 12402
rect 2382 12238 2434 12290
rect 6190 12238 6242 12290
rect 20526 12238 20578 12290
rect 27358 12238 27410 12290
rect 4622 12126 4674 12178
rect 5294 12126 5346 12178
rect 8430 12126 8482 12178
rect 9102 12126 9154 12178
rect 14590 12126 14642 12178
rect 22878 12126 22930 12178
rect 23438 12126 23490 12178
rect 24558 12126 24610 12178
rect 10782 12014 10834 12066
rect 25342 12014 25394 12066
rect 26462 12014 26514 12066
rect 1598 11902 1650 11954
rect 24110 11902 24162 11954
rect 4616 11734 4668 11786
rect 4720 11734 4772 11786
rect 4824 11734 4876 11786
rect 11420 11734 11472 11786
rect 11524 11734 11576 11786
rect 11628 11734 11680 11786
rect 18224 11734 18276 11786
rect 18328 11734 18380 11786
rect 18432 11734 18484 11786
rect 25028 11734 25080 11786
rect 25132 11734 25184 11786
rect 25236 11734 25288 11786
rect 3838 11454 3890 11506
rect 18062 11454 18114 11506
rect 1822 11342 1874 11394
rect 6302 11342 6354 11394
rect 7310 11342 7362 11394
rect 7758 11342 7810 11394
rect 8094 11342 8146 11394
rect 14142 11342 14194 11394
rect 14478 11342 14530 11394
rect 20302 11342 20354 11394
rect 21982 11342 22034 11394
rect 27358 11342 27410 11394
rect 2718 11230 2770 11282
rect 10446 11230 10498 11282
rect 13806 11230 13858 11282
rect 24334 11230 24386 11282
rect 2046 11118 2098 11170
rect 6862 11118 6914 11170
rect 11230 11118 11282 11170
rect 20750 11118 20802 11170
rect 26910 11118 26962 11170
rect 8018 10950 8070 11002
rect 8122 10950 8174 11002
rect 8226 10950 8278 11002
rect 14822 10950 14874 11002
rect 14926 10950 14978 11002
rect 15030 10950 15082 11002
rect 21626 10950 21678 11002
rect 21730 10950 21782 11002
rect 21834 10950 21886 11002
rect 28430 10950 28482 11002
rect 28534 10950 28586 11002
rect 28638 10950 28690 11002
rect 1822 10782 1874 10834
rect 6974 10782 7026 10834
rect 8094 10782 8146 10834
rect 22318 10782 22370 10834
rect 23774 10782 23826 10834
rect 15822 10670 15874 10722
rect 23102 10670 23154 10722
rect 27246 10670 27298 10722
rect 2942 10558 2994 10610
rect 3278 10558 3330 10610
rect 4286 10558 4338 10610
rect 4734 10558 4786 10610
rect 8542 10558 8594 10610
rect 13470 10558 13522 10610
rect 18286 10558 18338 10610
rect 19630 10558 19682 10610
rect 19966 10558 20018 10610
rect 23886 10558 23938 10610
rect 3726 10446 3778 10498
rect 9886 10446 9938 10498
rect 14814 10446 14866 10498
rect 24334 10446 24386 10498
rect 26238 10446 26290 10498
rect 7758 10334 7810 10386
rect 18062 10334 18114 10386
rect 4616 10166 4668 10218
rect 4720 10166 4772 10218
rect 4824 10166 4876 10218
rect 11420 10166 11472 10218
rect 11524 10166 11576 10218
rect 11628 10166 11680 10218
rect 18224 10166 18276 10218
rect 18328 10166 18380 10218
rect 18432 10166 18484 10218
rect 25028 10166 25080 10218
rect 25132 10166 25184 10218
rect 25236 10166 25288 10218
rect 12686 9998 12738 10050
rect 17502 9998 17554 10050
rect 3838 9886 3890 9938
rect 6638 9886 6690 9938
rect 8430 9886 8482 9938
rect 8990 9886 9042 9938
rect 19070 9886 19122 9938
rect 27470 9886 27522 9938
rect 6190 9774 6242 9826
rect 10334 9774 10386 9826
rect 14142 9774 14194 9826
rect 21534 9774 21586 9826
rect 21982 9774 22034 9826
rect 4958 9662 5010 9714
rect 7534 9662 7586 9714
rect 20414 9662 20466 9714
rect 26350 9662 26402 9714
rect 5630 9550 5682 9602
rect 24446 9550 24498 9602
rect 25006 9550 25058 9602
rect 25342 9550 25394 9602
rect 8018 9382 8070 9434
rect 8122 9382 8174 9434
rect 8226 9382 8278 9434
rect 14822 9382 14874 9434
rect 14926 9382 14978 9434
rect 15030 9382 15082 9434
rect 21626 9382 21678 9434
rect 21730 9382 21782 9434
rect 21834 9382 21886 9434
rect 28430 9382 28482 9434
rect 28534 9382 28586 9434
rect 28638 9382 28690 9434
rect 5630 9214 5682 9266
rect 15374 9214 15426 9266
rect 16270 9214 16322 9266
rect 20190 9102 20242 9154
rect 21870 9102 21922 9154
rect 27246 9102 27298 9154
rect 2718 8990 2770 9042
rect 3390 8990 3442 9042
rect 12238 8990 12290 9042
rect 12910 8990 12962 9042
rect 15934 8990 15986 9042
rect 17278 8990 17330 9042
rect 17950 8990 18002 9042
rect 24110 8990 24162 9042
rect 24670 8990 24722 9042
rect 16158 8878 16210 8930
rect 25342 8878 25394 8930
rect 26238 8878 26290 8930
rect 6414 8766 6466 8818
rect 20974 8766 21026 8818
rect 21086 8766 21138 8818
rect 4616 8598 4668 8650
rect 4720 8598 4772 8650
rect 4824 8598 4876 8650
rect 11420 8598 11472 8650
rect 11524 8598 11576 8650
rect 11628 8598 11680 8650
rect 18224 8598 18276 8650
rect 18328 8598 18380 8650
rect 18432 8598 18484 8650
rect 25028 8598 25080 8650
rect 25132 8598 25184 8650
rect 25236 8598 25288 8650
rect 4510 8430 4562 8482
rect 22766 8430 22818 8482
rect 5854 8318 5906 8370
rect 6750 8318 6802 8370
rect 19294 8318 19346 8370
rect 23550 8318 23602 8370
rect 4846 8206 4898 8258
rect 14926 8206 14978 8258
rect 15374 8206 15426 8258
rect 19070 8206 19122 8258
rect 21422 8206 21474 8258
rect 22990 8206 23042 8258
rect 26686 8206 26738 8258
rect 27134 8206 27186 8258
rect 27470 8206 27522 8258
rect 7758 8094 7810 8146
rect 17838 7982 17890 8034
rect 18398 7982 18450 8034
rect 20750 7982 20802 8034
rect 21982 7982 22034 8034
rect 24222 7982 24274 8034
rect 27582 7982 27634 8034
rect 8018 7814 8070 7866
rect 8122 7814 8174 7866
rect 8226 7814 8278 7866
rect 14822 7814 14874 7866
rect 14926 7814 14978 7866
rect 15030 7814 15082 7866
rect 21626 7814 21678 7866
rect 21730 7814 21782 7866
rect 21834 7814 21886 7866
rect 28430 7814 28482 7866
rect 28534 7814 28586 7866
rect 28638 7814 28690 7866
rect 4734 7646 4786 7698
rect 5518 7646 5570 7698
rect 13694 7646 13746 7698
rect 18510 7646 18562 7698
rect 22206 7646 22258 7698
rect 27246 7534 27298 7586
rect 2046 7422 2098 7474
rect 2382 7422 2434 7474
rect 10782 7422 10834 7474
rect 11230 7422 11282 7474
rect 19294 7422 19346 7474
rect 19966 7422 20018 7474
rect 24334 7422 24386 7474
rect 23326 7310 23378 7362
rect 26238 7310 26290 7362
rect 28142 7310 28194 7362
rect 14254 7198 14306 7250
rect 22990 7198 23042 7250
rect 24558 7198 24610 7250
rect 4616 7030 4668 7082
rect 4720 7030 4772 7082
rect 4824 7030 4876 7082
rect 11420 7030 11472 7082
rect 11524 7030 11576 7082
rect 11628 7030 11680 7082
rect 18224 7030 18276 7082
rect 18328 7030 18380 7082
rect 18432 7030 18484 7082
rect 25028 7030 25080 7082
rect 25132 7030 25184 7082
rect 25236 7030 25288 7082
rect 14478 6750 14530 6802
rect 17278 6750 17330 6802
rect 22654 6638 22706 6690
rect 23326 6638 23378 6690
rect 27694 6638 27746 6690
rect 15486 6526 15538 6578
rect 18622 6526 18674 6578
rect 1710 6414 1762 6466
rect 25790 6414 25842 6466
rect 26350 6414 26402 6466
rect 26910 6414 26962 6466
rect 28142 6414 28194 6466
rect 8018 6246 8070 6298
rect 8122 6246 8174 6298
rect 8226 6246 8278 6298
rect 14822 6246 14874 6298
rect 14926 6246 14978 6298
rect 15030 6246 15082 6298
rect 21626 6246 21678 6298
rect 21730 6246 21782 6298
rect 21834 6246 21886 6298
rect 28430 6246 28482 6298
rect 28534 6246 28586 6298
rect 28638 6246 28690 6298
rect 20302 5966 20354 6018
rect 23102 5966 23154 6018
rect 24670 5966 24722 6018
rect 27246 5966 27298 6018
rect 24334 5854 24386 5906
rect 19518 5742 19570 5794
rect 22094 5742 22146 5794
rect 26238 5742 26290 5794
rect 4616 5462 4668 5514
rect 4720 5462 4772 5514
rect 4824 5462 4876 5514
rect 11420 5462 11472 5514
rect 11524 5462 11576 5514
rect 11628 5462 11680 5514
rect 18224 5462 18276 5514
rect 18328 5462 18380 5514
rect 18432 5462 18484 5514
rect 25028 5462 25080 5514
rect 25132 5462 25184 5514
rect 25236 5462 25288 5514
rect 26126 5294 26178 5346
rect 27694 5294 27746 5346
rect 28142 5182 28194 5234
rect 9998 5070 10050 5122
rect 12014 5070 12066 5122
rect 12686 5070 12738 5122
rect 18286 5070 18338 5122
rect 21870 5070 21922 5122
rect 22654 5070 22706 5122
rect 23102 5070 23154 5122
rect 26910 5070 26962 5122
rect 10558 4958 10610 5010
rect 10894 4958 10946 5010
rect 11230 4958 11282 5010
rect 13470 4958 13522 5010
rect 14478 4958 14530 5010
rect 25342 4958 25394 5010
rect 10222 4846 10274 4898
rect 11566 4846 11618 4898
rect 12238 4846 12290 4898
rect 12910 4846 12962 4898
rect 13806 4846 13858 4898
rect 14814 4846 14866 4898
rect 17838 4846 17890 4898
rect 18510 4846 18562 4898
rect 20750 4846 20802 4898
rect 22206 4846 22258 4898
rect 26574 4846 26626 4898
rect 8018 4678 8070 4730
rect 8122 4678 8174 4730
rect 8226 4678 8278 4730
rect 14822 4678 14874 4730
rect 14926 4678 14978 4730
rect 15030 4678 15082 4730
rect 21626 4678 21678 4730
rect 21730 4678 21782 4730
rect 21834 4678 21886 4730
rect 28430 4678 28482 4730
rect 28534 4678 28586 4730
rect 28638 4678 28690 4730
rect 10334 4510 10386 4562
rect 12126 4510 12178 4562
rect 13694 4510 13746 4562
rect 15262 4510 15314 4562
rect 18062 4510 18114 4562
rect 18734 4510 18786 4562
rect 24222 4510 24274 4562
rect 24782 4510 24834 4562
rect 8654 4398 8706 4450
rect 9662 4398 9714 4450
rect 9998 4398 10050 4450
rect 17390 4398 17442 4450
rect 20414 4398 20466 4450
rect 20750 4398 20802 4450
rect 21086 4398 21138 4450
rect 21758 4398 21810 4450
rect 22430 4398 22482 4450
rect 22766 4398 22818 4450
rect 23102 4398 23154 4450
rect 23438 4398 23490 4450
rect 27470 4398 27522 4450
rect 10558 4286 10610 4338
rect 14926 4286 14978 4338
rect 15598 4286 15650 4338
rect 17614 4286 17666 4338
rect 18286 4286 18338 4338
rect 19070 4286 19122 4338
rect 20190 4286 20242 4338
rect 21534 4286 21586 4338
rect 22206 4286 22258 4338
rect 9102 4174 9154 4226
rect 11342 4174 11394 4226
rect 11790 4174 11842 4226
rect 12798 4174 12850 4226
rect 14142 4174 14194 4226
rect 16830 4174 16882 4226
rect 26462 4174 26514 4226
rect 4616 3894 4668 3946
rect 4720 3894 4772 3946
rect 4824 3894 4876 3946
rect 11420 3894 11472 3946
rect 11524 3894 11576 3946
rect 11628 3894 11680 3946
rect 18224 3894 18276 3946
rect 18328 3894 18380 3946
rect 18432 3894 18484 3946
rect 25028 3894 25080 3946
rect 25132 3894 25184 3946
rect 25236 3894 25288 3946
rect 27358 3726 27410 3778
rect 15598 3614 15650 3666
rect 17390 3614 17442 3666
rect 19406 3614 19458 3666
rect 23214 3614 23266 3666
rect 24670 3614 24722 3666
rect 25678 3614 25730 3666
rect 8654 3502 8706 3554
rect 10446 3502 10498 3554
rect 11230 3502 11282 3554
rect 11790 3502 11842 3554
rect 13582 3502 13634 3554
rect 15150 3502 15202 3554
rect 16942 3502 16994 3554
rect 18958 3502 19010 3554
rect 20862 3502 20914 3554
rect 21534 3502 21586 3554
rect 22430 3502 22482 3554
rect 22878 3502 22930 3554
rect 25006 3502 25058 3554
rect 26574 3502 26626 3554
rect 10894 3390 10946 3442
rect 12238 3390 12290 3442
rect 12574 3390 12626 3442
rect 13246 3390 13298 3442
rect 18398 3390 18450 3442
rect 20302 3390 20354 3442
rect 21086 3390 21138 3442
rect 21758 3390 21810 3442
rect 22094 3390 22146 3442
rect 24110 3390 24162 3442
rect 6750 3278 6802 3330
rect 7198 3278 7250 3330
rect 7982 3278 8034 3330
rect 9774 3278 9826 3330
rect 11566 3278 11618 3330
rect 14366 3278 14418 3330
rect 8018 3110 8070 3162
rect 8122 3110 8174 3162
rect 8226 3110 8278 3162
rect 14822 3110 14874 3162
rect 14926 3110 14978 3162
rect 15030 3110 15082 3162
rect 21626 3110 21678 3162
rect 21730 3110 21782 3162
rect 21834 3110 21886 3162
rect 28430 3110 28482 3162
rect 28534 3110 28586 3162
rect 28638 3110 28690 3162
<< metal2 >>
rect 1344 29200 1456 30000
rect 2016 29200 2128 30000
rect 2688 29200 2800 30000
rect 3360 29200 3472 30000
rect 4032 29200 4144 30000
rect 4704 29200 4816 30000
rect 5376 29200 5488 30000
rect 6048 29200 6160 30000
rect 6720 29200 6832 30000
rect 7392 29200 7504 30000
rect 8064 29200 8176 30000
rect 8736 29200 8848 30000
rect 9408 29200 9520 30000
rect 10080 29200 10192 30000
rect 10752 29200 10864 30000
rect 11424 29200 11536 30000
rect 12096 29200 12208 30000
rect 12768 29200 12880 30000
rect 13440 29200 13552 30000
rect 14112 29200 14224 30000
rect 14784 29200 14896 30000
rect 15456 29200 15568 30000
rect 16128 29200 16240 30000
rect 16800 29200 16912 30000
rect 17472 29200 17584 30000
rect 18144 29200 18256 30000
rect 18816 29200 18928 30000
rect 19488 29200 19600 30000
rect 20160 29200 20272 30000
rect 20832 29200 20944 30000
rect 21504 29200 21616 30000
rect 22176 29200 22288 30000
rect 22848 29200 22960 30000
rect 23520 29200 23632 30000
rect 24192 29200 24304 30000
rect 24444 29652 24500 29662
rect 1372 26404 1428 29200
rect 2044 26850 2100 29200
rect 2044 26798 2046 26850
rect 2098 26798 2100 26850
rect 2044 26786 2100 26798
rect 2604 26850 2660 26862
rect 2604 26798 2606 26850
rect 2658 26798 2660 26850
rect 1372 26348 1876 26404
rect 1820 25618 1876 26348
rect 2604 26402 2660 26798
rect 2604 26350 2606 26402
rect 2658 26350 2660 26402
rect 2604 26338 2660 26350
rect 1820 25566 1822 25618
rect 1874 25566 1876 25618
rect 1820 24722 1876 25566
rect 2156 25284 2212 25294
rect 2156 25190 2212 25228
rect 2716 25172 2772 29200
rect 3388 26908 3444 29200
rect 3388 26852 3556 26908
rect 3388 26292 3444 26302
rect 3388 26198 3444 26236
rect 3500 25508 3556 26852
rect 4060 26290 4116 29200
rect 4060 26238 4062 26290
rect 4114 26238 4116 26290
rect 4060 25956 4116 26238
rect 4284 26402 4340 26414
rect 4284 26350 4286 26402
rect 4338 26350 4340 26402
rect 4284 26180 4340 26350
rect 4732 26290 4788 29200
rect 4732 26238 4734 26290
rect 4786 26238 4788 26290
rect 4732 26180 4788 26238
rect 4956 26402 5012 26414
rect 4956 26350 4958 26402
rect 5010 26350 5012 26402
rect 4956 26292 5012 26350
rect 4956 26236 5236 26292
rect 4732 26124 5012 26180
rect 4284 26114 4340 26124
rect 4060 25900 4452 25956
rect 3948 25732 4004 25742
rect 3612 25508 3668 25518
rect 3276 25506 3668 25508
rect 3276 25454 3614 25506
rect 3666 25454 3668 25506
rect 3276 25452 3668 25454
rect 2940 25284 2996 25294
rect 2940 25190 2996 25228
rect 2716 25106 2772 25116
rect 3276 24946 3332 25452
rect 3612 25442 3668 25452
rect 3948 25394 4004 25676
rect 3948 25342 3950 25394
rect 4002 25342 4004 25394
rect 3948 25330 4004 25342
rect 4284 25394 4340 25406
rect 4284 25342 4286 25394
rect 4338 25342 4340 25394
rect 3276 24894 3278 24946
rect 3330 24894 3332 24946
rect 3276 24882 3332 24894
rect 3500 25284 3556 25294
rect 3500 24946 3556 25228
rect 3500 24894 3502 24946
rect 3554 24894 3556 24946
rect 3500 24882 3556 24894
rect 4284 25172 4340 25342
rect 4284 24946 4340 25116
rect 4284 24894 4286 24946
rect 4338 24894 4340 24946
rect 4284 24882 4340 24894
rect 4396 24948 4452 25900
rect 4614 25900 4878 25910
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4614 25834 4878 25844
rect 4956 25620 5012 26124
rect 5068 25620 5124 25630
rect 4956 25618 5124 25620
rect 4956 25566 5070 25618
rect 5122 25566 5124 25618
rect 4956 25564 5124 25566
rect 5068 25554 5124 25564
rect 5180 25396 5236 26236
rect 5404 26180 5460 29200
rect 6076 26908 6132 29200
rect 6748 26908 6804 29200
rect 7420 26908 7476 29200
rect 8092 27748 8148 29200
rect 7868 27692 8148 27748
rect 6076 26852 6356 26908
rect 6748 26852 7028 26908
rect 7420 26852 7700 26908
rect 5852 26180 5908 26190
rect 5404 26178 5908 26180
rect 5404 26126 5854 26178
rect 5906 26126 5908 26178
rect 5404 26124 5908 26126
rect 5852 26114 5908 26124
rect 6076 25620 6132 25630
rect 6076 25526 6132 25564
rect 6300 25508 6356 26852
rect 6860 26290 6916 26302
rect 6860 26238 6862 26290
rect 6914 26238 6916 26290
rect 4956 25340 5236 25396
rect 6188 25506 6356 25508
rect 6188 25454 6302 25506
rect 6354 25454 6356 25506
rect 6188 25452 6356 25454
rect 4620 25284 4676 25294
rect 4620 25190 4676 25228
rect 4732 24948 4788 24958
rect 4396 24946 4788 24948
rect 4396 24894 4734 24946
rect 4786 24894 4788 24946
rect 4396 24892 4788 24894
rect 4732 24882 4788 24892
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 24658 1876 24670
rect 2044 24834 2100 24846
rect 2044 24782 2046 24834
rect 2098 24782 2100 24834
rect 2044 24164 2100 24782
rect 2380 24834 2436 24846
rect 2380 24782 2382 24834
rect 2434 24782 2436 24834
rect 2380 24276 2436 24782
rect 2380 24210 2436 24220
rect 3724 24722 3780 24734
rect 3724 24670 3726 24722
rect 3778 24670 3780 24722
rect 2044 24098 2100 24108
rect 1708 23826 1764 23838
rect 1708 23774 1710 23826
rect 1762 23774 1764 23826
rect 1708 23604 1764 23774
rect 2044 23828 2100 23838
rect 2044 23734 2100 23772
rect 3724 23828 3780 24670
rect 4614 24332 4878 24342
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4614 24266 4878 24276
rect 3724 23762 3780 23772
rect 1708 23538 1764 23548
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 4956 23268 5012 25340
rect 6076 24948 6132 24958
rect 6188 24948 6244 25452
rect 6300 25442 6356 25452
rect 6636 25508 6692 25518
rect 6636 25394 6692 25452
rect 6636 25342 6638 25394
rect 6690 25342 6692 25394
rect 6636 25330 6692 25342
rect 6076 24946 6244 24948
rect 6076 24894 6078 24946
rect 6130 24894 6244 24946
rect 6076 24892 6244 24894
rect 6076 24882 6132 24892
rect 6860 23828 6916 26238
rect 6972 25620 7028 26852
rect 6972 25506 7028 25564
rect 6972 25454 6974 25506
rect 7026 25454 7028 25506
rect 6972 25442 7028 25454
rect 7308 25620 7364 25630
rect 7308 25394 7364 25564
rect 7644 25508 7700 26852
rect 7868 26402 7924 27692
rect 8016 26684 8280 26694
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8016 26618 8280 26628
rect 7868 26350 7870 26402
rect 7922 26350 7924 26402
rect 7868 26338 7924 26350
rect 7308 25342 7310 25394
rect 7362 25342 7364 25394
rect 7308 25330 7364 25342
rect 7420 25506 7700 25508
rect 7420 25454 7646 25506
rect 7698 25454 7700 25506
rect 7420 25452 7700 25454
rect 7420 24946 7476 25452
rect 7644 25442 7700 25452
rect 8540 26290 8596 26302
rect 8540 26238 8542 26290
rect 8594 26238 8596 26290
rect 7980 25396 8036 25406
rect 7980 25302 8036 25340
rect 8428 25284 8484 25294
rect 8016 25116 8280 25126
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8016 25050 8280 25060
rect 7420 24894 7422 24946
rect 7474 24894 7476 24946
rect 7420 24882 7476 24894
rect 8428 23938 8484 25228
rect 8428 23886 8430 23938
rect 8482 23886 8484 23938
rect 8428 23874 8484 23886
rect 6860 23762 6916 23772
rect 8540 23604 8596 26238
rect 8764 25620 8820 29200
rect 9212 25732 9268 25742
rect 8764 25618 9044 25620
rect 8764 25566 8766 25618
rect 8818 25566 9044 25618
rect 8764 25564 9044 25566
rect 8764 25554 8820 25564
rect 8988 25506 9044 25564
rect 8988 25454 8990 25506
rect 9042 25454 9044 25506
rect 8988 25442 9044 25454
rect 8876 24836 8932 24846
rect 8652 24780 8876 24836
rect 8652 23826 8708 24780
rect 8876 24770 8932 24780
rect 9212 23938 9268 25676
rect 9324 25284 9380 25294
rect 9324 25190 9380 25228
rect 9436 24948 9492 29200
rect 10108 27300 10164 29200
rect 10108 27244 10612 27300
rect 9436 24882 9492 24892
rect 9548 26292 9604 26302
rect 9212 23886 9214 23938
rect 9266 23886 9268 23938
rect 9212 23874 9268 23886
rect 8652 23774 8654 23826
rect 8706 23774 8708 23826
rect 8652 23762 8708 23774
rect 8988 23714 9044 23726
rect 8988 23662 8990 23714
rect 9042 23662 9044 23714
rect 8988 23604 9044 23662
rect 8016 23548 8280 23558
rect 8540 23548 9044 23604
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8016 23482 8280 23492
rect 9548 23378 9604 26236
rect 9996 26292 10052 26302
rect 9996 26290 10388 26292
rect 9996 26238 9998 26290
rect 10050 26238 10388 26290
rect 9996 26236 10388 26238
rect 9996 26226 10052 26236
rect 9772 25508 9828 25518
rect 9660 24836 9716 24874
rect 9660 24770 9716 24780
rect 9660 24164 9716 24174
rect 9660 23938 9716 24108
rect 9660 23886 9662 23938
rect 9714 23886 9716 23938
rect 9660 23874 9716 23886
rect 9548 23326 9550 23378
rect 9602 23326 9604 23378
rect 9548 23314 9604 23326
rect 4956 23202 5012 23212
rect 9772 23154 9828 25452
rect 9996 25508 10052 25518
rect 9996 23826 10052 25452
rect 9996 23774 9998 23826
rect 10050 23774 10052 23826
rect 9996 23762 10052 23774
rect 10332 23826 10388 26236
rect 10556 25730 10612 27244
rect 10780 26908 10836 29200
rect 10668 26852 10836 26908
rect 10668 26402 10724 26852
rect 10668 26350 10670 26402
rect 10722 26350 10724 26402
rect 10668 26338 10724 26350
rect 11340 26292 11396 26302
rect 11228 26290 11396 26292
rect 11228 26238 11342 26290
rect 11394 26238 11396 26290
rect 11228 26236 11396 26238
rect 10556 25678 10558 25730
rect 10610 25678 10612 25730
rect 10556 25666 10612 25678
rect 10668 26180 10724 26190
rect 10444 24948 10500 24958
rect 10444 24854 10500 24892
rect 10668 23938 10724 26124
rect 10668 23886 10670 23938
rect 10722 23886 10724 23938
rect 10668 23874 10724 23886
rect 10780 25620 10836 25630
rect 10332 23774 10334 23826
rect 10386 23774 10388 23826
rect 10332 23762 10388 23774
rect 10556 23492 10612 23502
rect 10556 23378 10612 23436
rect 10556 23326 10558 23378
rect 10610 23326 10612 23378
rect 10556 23314 10612 23326
rect 10220 23268 10276 23278
rect 10220 23174 10276 23212
rect 9772 23102 9774 23154
rect 9826 23102 9828 23154
rect 9772 23090 9828 23102
rect 10780 23156 10836 25564
rect 11004 25060 11060 25070
rect 10892 24500 10948 24510
rect 10892 23378 10948 24444
rect 11004 23938 11060 25004
rect 11004 23886 11006 23938
rect 11058 23886 11060 23938
rect 11004 23874 11060 23886
rect 11228 23828 11284 26236
rect 11340 26226 11396 26236
rect 11452 26068 11508 29200
rect 12124 26908 12180 29200
rect 12124 26852 12292 26908
rect 12236 26402 12292 26852
rect 12236 26350 12238 26402
rect 12290 26350 12292 26402
rect 12236 26338 12292 26350
rect 11452 26002 11508 26012
rect 12124 26068 12180 26078
rect 11418 25900 11682 25910
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11418 25834 11682 25844
rect 12124 25618 12180 26012
rect 12796 25732 12852 29200
rect 13468 26850 13524 29200
rect 14140 27076 14196 29200
rect 14140 27020 14644 27076
rect 13468 26798 13470 26850
rect 13522 26798 13524 26850
rect 13468 26786 13524 26798
rect 14140 26850 14196 26862
rect 14140 26798 14142 26850
rect 14194 26798 14196 26850
rect 13692 26292 13748 26302
rect 12796 25666 12852 25676
rect 13580 26290 13748 26292
rect 13580 26238 13694 26290
rect 13746 26238 13748 26290
rect 13580 26236 13748 26238
rect 12124 25566 12126 25618
rect 12178 25566 12180 25618
rect 12124 25554 12180 25566
rect 11788 25508 11844 25518
rect 11788 25414 11844 25452
rect 11900 25396 11956 25406
rect 11340 25282 11396 25294
rect 11340 25230 11342 25282
rect 11394 25230 11396 25282
rect 11340 24500 11396 25230
rect 11340 24434 11396 24444
rect 11418 24332 11682 24342
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11418 24266 11682 24276
rect 11900 23938 11956 25340
rect 13468 25282 13524 25294
rect 13468 25230 13470 25282
rect 13522 25230 13524 25282
rect 13468 24052 13524 25230
rect 11900 23886 11902 23938
rect 11954 23886 11956 23938
rect 11900 23874 11956 23886
rect 13356 23996 13524 24052
rect 11340 23828 11396 23838
rect 11228 23826 11396 23828
rect 11228 23774 11342 23826
rect 11394 23774 11396 23826
rect 11228 23772 11396 23774
rect 11340 23762 11396 23772
rect 11676 23828 11732 23838
rect 11676 23734 11732 23772
rect 13356 23492 13412 23996
rect 13468 23828 13524 23838
rect 13580 23828 13636 26236
rect 13692 26226 13748 26236
rect 14140 26178 14196 26798
rect 14140 26126 14142 26178
rect 14194 26126 14196 26178
rect 14140 26114 14196 26126
rect 13916 25732 13972 25742
rect 13916 25618 13972 25676
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 13916 25554 13972 25566
rect 14364 24836 14420 24846
rect 13804 24834 14420 24836
rect 13804 24782 14366 24834
rect 14418 24782 14420 24834
rect 13804 24780 14420 24782
rect 13804 23938 13860 24780
rect 14364 24770 14420 24780
rect 14588 24724 14644 27020
rect 14812 26908 14868 29200
rect 14700 26852 14868 26908
rect 14700 25620 14756 26852
rect 14820 26684 15084 26694
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 14820 26618 15084 26628
rect 15484 26628 15540 29200
rect 15484 26572 15988 26628
rect 15484 26514 15540 26572
rect 15484 26462 15486 26514
rect 15538 26462 15540 26514
rect 15484 26450 15540 26462
rect 15708 26404 15764 26414
rect 15596 26402 15764 26404
rect 15596 26350 15710 26402
rect 15762 26350 15764 26402
rect 15596 26348 15764 26350
rect 14812 25620 14868 25630
rect 14700 25618 15092 25620
rect 14700 25566 14814 25618
rect 14866 25566 15092 25618
rect 14700 25564 15092 25566
rect 14812 25554 14868 25564
rect 15036 25506 15092 25564
rect 15596 25508 15652 26348
rect 15708 26338 15764 26348
rect 15932 26290 15988 26572
rect 16156 26516 16212 29200
rect 16156 26450 16212 26460
rect 15932 26238 15934 26290
rect 15986 26238 15988 26290
rect 15932 26226 15988 26238
rect 15036 25454 15038 25506
rect 15090 25454 15092 25506
rect 15036 25442 15092 25454
rect 15148 25452 15652 25508
rect 15932 25844 15988 25854
rect 14820 25116 15084 25126
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 14820 25050 15084 25060
rect 15148 24948 15204 25452
rect 14476 24722 14644 24724
rect 14476 24670 14590 24722
rect 14642 24670 14644 24722
rect 14476 24668 14644 24670
rect 14140 24612 14196 24622
rect 14476 24612 14532 24668
rect 14588 24658 14644 24668
rect 15036 24892 15204 24948
rect 15260 25284 15316 25294
rect 14140 24610 14532 24612
rect 14140 24558 14142 24610
rect 14194 24558 14532 24610
rect 14140 24556 14532 24558
rect 14140 24546 14196 24556
rect 13804 23886 13806 23938
rect 13858 23886 13860 23938
rect 13804 23874 13860 23886
rect 15036 23938 15092 24892
rect 15036 23886 15038 23938
rect 15090 23886 15092 23938
rect 15036 23874 15092 23886
rect 13468 23826 13636 23828
rect 13468 23774 13470 23826
rect 13522 23774 13636 23826
rect 13468 23772 13636 23774
rect 15260 23826 15316 25228
rect 15372 25284 15428 25294
rect 15372 25282 15652 25284
rect 15372 25230 15374 25282
rect 15426 25230 15652 25282
rect 15372 25228 15652 25230
rect 15372 25218 15428 25228
rect 15596 23938 15652 25228
rect 15596 23886 15598 23938
rect 15650 23886 15652 23938
rect 15596 23874 15652 23886
rect 15260 23774 15262 23826
rect 15314 23774 15316 23826
rect 13468 23762 13524 23772
rect 15260 23762 15316 23774
rect 15932 23826 15988 25788
rect 16828 25620 16884 29200
rect 17500 26852 17556 29200
rect 17500 26786 17556 26796
rect 18172 26628 18228 29200
rect 18844 26850 18900 29200
rect 18844 26798 18846 26850
rect 18898 26798 18900 26850
rect 18844 26786 18900 26798
rect 18956 26852 19012 26862
rect 18172 26562 18228 26572
rect 18844 26628 18900 26638
rect 17388 26516 17444 26526
rect 16940 26290 16996 26302
rect 16940 26238 16942 26290
rect 16994 26238 16996 26290
rect 16940 25844 16996 26238
rect 17388 26178 17444 26460
rect 17388 26126 17390 26178
rect 17442 26126 17444 26178
rect 17388 26114 17444 26126
rect 18620 26290 18676 26302
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18222 25900 18486 25910
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18222 25834 18486 25844
rect 16940 25778 16996 25788
rect 16828 25618 17332 25620
rect 16828 25566 16830 25618
rect 16882 25566 17332 25618
rect 16828 25564 17332 25566
rect 16828 25554 16884 25564
rect 17276 25506 17332 25564
rect 17276 25454 17278 25506
rect 17330 25454 17332 25506
rect 17276 25442 17332 25454
rect 18508 25508 18564 25518
rect 18508 25414 18564 25452
rect 16828 25396 16884 25406
rect 16492 25284 16548 25294
rect 16492 23938 16548 25228
rect 16492 23886 16494 23938
rect 16546 23886 16548 23938
rect 16492 23874 16548 23886
rect 15932 23774 15934 23826
rect 15986 23774 15988 23826
rect 15932 23762 15988 23774
rect 16828 23826 16884 25340
rect 18620 25396 18676 26238
rect 18844 25618 18900 26572
rect 18956 26178 19012 26796
rect 18956 26126 18958 26178
rect 19010 26126 19012 26178
rect 18956 26114 19012 26126
rect 18844 25566 18846 25618
rect 18898 25566 18900 25618
rect 18844 25554 18900 25566
rect 19516 25620 19572 29200
rect 20076 26850 20132 26862
rect 20076 26798 20078 26850
rect 20130 26798 20132 26850
rect 20076 26514 20132 26798
rect 20188 26852 20244 29200
rect 20300 26852 20356 26862
rect 20188 26850 20356 26852
rect 20188 26798 20302 26850
rect 20354 26798 20356 26850
rect 20188 26796 20356 26798
rect 20300 26786 20356 26796
rect 20076 26462 20078 26514
rect 20130 26462 20132 26514
rect 20076 26450 20132 26462
rect 20748 26292 20804 26302
rect 20132 26290 20804 26292
rect 20132 26238 20750 26290
rect 20802 26238 20804 26290
rect 20132 26236 20804 26238
rect 20132 26180 20188 26236
rect 20748 26226 20804 26236
rect 20076 26124 20188 26180
rect 19628 25620 19684 25630
rect 19516 25564 19628 25620
rect 19628 25526 19684 25564
rect 18620 25330 18676 25340
rect 17052 25284 17108 25294
rect 19964 25284 20020 25294
rect 17052 25190 17108 25228
rect 19852 25282 20020 25284
rect 19852 25230 19966 25282
rect 20018 25230 20020 25282
rect 19852 25228 20020 25230
rect 18222 24332 18486 24342
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18222 24266 18486 24276
rect 19852 23938 19908 25228
rect 19964 25218 20020 25228
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23874 19908 23886
rect 16828 23774 16830 23826
rect 16882 23774 16884 23826
rect 16828 23762 16884 23774
rect 20076 23826 20132 26124
rect 20188 25620 20244 25630
rect 20188 25506 20244 25564
rect 20860 25620 20916 29200
rect 21196 26850 21252 26862
rect 21196 26798 21198 26850
rect 21250 26798 21252 26850
rect 21196 26178 21252 26798
rect 21532 26852 21588 29200
rect 21532 26786 21588 26796
rect 22204 26850 22260 29200
rect 22876 27188 22932 29200
rect 22876 27132 23044 27188
rect 22204 26798 22206 26850
rect 22258 26798 22260 26850
rect 22204 26786 22260 26798
rect 22764 26852 22820 26862
rect 21624 26684 21888 26694
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21624 26618 21888 26628
rect 22428 26292 22484 26302
rect 22428 26290 22596 26292
rect 22428 26238 22430 26290
rect 22482 26238 22596 26290
rect 22428 26236 22596 26238
rect 22428 26226 22484 26236
rect 21196 26126 21198 26178
rect 21250 26126 21252 26178
rect 21196 26114 21252 26126
rect 20860 25618 21364 25620
rect 20860 25566 20862 25618
rect 20914 25566 21364 25618
rect 20860 25564 21364 25566
rect 20860 25554 20916 25564
rect 20188 25454 20190 25506
rect 20242 25454 20244 25506
rect 20188 25442 20244 25454
rect 21308 25506 21364 25564
rect 21308 25454 21310 25506
rect 21362 25454 21364 25506
rect 21308 25442 21364 25454
rect 20748 25396 20804 25406
rect 20524 25284 20580 25294
rect 20524 23938 20580 25228
rect 20524 23886 20526 23938
rect 20578 23886 20580 23938
rect 20524 23874 20580 23886
rect 20076 23774 20078 23826
rect 20130 23774 20132 23826
rect 20076 23762 20132 23774
rect 20748 23826 20804 25340
rect 21644 25284 21700 25294
rect 22428 25284 22484 25294
rect 21420 25282 21700 25284
rect 21420 25230 21646 25282
rect 21698 25230 21700 25282
rect 21420 25228 21700 25230
rect 20748 23774 20750 23826
rect 20802 23774 20804 23826
rect 20748 23762 20804 23774
rect 20860 24724 20916 24734
rect 14820 23548 15084 23558
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 14820 23482 15084 23492
rect 13356 23426 13412 23436
rect 10892 23326 10894 23378
rect 10946 23326 10948 23378
rect 10892 23314 10948 23326
rect 20860 23378 20916 24668
rect 21420 23938 21476 25228
rect 21644 25218 21700 25228
rect 21980 25282 22484 25284
rect 21980 25230 22430 25282
rect 22482 25230 22484 25282
rect 21980 25228 22484 25230
rect 21624 25116 21888 25126
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21624 25050 21888 25060
rect 21980 24948 22036 25228
rect 22428 25218 22484 25228
rect 21420 23886 21422 23938
rect 21474 23886 21476 23938
rect 21420 23874 21476 23886
rect 21644 24892 22036 24948
rect 21644 23826 21700 24892
rect 22540 24724 22596 26236
rect 22764 26178 22820 26796
rect 22764 26126 22766 26178
rect 22818 26126 22820 26178
rect 22764 26114 22820 26126
rect 22876 26850 22932 26862
rect 22876 26798 22878 26850
rect 22930 26798 22932 26850
rect 22876 25618 22932 26798
rect 22988 26852 23044 27132
rect 22988 26786 23044 26796
rect 22876 25566 22878 25618
rect 22930 25566 22932 25618
rect 22876 25554 22932 25566
rect 23548 25508 23604 29200
rect 24220 26850 24276 29200
rect 24220 26798 24222 26850
rect 24274 26798 24276 26850
rect 24108 26516 24164 26526
rect 24220 26516 24276 26798
rect 24108 26514 24276 26516
rect 24108 26462 24110 26514
rect 24162 26462 24276 26514
rect 24108 26460 24276 26462
rect 24108 26450 24164 26460
rect 23660 25508 23716 25518
rect 24220 25508 24276 25518
rect 23548 25506 24276 25508
rect 23548 25454 23662 25506
rect 23714 25454 24222 25506
rect 24274 25454 24276 25506
rect 23548 25452 24276 25454
rect 23660 25442 23716 25452
rect 24220 25442 24276 25452
rect 23996 25284 24052 25294
rect 23996 25190 24052 25228
rect 22540 24658 22596 24668
rect 23100 25172 23156 25182
rect 23100 24722 23156 25116
rect 23660 25172 23716 25182
rect 23100 24670 23102 24722
rect 23154 24670 23156 24722
rect 23100 24658 23156 24670
rect 23324 24834 23380 24846
rect 23324 24782 23326 24834
rect 23378 24782 23380 24834
rect 22764 24612 22820 24622
rect 22764 24518 22820 24556
rect 23324 23940 23380 24782
rect 23660 24050 23716 25116
rect 24444 25172 24500 29596
rect 24864 29200 24976 30000
rect 24780 26850 24836 26862
rect 24780 26798 24782 26850
rect 24834 26798 24836 26850
rect 24556 26290 24612 26302
rect 24556 26238 24558 26290
rect 24610 26238 24612 26290
rect 24556 25396 24612 26238
rect 24780 25508 24836 26798
rect 24892 26516 24948 29200
rect 27804 28980 27860 28990
rect 25116 28308 25172 28318
rect 24892 26450 24948 26460
rect 25004 26852 25060 26862
rect 25004 26178 25060 26796
rect 25004 26126 25006 26178
rect 25058 26126 25060 26178
rect 25004 26114 25060 26126
rect 25116 26068 25172 28252
rect 27468 27636 27524 27646
rect 25900 26964 25956 26974
rect 25116 26012 25508 26068
rect 25026 25900 25290 25910
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25026 25834 25290 25844
rect 24892 25508 24948 25518
rect 24780 25506 24948 25508
rect 24780 25454 24894 25506
rect 24946 25454 24948 25506
rect 24780 25452 24948 25454
rect 24892 25442 24948 25452
rect 24556 25330 24612 25340
rect 24668 25284 24724 25294
rect 25340 25284 25396 25294
rect 24668 25190 24724 25228
rect 25116 25282 25396 25284
rect 25116 25230 25342 25282
rect 25394 25230 25396 25282
rect 25116 25228 25396 25230
rect 24444 25106 24500 25116
rect 23772 24948 23828 24958
rect 23772 24722 23828 24892
rect 23996 24836 24052 24846
rect 24332 24836 24388 24846
rect 23996 24742 24052 24780
rect 24108 24834 24388 24836
rect 24108 24782 24334 24834
rect 24386 24782 24388 24834
rect 24108 24780 24388 24782
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23772 24658 23828 24670
rect 23660 23998 23662 24050
rect 23714 23998 23716 24050
rect 23660 23986 23716 23998
rect 23324 23874 23380 23884
rect 23996 23940 24052 23950
rect 24108 23940 24164 24780
rect 24332 24770 24388 24780
rect 24668 24722 24724 24734
rect 24668 24670 24670 24722
rect 24722 24670 24724 24722
rect 24668 24612 24724 24670
rect 23996 23938 24164 23940
rect 23996 23886 23998 23938
rect 24050 23886 24164 23938
rect 23996 23884 24164 23886
rect 24220 24164 24276 24174
rect 23996 23874 24052 23884
rect 21644 23774 21646 23826
rect 21698 23774 21700 23826
rect 21644 23762 21700 23774
rect 24220 23826 24276 24108
rect 24220 23774 24222 23826
rect 24274 23774 24276 23826
rect 24220 23762 24276 23774
rect 24556 23826 24612 23838
rect 24556 23774 24558 23826
rect 24610 23774 24612 23826
rect 21624 23548 21888 23558
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21624 23482 21888 23492
rect 20860 23326 20862 23378
rect 20914 23326 20916 23378
rect 20860 23314 20916 23326
rect 20636 23268 20692 23278
rect 11116 23156 11172 23166
rect 10780 23154 11172 23156
rect 10780 23102 11118 23154
rect 11170 23102 11172 23154
rect 10780 23100 11172 23102
rect 11116 23090 11172 23100
rect 20636 23154 20692 23212
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20636 23090 20692 23102
rect 24444 23154 24500 23166
rect 24444 23102 24446 23154
rect 24498 23102 24500 23154
rect 4614 22764 4878 22774
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4614 22698 4878 22708
rect 11418 22764 11682 22774
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11418 22698 11682 22708
rect 18222 22764 18486 22774
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18222 22698 18486 22708
rect 8016 21980 8280 21990
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8016 21914 8280 21924
rect 14820 21980 15084 21990
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 14820 21914 15084 21924
rect 21624 21980 21888 21990
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21624 21914 21888 21924
rect 13020 21700 13076 21710
rect 12348 21476 12404 21486
rect 4614 21196 4878 21206
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4614 21130 4878 21140
rect 11418 21196 11682 21206
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11418 21130 11682 21140
rect 8016 20412 8280 20422
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8016 20346 8280 20356
rect 9884 20018 9940 20030
rect 9884 19966 9886 20018
rect 9938 19966 9940 20018
rect 8540 19796 8596 19806
rect 4614 19628 4878 19638
rect 4284 19572 4340 19582
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4614 19562 4878 19572
rect 3948 17442 4004 17454
rect 3948 17390 3950 17442
rect 4002 17390 4004 17442
rect 2268 17106 2324 17118
rect 2268 17054 2270 17106
rect 2322 17054 2324 17106
rect 1596 16660 1652 16670
rect 1596 16566 1652 16604
rect 2044 15202 2100 15214
rect 2044 15150 2046 15202
rect 2098 15150 2100 15202
rect 2044 14530 2100 15150
rect 2268 14754 2324 17054
rect 3612 16884 3668 16894
rect 2716 16660 2772 16670
rect 2716 15986 2772 16604
rect 2716 15934 2718 15986
rect 2770 15934 2772 15986
rect 2716 15922 2772 15934
rect 2716 15314 2772 15326
rect 2716 15262 2718 15314
rect 2770 15262 2772 15314
rect 2268 14702 2270 14754
rect 2322 14702 2324 14754
rect 2268 14690 2324 14702
rect 2604 15202 2660 15214
rect 2604 15150 2606 15202
rect 2658 15150 2660 15202
rect 2044 14478 2046 14530
rect 2098 14478 2100 14530
rect 2044 14308 2100 14478
rect 2044 14242 2100 14252
rect 2604 13970 2660 15150
rect 2716 14308 2772 15262
rect 3612 15314 3668 16828
rect 3948 16660 4004 17390
rect 3948 16594 4004 16604
rect 3612 15262 3614 15314
rect 3666 15262 3668 15314
rect 3612 15250 3668 15262
rect 3948 16210 4004 16222
rect 3948 16158 3950 16210
rect 4002 16158 4004 16210
rect 3948 15314 4004 16158
rect 3948 15262 3950 15314
rect 4002 15262 4004 15314
rect 3948 15250 4004 15262
rect 4060 14642 4116 14654
rect 4060 14590 4062 14642
rect 4114 14590 4116 14642
rect 3052 14420 3108 14430
rect 3052 14326 3108 14364
rect 2716 14242 2772 14252
rect 3388 14308 3444 14318
rect 2604 13918 2606 13970
rect 2658 13918 2660 13970
rect 2604 13906 2660 13918
rect 2044 13522 2100 13534
rect 2044 13470 2046 13522
rect 2098 13470 2100 13522
rect 2044 12852 2100 13470
rect 2716 12852 2772 12862
rect 2044 12850 2772 12852
rect 2044 12798 2718 12850
rect 2770 12798 2772 12850
rect 2044 12796 2772 12798
rect 2716 12786 2772 12796
rect 2380 12290 2436 12302
rect 2380 12238 2382 12290
rect 2434 12238 2436 12290
rect 1596 11954 1652 11966
rect 1596 11902 1598 11954
rect 1650 11902 1652 11954
rect 1596 11284 1652 11902
rect 1596 11218 1652 11228
rect 1820 11394 1876 11406
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 10836 1876 11342
rect 1820 10742 1876 10780
rect 2044 11170 2100 11182
rect 2044 11118 2046 11170
rect 2098 11118 2100 11170
rect 2044 8428 2100 11118
rect 2380 10388 2436 12238
rect 3388 11396 3444 14252
rect 4060 13748 4116 14590
rect 4060 13682 4116 13692
rect 4060 13074 4116 13086
rect 4060 13022 4062 13074
rect 4114 13022 4116 13074
rect 4060 12740 4116 13022
rect 4284 12964 4340 19516
rect 6076 19348 6132 19358
rect 5516 18450 5572 18462
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 4614 18060 4878 18070
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4614 17994 4878 18004
rect 4508 17666 4564 17678
rect 4508 17614 4510 17666
rect 4562 17614 4564 17666
rect 4508 17444 4564 17614
rect 5516 17668 5572 18398
rect 6076 18450 6132 19292
rect 7644 19348 7700 19358
rect 7644 19254 7700 19292
rect 8016 18844 8280 18854
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8016 18778 8280 18788
rect 8540 18674 8596 19740
rect 9548 19796 9604 19806
rect 9548 19702 9604 19740
rect 9548 19234 9604 19246
rect 9548 19182 9550 19234
rect 9602 19182 9604 19234
rect 8540 18622 8542 18674
rect 8594 18622 8596 18674
rect 8540 18610 8596 18622
rect 8988 19122 9044 19134
rect 8988 19070 8990 19122
rect 9042 19070 9044 19122
rect 6076 18398 6078 18450
rect 6130 18398 6132 18450
rect 6076 18386 6132 18398
rect 4956 17444 5012 17454
rect 4508 17388 4956 17444
rect 4620 16884 4676 16894
rect 4284 12898 4340 12908
rect 4396 16882 4676 16884
rect 4396 16830 4622 16882
rect 4674 16830 4676 16882
rect 4396 16828 4676 16830
rect 4396 12740 4452 16828
rect 4620 16818 4676 16828
rect 4614 16492 4878 16502
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4614 16426 4878 16436
rect 4614 14924 4878 14934
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4614 14858 4878 14868
rect 4508 14308 4564 14318
rect 4956 14308 5012 17388
rect 5068 16884 5124 16894
rect 5068 16790 5124 16828
rect 5516 16884 5572 17612
rect 5628 17666 5684 17678
rect 5628 17614 5630 17666
rect 5682 17614 5684 17666
rect 5628 17444 5684 17614
rect 7532 17668 7588 17678
rect 7532 17574 7588 17612
rect 8204 17666 8260 17678
rect 8204 17614 8206 17666
rect 8258 17614 8260 17666
rect 5628 17378 5684 17388
rect 6188 17444 6244 17454
rect 6636 17444 6692 17454
rect 6188 17442 6356 17444
rect 6188 17390 6190 17442
rect 6242 17390 6356 17442
rect 6188 17388 6356 17390
rect 6188 17378 6244 17388
rect 5516 16790 5572 16828
rect 6076 16882 6132 16894
rect 6076 16830 6078 16882
rect 6130 16830 6132 16882
rect 5852 16660 5908 16670
rect 5852 15148 5908 16604
rect 6076 16212 6132 16830
rect 6076 16146 6132 16156
rect 6300 15538 6356 17388
rect 8204 17444 8260 17614
rect 8204 17388 8484 17444
rect 6636 17350 6692 17388
rect 8016 17276 8280 17286
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8016 17210 8280 17220
rect 8316 16994 8372 17006
rect 8316 16942 8318 16994
rect 8370 16942 8372 16994
rect 6972 16212 7028 16222
rect 6972 16118 7028 16156
rect 8316 16100 8372 16942
rect 8428 16772 8484 17388
rect 8988 17108 9044 19070
rect 9548 18452 9604 19182
rect 9100 18228 9156 18238
rect 9100 18226 9268 18228
rect 9100 18174 9102 18226
rect 9154 18174 9268 18226
rect 9100 18172 9268 18174
rect 9100 18162 9156 18172
rect 9100 17108 9156 17118
rect 8988 17106 9156 17108
rect 8988 17054 9102 17106
rect 9154 17054 9156 17106
rect 8988 17052 9156 17054
rect 9100 17042 9156 17052
rect 8428 16706 8484 16716
rect 8316 16044 8484 16100
rect 7980 15988 8036 15998
rect 6300 15486 6302 15538
rect 6354 15486 6356 15538
rect 6300 15474 6356 15486
rect 7084 15986 8036 15988
rect 7084 15934 7982 15986
rect 8034 15934 8036 15986
rect 7084 15932 8036 15934
rect 7084 15538 7140 15932
rect 7980 15922 8036 15932
rect 8016 15708 8280 15718
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8016 15642 8280 15652
rect 7084 15486 7086 15538
rect 7138 15486 7140 15538
rect 7084 15474 7140 15486
rect 8428 15538 8484 16044
rect 9212 15988 9268 18172
rect 9212 15922 9268 15932
rect 9548 17668 9604 18396
rect 9884 18450 9940 19966
rect 11900 20018 11956 20030
rect 11900 19966 11902 20018
rect 11954 19966 11956 20018
rect 11418 19628 11682 19638
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11418 19562 11682 19572
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9884 17668 9940 18398
rect 9996 19234 10052 19246
rect 9996 19182 9998 19234
rect 10050 19182 10052 19234
rect 9996 18340 10052 19182
rect 9996 18274 10052 18284
rect 11228 18564 11284 18574
rect 10220 18228 10276 18238
rect 10220 18226 10500 18228
rect 10220 18174 10222 18226
rect 10274 18174 10500 18226
rect 10220 18172 10500 18174
rect 10220 18162 10276 18172
rect 9996 17668 10052 17678
rect 9884 17612 9996 17668
rect 9548 16996 9604 17612
rect 9996 17602 10052 17612
rect 10444 17554 10500 18172
rect 11228 17890 11284 18508
rect 11900 18452 11956 19966
rect 12348 20018 12404 21420
rect 12348 19966 12350 20018
rect 12402 19966 12404 20018
rect 12348 19954 12404 19966
rect 13020 19458 13076 21644
rect 14812 21700 14868 21710
rect 14812 21606 14868 21644
rect 24444 21700 24500 23102
rect 24444 21634 24500 21644
rect 13804 21476 13860 21486
rect 13804 21382 13860 21420
rect 18222 21196 18486 21206
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18222 21130 18486 21140
rect 16268 20914 16324 20926
rect 16268 20862 16270 20914
rect 16322 20862 16324 20914
rect 15372 20692 15428 20702
rect 14820 20412 15084 20422
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 14820 20346 15084 20356
rect 14924 20244 14980 20254
rect 14588 20132 14644 20142
rect 13020 19406 13022 19458
rect 13074 19406 13076 19458
rect 13020 19394 13076 19406
rect 14028 20130 14644 20132
rect 14028 20078 14590 20130
rect 14642 20078 14644 20130
rect 14028 20076 14644 20078
rect 14028 19458 14084 20076
rect 14588 20066 14644 20076
rect 14028 19406 14030 19458
rect 14082 19406 14084 19458
rect 14028 19394 14084 19406
rect 13468 19234 13524 19246
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 12236 19012 12292 19022
rect 11900 18386 11956 18396
rect 12012 19010 12292 19012
rect 12012 18958 12238 19010
rect 12290 18958 12292 19010
rect 12012 18956 12292 18958
rect 11564 18340 11620 18350
rect 11564 18246 11620 18284
rect 11418 18060 11682 18070
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11418 17994 11682 18004
rect 11228 17838 11230 17890
rect 11282 17838 11284 17890
rect 11228 17826 11284 17838
rect 12012 17890 12068 18956
rect 12236 18946 12292 18956
rect 12572 18564 12628 18574
rect 12572 18470 12628 18508
rect 12012 17838 12014 17890
rect 12066 17838 12068 17890
rect 12012 17826 12068 17838
rect 12460 18452 12516 18462
rect 10444 17502 10446 17554
rect 10498 17502 10500 17554
rect 10444 17490 10500 17502
rect 11676 17668 11732 17678
rect 9772 16996 9828 17006
rect 9548 16994 9828 16996
rect 9548 16942 9774 16994
rect 9826 16942 9828 16994
rect 9548 16940 9828 16942
rect 8428 15486 8430 15538
rect 8482 15486 8484 15538
rect 8428 15474 8484 15486
rect 8988 15316 9044 15326
rect 8988 15222 9044 15260
rect 5852 15092 6132 15148
rect 5516 14420 5572 14430
rect 5516 14326 5572 14364
rect 4564 14252 5012 14308
rect 6076 14306 6132 15092
rect 8652 14644 8708 14654
rect 8652 14530 8708 14588
rect 8652 14478 8654 14530
rect 8706 14478 8708 14530
rect 8652 14466 8708 14478
rect 9212 14532 9268 14542
rect 9548 14532 9604 16940
rect 9772 16930 9828 16940
rect 9772 16772 9828 16782
rect 11676 16772 11732 17612
rect 11676 16716 11844 16772
rect 9772 16210 9828 16716
rect 11418 16492 11682 16502
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11418 16426 11682 16436
rect 9772 16158 9774 16210
rect 9826 16158 9828 16210
rect 9772 16146 9828 16158
rect 10780 15988 10836 15998
rect 10780 15894 10836 15932
rect 11452 15316 11508 15326
rect 11452 15148 11508 15260
rect 11788 15148 11844 16716
rect 12012 15988 12068 15998
rect 12012 15538 12068 15932
rect 12012 15486 12014 15538
rect 12066 15486 12068 15538
rect 12012 15474 12068 15486
rect 11228 15090 11284 15102
rect 11452 15092 11844 15148
rect 12460 15148 12516 18396
rect 13244 18452 13300 18462
rect 13244 18358 13300 18396
rect 13468 17668 13524 19182
rect 14252 19234 14308 19246
rect 14252 19182 14254 19234
rect 14306 19182 14308 19234
rect 14252 18564 14308 19182
rect 14924 19234 14980 20188
rect 15372 20130 15428 20636
rect 16268 20244 16324 20862
rect 22876 20916 22932 20926
rect 17276 20692 17332 20702
rect 17276 20598 17332 20636
rect 21624 20412 21888 20422
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21624 20346 21888 20356
rect 16268 20178 16324 20188
rect 20524 20242 20580 20254
rect 20524 20190 20526 20242
rect 20578 20190 20580 20242
rect 20524 20188 20580 20190
rect 20524 20132 21364 20188
rect 15372 20078 15374 20130
rect 15426 20078 15428 20130
rect 15372 20066 15428 20078
rect 15820 20020 15876 20030
rect 14924 19182 14926 19234
rect 14978 19182 14980 19234
rect 14924 19170 14980 19182
rect 15708 20018 15876 20020
rect 15708 19966 15822 20018
rect 15874 19966 15876 20018
rect 15708 19964 15876 19966
rect 14820 18844 15084 18854
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 14820 18778 15084 18788
rect 14252 18498 14308 18508
rect 13916 18450 13972 18462
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13692 17668 13748 17678
rect 13524 17666 13748 17668
rect 13524 17614 13694 17666
rect 13746 17614 13748 17666
rect 13524 17612 13748 17614
rect 13468 17602 13524 17612
rect 13692 17602 13748 17612
rect 12796 17444 12852 17454
rect 12796 15538 12852 17388
rect 13804 17444 13860 17454
rect 13804 17350 13860 17388
rect 13916 17332 13972 18398
rect 15708 17668 15764 19964
rect 15820 19954 15876 19964
rect 17612 20018 17668 20030
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 16380 19794 16436 19806
rect 16380 19742 16382 19794
rect 16434 19742 16436 19794
rect 16380 19124 16436 19742
rect 16380 19058 16436 19068
rect 17164 19124 17220 19134
rect 17164 19030 17220 19068
rect 16156 18564 16212 18574
rect 15820 18562 16212 18564
rect 15820 18510 16158 18562
rect 16210 18510 16212 18562
rect 15820 18508 16212 18510
rect 15820 17890 15876 18508
rect 16156 18498 16212 18508
rect 16940 18564 16996 18574
rect 16940 18450 16996 18508
rect 16940 18398 16942 18450
rect 16994 18398 16996 18450
rect 16940 18386 16996 18398
rect 16940 18228 16996 18238
rect 15820 17838 15822 17890
rect 15874 17838 15876 17890
rect 15820 17826 15876 17838
rect 16828 18172 16940 18228
rect 16156 17668 16212 17678
rect 15708 17574 15764 17612
rect 16044 17666 16212 17668
rect 16044 17614 16158 17666
rect 16210 17614 16212 17666
rect 16044 17612 16212 17614
rect 13916 17276 14756 17332
rect 14588 16882 14644 16894
rect 14588 16830 14590 16882
rect 14642 16830 14644 16882
rect 13580 15988 13636 15998
rect 13580 15894 13636 15932
rect 12796 15486 12798 15538
rect 12850 15486 12852 15538
rect 12796 15474 12852 15486
rect 12460 15092 12628 15148
rect 11228 15038 11230 15090
rect 11282 15038 11284 15090
rect 9212 14530 9604 14532
rect 9212 14478 9214 14530
rect 9266 14478 9550 14530
rect 9602 14478 9604 14530
rect 9212 14476 9604 14478
rect 9212 14466 9268 14476
rect 9548 14466 9604 14476
rect 9884 14530 9940 14542
rect 9884 14478 9886 14530
rect 9938 14478 9940 14530
rect 6076 14254 6078 14306
rect 6130 14254 6132 14306
rect 4508 14214 4564 14252
rect 6076 14242 6132 14254
rect 8016 14140 8280 14150
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8016 14074 8280 14084
rect 7980 13972 8036 13982
rect 6972 13858 7028 13870
rect 6972 13806 6974 13858
rect 7026 13806 7028 13858
rect 5068 13748 5124 13758
rect 5068 13654 5124 13692
rect 5740 13746 5796 13758
rect 5740 13694 5742 13746
rect 5794 13694 5796 13746
rect 4614 13356 4878 13366
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4614 13290 4878 13300
rect 4060 12684 4452 12740
rect 5404 12404 5460 12414
rect 5628 12404 5684 12414
rect 5404 12402 5628 12404
rect 5404 12350 5406 12402
rect 5458 12350 5628 12402
rect 5404 12348 5628 12350
rect 5404 12338 5460 12348
rect 5628 12338 5684 12348
rect 4620 12180 4676 12190
rect 3948 12178 4676 12180
rect 3948 12126 4622 12178
rect 4674 12126 4676 12178
rect 3948 12124 4676 12126
rect 3836 11508 3892 11518
rect 2716 11284 2772 11294
rect 2716 11190 2772 11228
rect 2380 10322 2436 10332
rect 2716 10612 2772 10622
rect 2716 9042 2772 10556
rect 2940 10612 2996 10622
rect 3276 10612 3332 10622
rect 2940 10610 3332 10612
rect 2940 10558 2942 10610
rect 2994 10558 3278 10610
rect 3330 10558 3332 10610
rect 2940 10556 3332 10558
rect 2940 10546 2996 10556
rect 3276 10500 3332 10556
rect 3276 10434 3332 10444
rect 3388 10500 3444 11340
rect 3388 10434 3444 10444
rect 3500 11506 3892 11508
rect 3500 11454 3838 11506
rect 3890 11454 3892 11506
rect 3500 11452 3892 11454
rect 2716 8990 2718 9042
rect 2770 8990 2772 9042
rect 2044 8372 2436 8428
rect 2044 7474 2100 7486
rect 2044 7422 2046 7474
rect 2098 7422 2100 7474
rect 2044 7252 2100 7422
rect 2380 7474 2436 8372
rect 2380 7422 2382 7474
rect 2434 7422 2436 7474
rect 2380 7410 2436 7422
rect 2716 7252 2772 8990
rect 3388 9044 3444 9054
rect 3500 9044 3556 11452
rect 3836 11442 3892 11452
rect 3388 9042 3556 9044
rect 3388 8990 3390 9042
rect 3442 8990 3556 9042
rect 3388 8988 3556 8990
rect 3724 10498 3780 10510
rect 3724 10446 3726 10498
rect 3778 10446 3780 10498
rect 3388 8978 3444 8988
rect 3724 7812 3780 10446
rect 3836 9940 3892 9950
rect 3948 9940 4004 12124
rect 4620 12114 4676 12124
rect 5292 12178 5348 12190
rect 5292 12126 5294 12178
rect 5346 12126 5348 12178
rect 5292 12068 5348 12126
rect 4614 11788 4878 11798
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4614 11722 4878 11732
rect 4284 10612 4340 10622
rect 4284 10518 4340 10556
rect 4732 10612 4788 10622
rect 5292 10612 5348 12012
rect 5740 12068 5796 13694
rect 6972 13188 7028 13806
rect 7980 13634 8036 13916
rect 9884 13972 9940 14478
rect 9884 13906 9940 13916
rect 7980 13582 7982 13634
rect 8034 13582 8036 13634
rect 7980 13570 8036 13582
rect 10108 13748 10164 13758
rect 10892 13748 10948 13758
rect 10108 13746 10948 13748
rect 10108 13694 10110 13746
rect 10162 13694 10894 13746
rect 10946 13694 10948 13746
rect 10108 13692 10948 13694
rect 9884 13524 9940 13534
rect 6972 13122 7028 13132
rect 9100 13188 9156 13198
rect 9100 13094 9156 13132
rect 7868 13074 7924 13086
rect 7868 13022 7870 13074
rect 7922 13022 7924 13074
rect 6524 12850 6580 12862
rect 6524 12798 6526 12850
rect 6578 12798 6580 12850
rect 6524 12404 6580 12798
rect 6524 12338 6580 12348
rect 5740 12002 5796 12012
rect 6188 12290 6244 12302
rect 6188 12238 6190 12290
rect 6242 12238 6244 12290
rect 6188 10836 6244 12238
rect 7756 12068 7812 12078
rect 6188 10770 6244 10780
rect 6300 11396 6356 11406
rect 4732 10610 5012 10612
rect 4732 10558 4734 10610
rect 4786 10558 5012 10610
rect 4732 10556 5012 10558
rect 4732 10546 4788 10556
rect 3836 9938 4004 9940
rect 3836 9886 3838 9938
rect 3890 9886 4004 9938
rect 3836 9884 4004 9886
rect 4396 10388 4452 10398
rect 3836 9874 3892 9884
rect 4396 8484 4452 10332
rect 4614 10220 4878 10230
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4614 10154 4878 10164
rect 4956 10052 5012 10556
rect 5292 10546 5348 10556
rect 4844 9996 5012 10052
rect 4844 9380 4900 9996
rect 6300 9940 6356 11340
rect 7308 11396 7364 11406
rect 7308 11302 7364 11340
rect 7756 11394 7812 12012
rect 7756 11342 7758 11394
rect 7810 11342 7812 11394
rect 7756 11330 7812 11342
rect 7868 11396 7924 13022
rect 9884 12850 9940 13468
rect 9884 12798 9886 12850
rect 9938 12798 9940 12850
rect 9884 12786 9940 12798
rect 8016 12572 8280 12582
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8016 12506 8280 12516
rect 8428 12178 8484 12190
rect 8428 12126 8430 12178
rect 8482 12126 8484 12178
rect 8092 11396 8148 11406
rect 7868 11394 8148 11396
rect 7868 11342 8094 11394
rect 8146 11342 8148 11394
rect 7868 11340 8148 11342
rect 8092 11330 8148 11340
rect 6860 11172 6916 11182
rect 6860 11170 7028 11172
rect 6860 11118 6862 11170
rect 6914 11118 7028 11170
rect 6860 11116 7028 11118
rect 6860 11106 6916 11116
rect 6972 10834 7028 11116
rect 8016 11004 8280 11014
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8016 10938 8280 10948
rect 6972 10782 6974 10834
rect 7026 10782 7028 10834
rect 6972 10770 7028 10782
rect 8092 10836 8148 10846
rect 8092 10742 8148 10780
rect 7756 10388 7812 10398
rect 7532 10386 7812 10388
rect 7532 10334 7758 10386
rect 7810 10334 7812 10386
rect 7532 10332 7812 10334
rect 6636 9940 6692 9950
rect 6300 9938 6692 9940
rect 6300 9886 6638 9938
rect 6690 9886 6692 9938
rect 6300 9884 6692 9886
rect 6188 9828 6244 9838
rect 6300 9828 6356 9884
rect 6636 9874 6692 9884
rect 5852 9826 6356 9828
rect 5852 9774 6190 9826
rect 6242 9774 6356 9826
rect 5852 9772 6356 9774
rect 4844 9314 4900 9324
rect 4956 9714 5012 9726
rect 4956 9662 4958 9714
rect 5010 9662 5012 9714
rect 4614 8652 4878 8662
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4614 8586 4878 8596
rect 4508 8484 4564 8494
rect 4396 8482 4564 8484
rect 4396 8430 4510 8482
rect 4562 8430 4564 8482
rect 4396 8428 4564 8430
rect 4508 8418 4564 8428
rect 4844 8372 4900 8382
rect 4956 8372 5012 9662
rect 5628 9602 5684 9614
rect 5628 9550 5630 9602
rect 5682 9550 5684 9602
rect 5628 9266 5684 9550
rect 5628 9214 5630 9266
rect 5682 9214 5684 9266
rect 5628 9202 5684 9214
rect 5852 8372 5908 9772
rect 6188 9762 6244 9772
rect 7532 9714 7588 10332
rect 7756 10322 7812 10332
rect 8428 9938 8484 12126
rect 9100 12178 9156 12190
rect 9100 12126 9102 12178
rect 9154 12126 9156 12178
rect 9100 12068 9156 12126
rect 9100 12002 9156 12012
rect 8540 11396 8596 11406
rect 8540 10612 8596 11340
rect 8540 10610 9044 10612
rect 8540 10558 8542 10610
rect 8594 10558 9044 10610
rect 8540 10556 9044 10558
rect 8540 10546 8596 10556
rect 8428 9886 8430 9938
rect 8482 9886 8484 9938
rect 8428 9874 8484 9886
rect 8988 10500 9044 10556
rect 8988 9938 9044 10444
rect 9884 10500 9940 10510
rect 10108 10500 10164 13692
rect 10892 13682 10948 13692
rect 10444 13522 10500 13534
rect 10444 13470 10446 13522
rect 10498 13470 10500 13522
rect 10444 11282 10500 13470
rect 11228 13524 11284 15038
rect 11418 14924 11682 14934
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11418 14858 11682 14868
rect 11228 13458 11284 13468
rect 11788 13412 11844 15092
rect 11418 13356 11682 13366
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11788 13346 11844 13356
rect 12460 14306 12516 14318
rect 12460 14254 12462 14306
rect 12514 14254 12516 14306
rect 11418 13290 11682 13300
rect 12460 13188 12516 14254
rect 12460 13122 12516 13132
rect 12236 12962 12292 12974
rect 12236 12910 12238 12962
rect 12290 12910 12292 12962
rect 10444 11230 10446 11282
rect 10498 11230 10500 11282
rect 10444 11218 10500 11230
rect 10780 12068 10836 12078
rect 9940 10444 10164 10500
rect 9884 10406 9940 10444
rect 8988 9886 8990 9938
rect 9042 9886 9044 9938
rect 8988 9874 9044 9886
rect 10332 9828 10388 9838
rect 7532 9662 7534 9714
rect 7586 9662 7588 9714
rect 7532 9650 7588 9662
rect 10108 9826 10388 9828
rect 10108 9774 10334 9826
rect 10386 9774 10388 9826
rect 10108 9772 10388 9774
rect 8016 9436 8280 9446
rect 6636 9380 6692 9390
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8016 9370 8280 9380
rect 4956 8316 5572 8372
rect 4844 8258 4900 8316
rect 4844 8206 4846 8258
rect 4898 8206 4900 8258
rect 4844 8194 4900 8206
rect 3724 7756 4788 7812
rect 4732 7698 4788 7756
rect 4732 7646 4734 7698
rect 4786 7646 4788 7698
rect 4732 7634 4788 7646
rect 5516 7698 5572 8316
rect 5852 8278 5908 8316
rect 6412 8818 6468 8830
rect 6412 8766 6414 8818
rect 6466 8766 6468 8818
rect 6412 8148 6468 8766
rect 6636 8484 6692 9324
rect 6636 8428 6804 8484
rect 6748 8370 6804 8428
rect 6748 8318 6750 8370
rect 6802 8318 6804 8370
rect 6748 8306 6804 8318
rect 6412 8082 6468 8092
rect 7756 8148 7812 8158
rect 7756 8054 7812 8092
rect 8016 7868 8280 7878
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8016 7802 8280 7812
rect 5516 7646 5518 7698
rect 5570 7646 5572 7698
rect 5516 7634 5572 7646
rect 2044 7196 2772 7252
rect 4614 7084 4878 7094
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4614 7018 4878 7028
rect 1708 6466 1764 6478
rect 1708 6414 1710 6466
rect 1762 6414 1764 6466
rect 1708 6132 1764 6414
rect 8016 6300 8280 6310
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8016 6234 8280 6244
rect 1708 6066 1764 6076
rect 4614 5516 4878 5526
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4614 5450 4878 5460
rect 10108 5348 10164 9772
rect 10332 9762 10388 9772
rect 10780 9044 10836 12012
rect 11418 11788 11682 11798
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11418 11722 11682 11732
rect 11228 11172 11284 11182
rect 11228 11078 11284 11116
rect 12236 10500 12292 12910
rect 12572 12962 12628 15092
rect 14476 14644 14532 14654
rect 14476 14550 14532 14588
rect 13020 14420 13076 14430
rect 13020 14326 13076 14364
rect 14476 13746 14532 13758
rect 14476 13694 14478 13746
rect 14530 13694 14532 13746
rect 13916 13522 13972 13534
rect 13916 13470 13918 13522
rect 13970 13470 13972 13522
rect 13916 13412 13972 13470
rect 13468 13188 13524 13198
rect 13468 13094 13524 13132
rect 12572 12910 12574 12962
rect 12626 12910 12628 12962
rect 12572 12898 12628 12910
rect 13916 12962 13972 13356
rect 13916 12910 13918 12962
rect 13970 12910 13972 12962
rect 13916 12898 13972 12910
rect 14140 11396 14196 11406
rect 14476 11396 14532 13694
rect 14588 13076 14644 16830
rect 14700 16210 14756 17276
rect 14820 17276 15084 17286
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 14820 17210 15084 17220
rect 14700 16158 14702 16210
rect 14754 16158 14756 16210
rect 14700 16146 14756 16158
rect 16044 16884 16100 17612
rect 16156 17602 16212 17612
rect 16828 17666 16884 18172
rect 16940 18162 16996 18172
rect 16828 17614 16830 17666
rect 16882 17614 16884 17666
rect 16828 17602 16884 17614
rect 14820 15708 15084 15718
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 14820 15642 15084 15652
rect 15036 15316 15092 15326
rect 15036 15222 15092 15260
rect 15708 15316 15764 15326
rect 16044 15316 16100 16828
rect 17612 16884 17668 19966
rect 18060 20018 18116 20030
rect 18060 19966 18062 20018
rect 18114 19966 18116 20018
rect 18060 19348 18116 19966
rect 21084 20020 21140 20030
rect 21084 19926 21140 19964
rect 20748 19908 20804 19918
rect 18222 19628 18486 19638
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18222 19562 18486 19572
rect 18060 19282 18116 19292
rect 19180 19348 19236 19358
rect 19180 19254 19236 19292
rect 17948 19124 18004 19134
rect 17948 19030 18004 19068
rect 20188 19124 20244 19134
rect 20188 19030 20244 19068
rect 19404 18564 19460 18574
rect 19404 18470 19460 18508
rect 20188 18450 20244 18462
rect 20188 18398 20190 18450
rect 20242 18398 20244 18450
rect 18396 18338 18452 18350
rect 18396 18286 18398 18338
rect 18450 18286 18452 18338
rect 18396 18228 18452 18286
rect 18396 18162 18452 18172
rect 18222 18060 18486 18070
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18222 17994 18486 18004
rect 19292 17444 19348 17454
rect 19292 17350 19348 17388
rect 19852 17442 19908 17454
rect 19852 17390 19854 17442
rect 19906 17390 19908 17442
rect 17612 16818 17668 16828
rect 17948 16884 18004 16894
rect 17948 16790 18004 16828
rect 18620 16882 18676 16894
rect 18620 16830 18622 16882
rect 18674 16830 18676 16882
rect 18222 16492 18486 16502
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18222 16426 18486 16436
rect 18620 16212 18676 16830
rect 19292 16212 19348 16222
rect 18620 16210 19348 16212
rect 18620 16158 19294 16210
rect 19346 16158 19348 16210
rect 18620 16156 19348 16158
rect 19292 16146 19348 16156
rect 19852 15988 19908 17390
rect 20076 17444 20132 17454
rect 20076 17350 20132 17388
rect 19852 15922 19908 15932
rect 20076 16884 20132 16894
rect 20188 16884 20244 18398
rect 20748 18450 20804 19852
rect 21308 19458 21364 20132
rect 21308 19406 21310 19458
rect 21362 19406 21364 19458
rect 21308 19394 21364 19406
rect 21532 19906 21588 19918
rect 21532 19854 21534 19906
rect 21586 19854 21588 19906
rect 21532 19236 21588 19854
rect 20748 18398 20750 18450
rect 20802 18398 20804 18450
rect 20748 18386 20804 18398
rect 21420 19234 21588 19236
rect 21420 19182 21534 19234
rect 21586 19182 21588 19234
rect 21420 19180 21588 19182
rect 21868 19906 21924 19918
rect 21868 19854 21870 19906
rect 21922 19854 21924 19906
rect 21868 19236 21924 19854
rect 22316 19908 22372 19918
rect 22316 19814 22372 19852
rect 22428 19236 22484 19246
rect 21868 19234 22484 19236
rect 21868 19182 22430 19234
rect 22482 19182 22484 19234
rect 21868 19180 22484 19182
rect 21420 18340 21476 19180
rect 21532 19170 21588 19180
rect 21624 18844 21888 18854
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21624 18778 21888 18788
rect 21420 17778 21476 18284
rect 21420 17726 21422 17778
rect 21474 17726 21476 17778
rect 20132 16828 20244 16884
rect 20636 17668 20692 17678
rect 15708 15314 16100 15316
rect 15708 15262 15710 15314
rect 15762 15262 16046 15314
rect 16098 15262 16100 15314
rect 15708 15260 16100 15262
rect 15708 15250 15764 15260
rect 16044 15250 16100 15260
rect 20076 15314 20132 16828
rect 20300 15988 20356 15998
rect 20300 15894 20356 15932
rect 20076 15262 20078 15314
rect 20130 15262 20132 15314
rect 20076 15250 20132 15262
rect 20524 15316 20580 15326
rect 20524 15222 20580 15260
rect 18222 14924 18486 14934
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18222 14858 18486 14868
rect 20524 14532 20580 14542
rect 20636 14532 20692 17612
rect 21420 17668 21476 17726
rect 21420 17602 21476 17612
rect 21624 17276 21888 17286
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21624 17210 21888 17220
rect 21644 17108 21700 17118
rect 21644 17014 21700 17052
rect 20860 16994 20916 17006
rect 20860 16942 20862 16994
rect 20914 16942 20916 16994
rect 20748 14756 20804 14766
rect 20860 14756 20916 16942
rect 21980 16884 22036 16894
rect 22428 16884 22484 19180
rect 22876 19234 22932 20860
rect 24444 20916 24500 20926
rect 24444 20822 24500 20860
rect 23996 20578 24052 20590
rect 23996 20526 23998 20578
rect 24050 20526 24052 20578
rect 23548 20130 23604 20142
rect 23548 20078 23550 20130
rect 23602 20078 23604 20130
rect 23548 20020 23604 20078
rect 23548 19954 23604 19964
rect 23772 20020 23828 20030
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22876 19170 22932 19182
rect 23212 19796 23268 19806
rect 23212 18674 23268 19740
rect 23212 18622 23214 18674
rect 23266 18622 23268 18674
rect 23212 18610 23268 18622
rect 23772 18450 23828 19964
rect 23996 19908 24052 20526
rect 24556 20132 24612 23774
rect 24668 23828 24724 24556
rect 25116 24500 25172 25228
rect 25340 25218 25396 25228
rect 25452 24948 25508 26012
rect 25900 25618 25956 26908
rect 26124 26516 26180 26526
rect 26124 26422 26180 26460
rect 25900 25566 25902 25618
rect 25954 25566 25956 25618
rect 25900 25554 25956 25566
rect 26124 26292 26180 26302
rect 26572 26292 26628 26302
rect 25452 24854 25508 24892
rect 25564 25284 25620 25294
rect 24668 23762 24724 23772
rect 24892 24444 25172 24500
rect 24892 23826 24948 24444
rect 25026 24332 25290 24342
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25026 24266 25290 24276
rect 25228 23940 25284 23950
rect 25228 23846 25284 23884
rect 24892 23774 24894 23826
rect 24946 23774 24948 23826
rect 24892 23762 24948 23774
rect 25564 23826 25620 25228
rect 25900 24836 25956 24846
rect 25900 23938 25956 24780
rect 26124 24610 26180 26236
rect 26124 24558 26126 24610
rect 26178 24558 26180 24610
rect 26124 24546 26180 24558
rect 26236 26290 26628 26292
rect 26236 26238 26574 26290
rect 26626 26238 26628 26290
rect 26236 26236 26628 26238
rect 25900 23886 25902 23938
rect 25954 23886 25956 23938
rect 25900 23874 25956 23886
rect 25564 23774 25566 23826
rect 25618 23774 25620 23826
rect 25564 23762 25620 23774
rect 26236 23826 26292 26236
rect 26572 26226 26628 26236
rect 26908 25284 26964 25294
rect 26908 25190 26964 25228
rect 26236 23774 26238 23826
rect 26290 23774 26292 23826
rect 26236 23762 26292 23774
rect 26572 24722 26628 24734
rect 26572 24670 26574 24722
rect 26626 24670 26628 24722
rect 25788 23716 25844 23726
rect 25676 23660 25788 23716
rect 25564 23380 25620 23390
rect 25676 23380 25732 23660
rect 25788 23650 25844 23660
rect 25564 23378 25732 23380
rect 25564 23326 25566 23378
rect 25618 23326 25732 23378
rect 25564 23324 25732 23326
rect 25564 23314 25620 23324
rect 24668 23268 24724 23278
rect 24668 23174 24724 23212
rect 26236 23266 26292 23278
rect 26236 23214 26238 23266
rect 26290 23214 26292 23266
rect 25340 23156 25396 23166
rect 26012 23156 26068 23166
rect 25340 23154 25508 23156
rect 25340 23102 25342 23154
rect 25394 23102 25508 23154
rect 25340 23100 25508 23102
rect 25340 23090 25396 23100
rect 25026 22764 25290 22774
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25026 22698 25290 22708
rect 25452 21700 25508 23100
rect 26012 23154 26180 23156
rect 26012 23102 26014 23154
rect 26066 23102 26180 23154
rect 26012 23100 26180 23102
rect 26012 23090 26068 23100
rect 26124 22484 26180 23100
rect 26236 22820 26292 23214
rect 26236 22754 26292 22764
rect 26124 22428 26516 22484
rect 25676 22372 25732 22382
rect 25676 22370 25844 22372
rect 25676 22318 25678 22370
rect 25730 22318 25844 22370
rect 25676 22316 25844 22318
rect 25676 22306 25732 22316
rect 25452 21644 25620 21700
rect 25026 21196 25290 21206
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25026 21130 25290 21140
rect 25452 20690 25508 20702
rect 25452 20638 25454 20690
rect 25506 20638 25508 20690
rect 25452 20188 25508 20638
rect 24556 20066 24612 20076
rect 25340 20132 25508 20188
rect 23996 19842 24052 19852
rect 24444 20018 24500 20030
rect 24444 19966 24446 20018
rect 24498 19966 24500 20018
rect 24108 19796 24164 19806
rect 24108 19702 24164 19740
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 23772 18386 23828 18398
rect 23884 19012 23940 19022
rect 23100 18340 23156 18350
rect 23100 17780 23156 18284
rect 22652 17778 23156 17780
rect 22652 17726 23102 17778
rect 23154 17726 23156 17778
rect 22652 17724 23156 17726
rect 22652 17666 22708 17724
rect 23100 17714 23156 17724
rect 22652 17614 22654 17666
rect 22706 17614 22708 17666
rect 22652 17602 22708 17614
rect 22540 17444 22596 17454
rect 22540 17442 22820 17444
rect 22540 17390 22542 17442
rect 22594 17390 22820 17442
rect 22540 17388 22820 17390
rect 22540 17378 22596 17388
rect 22036 16882 22484 16884
rect 22036 16830 22430 16882
rect 22482 16830 22484 16882
rect 22036 16828 22484 16830
rect 21980 16790 22036 16828
rect 21980 16098 22036 16110
rect 21980 16046 21982 16098
rect 22034 16046 22036 16098
rect 21624 15708 21888 15718
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21624 15642 21888 15652
rect 20748 14754 20916 14756
rect 20748 14702 20750 14754
rect 20802 14702 20916 14754
rect 20748 14700 20916 14702
rect 20748 14690 20804 14700
rect 20524 14530 20692 14532
rect 20524 14478 20526 14530
rect 20578 14478 20692 14530
rect 20524 14476 20692 14478
rect 15484 14420 15540 14430
rect 15484 14326 15540 14364
rect 18060 14308 18116 14318
rect 14820 14140 15084 14150
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 14820 14074 15084 14084
rect 14588 12178 14644 13020
rect 16828 13076 16884 13086
rect 16828 12982 16884 13020
rect 15148 12964 15204 12974
rect 15204 12908 15316 12964
rect 15148 12870 15204 12908
rect 14820 12572 15084 12582
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 14820 12506 15084 12516
rect 15260 12402 15316 12908
rect 15260 12350 15262 12402
rect 15314 12350 15316 12402
rect 15260 12338 15316 12350
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 14588 12114 14644 12126
rect 18060 11506 18116 14252
rect 19852 14308 19908 14318
rect 20524 14308 20580 14476
rect 19908 14252 20580 14308
rect 19852 14214 19908 14252
rect 21624 14140 21888 14150
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21624 14074 21888 14084
rect 18844 13860 18900 13870
rect 18844 13858 19796 13860
rect 18844 13806 18846 13858
rect 18898 13806 19796 13858
rect 18844 13804 19796 13806
rect 18844 13794 18900 13804
rect 18222 13356 18486 13366
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18222 13290 18486 13300
rect 19740 12402 19796 13804
rect 21308 13746 21364 13758
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 19740 12350 19742 12402
rect 19794 12350 19796 12402
rect 19740 12338 19796 12350
rect 19852 13634 19908 13646
rect 19852 13582 19854 13634
rect 19906 13582 19908 13634
rect 19628 11844 19684 11854
rect 18222 11788 18486 11798
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18222 11722 18486 11732
rect 18060 11454 18062 11506
rect 18114 11454 18116 11506
rect 18060 11442 18116 11454
rect 14140 11394 14532 11396
rect 14140 11342 14142 11394
rect 14194 11342 14478 11394
rect 14530 11342 14532 11394
rect 14140 11340 14532 11342
rect 13804 11284 13860 11294
rect 13692 11282 13860 11284
rect 13692 11230 13806 11282
rect 13858 11230 13860 11282
rect 13692 11228 13860 11230
rect 12236 10434 12292 10444
rect 12684 10612 12740 10622
rect 11418 10220 11682 10230
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11418 10154 11682 10164
rect 12684 10050 12740 10556
rect 13468 10612 13524 10622
rect 13468 10518 13524 10556
rect 12684 9998 12686 10050
rect 12738 9998 12740 10050
rect 12684 9986 12740 9998
rect 10780 7474 10836 8988
rect 12236 9044 12292 9054
rect 12236 8950 12292 8988
rect 12908 9042 12964 9054
rect 12908 8990 12910 9042
rect 12962 8990 12964 9042
rect 11418 8652 11682 8662
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11418 8586 11682 8596
rect 12908 7924 12964 8990
rect 12908 7858 12964 7868
rect 13692 7698 13748 11228
rect 13804 11218 13860 11228
rect 14140 10612 14196 11340
rect 14476 11330 14532 11340
rect 15820 11172 15876 11182
rect 14820 11004 15084 11014
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 14820 10938 15084 10948
rect 15820 10722 15876 11116
rect 15820 10670 15822 10722
rect 15874 10670 15876 10722
rect 15820 10658 15876 10670
rect 14140 9826 14196 10556
rect 17500 10612 17556 10622
rect 14812 10500 14868 10510
rect 14812 10406 14868 10444
rect 17500 10050 17556 10556
rect 18284 10612 18340 10622
rect 18284 10518 18340 10556
rect 19628 10610 19684 11788
rect 19628 10558 19630 10610
rect 19682 10558 19684 10610
rect 19628 10546 19684 10558
rect 19852 10612 19908 13582
rect 20524 12290 20580 12302
rect 20524 12238 20526 12290
rect 20578 12238 20580 12290
rect 20524 11508 20580 12238
rect 21308 11844 21364 13694
rect 21756 13748 21812 13758
rect 21756 13654 21812 13692
rect 21980 13076 22036 16046
rect 22428 15204 22484 16828
rect 22764 15538 22820 17388
rect 23324 17442 23380 17454
rect 23324 17390 23326 17442
rect 23378 17390 23380 17442
rect 23324 16996 23380 17390
rect 23884 17442 23940 18956
rect 24444 18450 24500 19966
rect 25340 20020 25396 20132
rect 25340 19954 25396 19964
rect 25452 19906 25508 19918
rect 25452 19854 25454 19906
rect 25506 19854 25508 19906
rect 25452 19794 25508 19854
rect 25452 19742 25454 19794
rect 25506 19742 25508 19794
rect 25026 19628 25290 19638
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25026 19562 25290 19572
rect 25116 19012 25172 19022
rect 24668 19010 25172 19012
rect 24668 18958 25118 19010
rect 25170 18958 25172 19010
rect 24668 18956 25172 18958
rect 24668 18674 24724 18956
rect 25116 18946 25172 18956
rect 24668 18622 24670 18674
rect 24722 18622 24724 18674
rect 24668 18610 24724 18622
rect 24444 18398 24446 18450
rect 24498 18398 24500 18450
rect 24444 18340 24500 18398
rect 24444 18274 24500 18284
rect 25340 18340 25396 18350
rect 25452 18340 25508 19742
rect 25396 18284 25508 18340
rect 25340 18246 25396 18284
rect 25026 18060 25290 18070
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25026 17994 25290 18004
rect 23884 17390 23886 17442
rect 23938 17390 23940 17442
rect 23884 17378 23940 17390
rect 23324 16930 23380 16940
rect 23996 16996 24052 17006
rect 23996 16902 24052 16940
rect 22764 15486 22766 15538
rect 22818 15486 22820 15538
rect 22764 15474 22820 15486
rect 22876 16770 22932 16782
rect 22876 16718 22878 16770
rect 22930 16718 22932 16770
rect 22876 15540 22932 16718
rect 25026 16492 25290 16502
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25026 16426 25290 16436
rect 22876 15474 22932 15484
rect 24556 15428 24612 15438
rect 24556 15314 24612 15372
rect 24556 15262 24558 15314
rect 24610 15262 24612 15314
rect 24556 15250 24612 15262
rect 25340 15428 25396 15438
rect 22092 15148 22428 15204
rect 22092 14530 22148 15148
rect 22428 15138 22484 15148
rect 23212 15204 23268 15214
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 22092 14466 22148 14478
rect 22540 14530 22596 14542
rect 22540 14478 22542 14530
rect 22594 14478 22596 14530
rect 22540 13636 22596 14478
rect 22540 13570 22596 13580
rect 21624 12572 21888 12582
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21624 12506 21888 12516
rect 21308 11778 21364 11788
rect 20524 11442 20580 11452
rect 20300 11394 20356 11406
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 19964 10612 20020 10622
rect 19852 10610 20020 10612
rect 19852 10558 19966 10610
rect 20018 10558 20020 10610
rect 19852 10556 20020 10558
rect 19964 10546 20020 10556
rect 20300 10612 20356 11342
rect 21980 11394 22036 13020
rect 23212 12962 23268 15148
rect 25340 15204 25396 15372
rect 25452 15204 25508 18284
rect 25564 17556 25620 21644
rect 25788 21252 25844 22316
rect 26236 22258 26292 22270
rect 26236 22206 26238 22258
rect 26290 22206 26292 22258
rect 25788 21186 25844 21196
rect 25900 22146 25956 22158
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25900 20804 25956 22094
rect 26236 21812 26292 22206
rect 26236 21746 26292 21756
rect 26460 21810 26516 22428
rect 26572 22258 26628 24670
rect 26908 24722 26964 24734
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26908 24164 26964 24670
rect 26908 24098 26964 24108
rect 26908 23716 26964 23726
rect 26908 23622 26964 23660
rect 26908 23268 26964 23278
rect 26908 23174 26964 23212
rect 27468 23042 27524 27580
rect 27692 26178 27748 26190
rect 27692 26126 27694 26178
rect 27746 26126 27748 26178
rect 27692 25620 27748 26126
rect 27692 25554 27748 25564
rect 27692 25282 27748 25294
rect 27692 25230 27694 25282
rect 27746 25230 27748 25282
rect 27692 24948 27748 25230
rect 27692 24882 27748 24892
rect 27692 24164 27748 24174
rect 27804 24164 27860 28924
rect 28428 26684 28692 26694
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28428 26618 28692 26628
rect 28428 25116 28692 25126
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28428 25050 28692 25060
rect 28028 24610 28084 24622
rect 28028 24558 28030 24610
rect 28082 24558 28084 24610
rect 28028 24276 28084 24558
rect 28028 24210 28084 24220
rect 27692 24162 27860 24164
rect 27692 24110 27694 24162
rect 27746 24110 27860 24162
rect 27692 24108 27860 24110
rect 27692 24098 27748 24108
rect 28428 23548 28692 23558
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28428 23482 28692 23492
rect 27468 22990 27470 23042
rect 27522 22990 27524 23042
rect 27468 22978 27524 22990
rect 28252 23042 28308 23054
rect 28252 22990 28254 23042
rect 28306 22990 28308 23042
rect 26572 22206 26574 22258
rect 26626 22206 26628 22258
rect 26572 22194 26628 22206
rect 26796 22932 26852 22942
rect 26460 21758 26462 21810
rect 26514 21758 26516 21810
rect 26460 21746 26516 21758
rect 26796 21698 26852 22876
rect 26908 22820 26964 22830
rect 26908 22370 26964 22764
rect 26908 22318 26910 22370
rect 26962 22318 26964 22370
rect 26908 22306 26964 22318
rect 28028 22260 28084 22270
rect 28028 22166 28084 22204
rect 27804 21812 27860 21822
rect 27804 21718 27860 21756
rect 26796 21646 26798 21698
rect 26850 21646 26852 21698
rect 26684 21588 26740 21598
rect 26236 21476 26292 21486
rect 26236 21382 26292 21420
rect 26684 20914 26740 21532
rect 26796 21476 26852 21646
rect 27132 21700 27188 21710
rect 27132 21606 27188 21644
rect 27468 21588 27524 21598
rect 27468 21494 27524 21532
rect 28140 21588 28196 21598
rect 28252 21588 28308 22990
rect 28428 21980 28692 21990
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28428 21914 28692 21924
rect 28140 21586 28308 21588
rect 28140 21534 28142 21586
rect 28194 21534 28308 21586
rect 28140 21532 28308 21534
rect 26796 21410 26852 21420
rect 26684 20862 26686 20914
rect 26738 20862 26740 20914
rect 26684 20850 26740 20862
rect 27468 21252 27524 21262
rect 25900 20738 25956 20748
rect 26908 20804 26964 20814
rect 26908 20710 26964 20748
rect 25900 19906 25956 19918
rect 25900 19854 25902 19906
rect 25954 19854 25956 19906
rect 25900 19794 25956 19854
rect 25900 19742 25902 19794
rect 25954 19742 25956 19794
rect 25900 19730 25956 19742
rect 26236 19908 26292 19918
rect 25900 19010 25956 19022
rect 25900 18958 25902 19010
rect 25954 18958 25956 19010
rect 25900 18562 25956 18958
rect 26124 19012 26180 19022
rect 26124 18918 26180 18956
rect 25900 18510 25902 18562
rect 25954 18510 25956 18562
rect 25900 18498 25956 18510
rect 26236 17892 26292 19852
rect 27468 19572 27524 21196
rect 28140 20916 28196 21532
rect 28140 20850 28196 20860
rect 28028 20690 28084 20702
rect 28028 20638 28030 20690
rect 28082 20638 28084 20690
rect 28028 20244 28084 20638
rect 28428 20412 28692 20422
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28428 20346 28692 20356
rect 28028 20178 28084 20188
rect 27804 20132 27860 20142
rect 27804 20038 27860 20076
rect 28140 20018 28196 20030
rect 28140 19966 28142 20018
rect 28194 19966 28196 20018
rect 27580 19908 27636 19918
rect 28140 19908 28196 19966
rect 27580 19906 28196 19908
rect 27580 19854 27582 19906
rect 27634 19854 28196 19906
rect 27580 19852 28196 19854
rect 27580 19842 27636 19852
rect 28140 19572 28196 19852
rect 27468 19516 27860 19572
rect 26348 19234 26404 19246
rect 26348 19182 26350 19234
rect 26402 19182 26404 19234
rect 26348 18340 26404 19182
rect 27804 19122 27860 19516
rect 28140 19506 28196 19516
rect 27804 19070 27806 19122
rect 27858 19070 27860 19122
rect 27804 19058 27860 19070
rect 28140 19122 28196 19134
rect 28140 19070 28142 19122
rect 28194 19070 28196 19122
rect 27580 19012 27636 19022
rect 27580 18918 27636 18956
rect 28140 19012 28196 19070
rect 28140 18946 28196 18956
rect 28428 18844 28692 18854
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28428 18778 28692 18788
rect 26348 18274 26404 18284
rect 27132 18338 27188 18350
rect 27132 18286 27134 18338
rect 27186 18286 27188 18338
rect 26236 17836 26516 17892
rect 26348 17668 26404 17678
rect 26460 17668 26516 17836
rect 27020 17668 27076 17678
rect 26460 17666 27076 17668
rect 26460 17614 27022 17666
rect 27074 17614 27076 17666
rect 26460 17612 27076 17614
rect 26348 17574 26404 17612
rect 25564 17490 25620 17500
rect 27020 17444 27076 17612
rect 27132 17668 27188 18286
rect 27692 18338 27748 18350
rect 27692 18286 27694 18338
rect 27746 18286 27748 18338
rect 27692 18228 27748 18286
rect 27692 18162 27748 18172
rect 28140 18228 28196 18238
rect 27132 17602 27188 17612
rect 28140 17666 28196 18172
rect 28140 17614 28142 17666
rect 28194 17614 28196 17666
rect 28140 17602 28196 17614
rect 27804 17556 27860 17566
rect 27804 17462 27860 17500
rect 27356 17444 27412 17454
rect 27020 17442 27412 17444
rect 27020 17390 27358 17442
rect 27410 17390 27412 17442
rect 27020 17388 27412 17390
rect 27244 17108 27300 17118
rect 26684 16770 26740 16782
rect 26684 16718 26686 16770
rect 26738 16718 26740 16770
rect 25788 15986 25844 15998
rect 25788 15934 25790 15986
rect 25842 15934 25844 15986
rect 25340 15202 25508 15204
rect 25340 15150 25342 15202
rect 25394 15150 25508 15202
rect 25340 15148 25508 15150
rect 25340 15138 25396 15148
rect 23548 15092 23604 15102
rect 23548 14998 23604 15036
rect 24444 15092 24500 15102
rect 24444 15090 24836 15092
rect 24444 15038 24446 15090
rect 24498 15038 24836 15090
rect 24444 15036 24836 15038
rect 24444 15026 24500 15036
rect 23212 12910 23214 12962
rect 23266 12910 23268 12962
rect 23212 12898 23268 12910
rect 23660 14756 23716 14766
rect 23660 12962 23716 14700
rect 24780 14418 24836 15036
rect 25026 14924 25290 14934
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25026 14858 25290 14868
rect 24780 14366 24782 14418
rect 24834 14366 24836 14418
rect 24780 14354 24836 14366
rect 25452 14532 25508 15148
rect 25564 15652 25620 15662
rect 25564 14754 25620 15596
rect 25788 15204 25844 15934
rect 25788 15110 25844 15148
rect 26236 15316 26292 15326
rect 26236 15202 26292 15260
rect 26236 15150 26238 15202
rect 26290 15150 26292 15202
rect 26236 15138 26292 15150
rect 25564 14702 25566 14754
rect 25618 14702 25620 14754
rect 25564 14690 25620 14702
rect 26684 14756 26740 16718
rect 27244 15426 27300 17052
rect 27244 15374 27246 15426
rect 27298 15374 27300 15426
rect 27244 15362 27300 15374
rect 27356 15204 27412 17388
rect 28428 17276 28692 17286
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28428 17210 28692 17220
rect 27692 16994 27748 17006
rect 27692 16942 27694 16994
rect 27746 16942 27748 16994
rect 27692 15652 27748 16942
rect 28428 15708 28692 15718
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28428 15642 28692 15652
rect 27692 15586 27748 15596
rect 27356 15138 27412 15148
rect 27692 15204 27748 15214
rect 26684 14690 26740 14700
rect 27244 15092 27300 15102
rect 24220 14308 24276 14318
rect 24220 13970 24276 14252
rect 24220 13918 24222 13970
rect 24274 13918 24276 13970
rect 24220 13906 24276 13918
rect 25452 13970 25508 14476
rect 25452 13918 25454 13970
rect 25506 13918 25508 13970
rect 25452 13906 25508 13918
rect 25900 14642 25956 14654
rect 25900 14590 25902 14642
rect 25954 14590 25956 14642
rect 24780 13524 24836 13534
rect 24780 13430 24836 13468
rect 25026 13356 25290 13366
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25026 13290 25290 13300
rect 23660 12910 23662 12962
rect 23714 12910 23716 12962
rect 23660 12898 23716 12910
rect 25900 12850 25956 14590
rect 26348 14532 26404 14542
rect 26348 14438 26404 14476
rect 27132 14532 27188 14542
rect 27132 14438 27188 14476
rect 26684 14308 26740 14318
rect 26684 14214 26740 14252
rect 27244 13858 27300 15036
rect 27244 13806 27246 13858
rect 27298 13806 27300 13858
rect 27244 13794 27300 13806
rect 27692 14306 27748 15148
rect 28140 14532 28196 14542
rect 28140 14438 28196 14476
rect 27692 14254 27694 14306
rect 27746 14254 27748 14306
rect 26460 13748 26516 13758
rect 25900 12798 25902 12850
rect 25954 12798 25956 12850
rect 25900 12786 25956 12798
rect 26012 13634 26068 13646
rect 26012 13582 26014 13634
rect 26066 13582 26068 13634
rect 22876 12178 22932 12190
rect 22876 12126 22878 12178
rect 22930 12126 22932 12178
rect 22876 11956 22932 12126
rect 22876 11890 22932 11900
rect 23436 12178 23492 12190
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 21980 11342 21982 11394
rect 22034 11342 22036 11394
rect 21980 11330 22036 11342
rect 23436 11732 23492 12126
rect 24556 12178 24612 12190
rect 24556 12126 24558 12178
rect 24610 12126 24612 12178
rect 23436 11284 23492 11676
rect 24108 11954 24164 11966
rect 24108 11902 24110 11954
rect 24162 11902 24164 11954
rect 23660 11508 23716 11518
rect 23716 11452 23828 11508
rect 23660 11442 23716 11452
rect 23436 11218 23492 11228
rect 20748 11172 20804 11182
rect 20748 11078 20804 11116
rect 22316 11172 22372 11182
rect 21624 11004 21888 11014
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21624 10938 21888 10948
rect 22316 10834 22372 11116
rect 22316 10782 22318 10834
rect 22370 10782 22372 10834
rect 22316 10770 22372 10782
rect 23772 10834 23828 11452
rect 23772 10782 23774 10834
rect 23826 10782 23828 10834
rect 23772 10770 23828 10782
rect 23100 10724 23156 10734
rect 23100 10630 23156 10668
rect 20300 10546 20356 10556
rect 23884 10612 23940 10622
rect 23884 10518 23940 10556
rect 21980 10500 22036 10510
rect 17500 9998 17502 10050
rect 17554 9998 17556 10050
rect 17500 9986 17556 9998
rect 18060 10386 18116 10398
rect 18060 10334 18062 10386
rect 18114 10334 18116 10386
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 14140 8820 14196 9774
rect 14820 9436 15084 9446
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 14820 9370 15084 9380
rect 15372 9268 15428 9278
rect 16268 9268 16324 9278
rect 15372 9266 16324 9268
rect 15372 9214 15374 9266
rect 15426 9214 16270 9266
rect 16322 9214 16324 9266
rect 15372 9212 16324 9214
rect 15372 9202 15428 9212
rect 16268 9202 16324 9212
rect 15932 9044 15988 9054
rect 15932 8950 15988 8988
rect 17276 9042 17332 9054
rect 17276 8990 17278 9042
rect 17330 8990 17332 9042
rect 14140 8754 14196 8764
rect 15372 8932 15428 8942
rect 14924 8260 14980 8270
rect 14924 8166 14980 8204
rect 15372 8258 15428 8876
rect 16156 8930 16212 8942
rect 16156 8878 16158 8930
rect 16210 8878 16212 8930
rect 16156 8820 16212 8878
rect 16156 8754 16212 8764
rect 15372 8206 15374 8258
rect 15426 8206 15428 8258
rect 15372 8194 15428 8206
rect 17276 8260 17332 8990
rect 17948 9042 18004 9054
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 8372 18004 8990
rect 17948 8306 18004 8316
rect 17276 8194 17332 8204
rect 17836 8036 17892 8046
rect 18060 8036 18116 10334
rect 18222 10220 18486 10230
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18222 10154 18486 10164
rect 19068 9938 19124 9950
rect 19068 9886 19070 9938
rect 19122 9886 19124 9938
rect 19068 8932 19124 9886
rect 20748 9828 20804 9838
rect 20412 9714 20468 9726
rect 20412 9662 20414 9714
rect 20466 9662 20468 9714
rect 19068 8866 19124 8876
rect 19292 9156 19348 9166
rect 18222 8652 18486 8662
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18222 8586 18486 8596
rect 19292 8370 19348 9100
rect 20188 9156 20244 9166
rect 20188 9062 20244 9100
rect 20412 9044 20468 9662
rect 20412 8978 20468 8988
rect 19292 8318 19294 8370
rect 19346 8318 19348 8370
rect 19292 8306 19348 8318
rect 19516 8372 19572 8382
rect 18508 8260 18564 8270
rect 17836 8034 18116 8036
rect 17836 7982 17838 8034
rect 17890 7982 18116 8034
rect 17836 7980 18116 7982
rect 18396 8034 18452 8046
rect 18396 7982 18398 8034
rect 18450 7982 18452 8034
rect 17836 7970 17892 7980
rect 13692 7646 13694 7698
rect 13746 7646 13748 7698
rect 13692 7634 13748 7646
rect 14476 7924 14532 7934
rect 10780 7422 10782 7474
rect 10834 7422 10836 7474
rect 10780 7410 10836 7422
rect 11228 7474 11284 7486
rect 11228 7422 11230 7474
rect 11282 7422 11284 7474
rect 11228 6804 11284 7422
rect 14252 7250 14308 7262
rect 14252 7198 14254 7250
rect 14306 7198 14308 7250
rect 11418 7084 11682 7094
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11418 7018 11682 7028
rect 11228 6738 11284 6748
rect 14252 6580 14308 7198
rect 14476 6802 14532 7868
rect 14820 7868 15084 7878
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 14820 7802 15084 7812
rect 18396 7252 18452 7982
rect 18508 7700 18564 8204
rect 19068 8258 19124 8270
rect 19068 8206 19070 8258
rect 19122 8206 19124 8258
rect 19068 8148 19124 8206
rect 19068 8082 19124 8092
rect 18508 7606 18564 7644
rect 19292 7700 19348 7710
rect 19292 7474 19348 7644
rect 19292 7422 19294 7474
rect 19346 7422 19348 7474
rect 19292 7410 19348 7422
rect 18060 7196 18452 7252
rect 14476 6750 14478 6802
rect 14530 6750 14532 6802
rect 14476 6738 14532 6750
rect 17276 6804 17332 6814
rect 17276 6710 17332 6748
rect 18060 6692 18116 7196
rect 18222 7084 18486 7094
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18222 7018 18486 7028
rect 18060 6626 18116 6636
rect 18620 6916 18676 6926
rect 14252 6514 14308 6524
rect 15484 6580 15540 6590
rect 15484 6486 15540 6524
rect 18620 6578 18676 6860
rect 18620 6526 18622 6578
rect 18674 6526 18676 6578
rect 18620 6514 18676 6526
rect 14820 6300 15084 6310
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 14820 6234 15084 6244
rect 19516 5794 19572 8316
rect 20748 8034 20804 9772
rect 21532 9828 21588 9838
rect 21532 9734 21588 9772
rect 21980 9826 22036 10444
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21980 9762 22036 9774
rect 21624 9436 21888 9446
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21624 9370 21888 9380
rect 24108 9380 24164 11902
rect 24332 11284 24388 11294
rect 24332 10498 24388 11228
rect 24332 10446 24334 10498
rect 24386 10446 24388 10498
rect 24332 9828 24388 10446
rect 24108 9324 24276 9380
rect 21868 9156 21924 9166
rect 23548 9156 23604 9166
rect 21868 9154 22820 9156
rect 21868 9102 21870 9154
rect 21922 9102 22820 9154
rect 21868 9100 22820 9102
rect 21868 9090 21924 9100
rect 20748 7982 20750 8034
rect 20802 7982 20804 8034
rect 20748 7700 20804 7982
rect 19516 5742 19518 5794
rect 19570 5742 19572 5794
rect 19516 5730 19572 5742
rect 19964 7474 20020 7486
rect 19964 7422 19966 7474
rect 20018 7422 20020 7474
rect 19964 5796 20020 7422
rect 20748 7364 20804 7644
rect 20748 7298 20804 7308
rect 20972 8818 21028 8830
rect 20972 8766 20974 8818
rect 21026 8766 21028 8818
rect 20972 7252 21028 8766
rect 20972 7186 21028 7196
rect 21084 8818 21140 8830
rect 21084 8766 21086 8818
rect 21138 8766 21140 8818
rect 21084 6916 21140 8766
rect 22764 8482 22820 9100
rect 22764 8430 22766 8482
rect 22818 8430 22820 8482
rect 22764 8418 22820 8430
rect 23548 8370 23604 9100
rect 24108 9042 24164 9054
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 24108 8820 24164 8990
rect 24108 8754 24164 8764
rect 23548 8318 23550 8370
rect 23602 8318 23604 8370
rect 23548 8306 23604 8318
rect 21420 8258 21476 8270
rect 21420 8206 21422 8258
rect 21474 8206 21476 8258
rect 21420 8148 21476 8206
rect 21420 8082 21476 8092
rect 22988 8258 23044 8270
rect 22988 8206 22990 8258
rect 23042 8206 23044 8258
rect 22988 8148 23044 8206
rect 22988 8082 23044 8092
rect 21980 8036 22036 8046
rect 21980 8034 22260 8036
rect 21980 7982 21982 8034
rect 22034 7982 22260 8034
rect 21980 7980 22260 7982
rect 21980 7970 22036 7980
rect 21624 7868 21888 7878
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21624 7802 21888 7812
rect 22204 7698 22260 7980
rect 24220 8034 24276 9324
rect 24332 9044 24388 9772
rect 24444 11172 24500 11182
rect 24444 9602 24500 11116
rect 24556 10612 24612 12126
rect 25340 12068 25396 12078
rect 26012 12068 26068 13582
rect 26236 13636 26292 13646
rect 26236 13542 26292 13580
rect 25340 12066 26068 12068
rect 25340 12014 25342 12066
rect 25394 12014 26068 12066
rect 25340 12012 26068 12014
rect 26348 13524 26404 13534
rect 25340 12002 25396 12012
rect 25026 11788 25290 11798
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25026 11722 25290 11732
rect 24556 10546 24612 10556
rect 25026 10220 25290 10230
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25026 10154 25290 10164
rect 25004 9604 25060 9614
rect 24444 9550 24446 9602
rect 24498 9550 24500 9602
rect 24444 9538 24500 9550
rect 24892 9602 25060 9604
rect 24892 9550 25006 9602
rect 25058 9550 25060 9602
rect 24892 9548 25060 9550
rect 24668 9044 24724 9054
rect 24332 8988 24668 9044
rect 24668 8950 24724 8988
rect 24220 7982 24222 8034
rect 24274 7982 24276 8034
rect 24220 7970 24276 7982
rect 24332 8148 24388 8158
rect 22204 7646 22206 7698
rect 22258 7646 22260 7698
rect 22204 7634 22260 7646
rect 24332 7474 24388 8092
rect 24892 7588 24948 9548
rect 25004 9538 25060 9548
rect 25340 9604 25396 9614
rect 25452 9604 25508 12012
rect 25340 9602 25508 9604
rect 25340 9550 25342 9602
rect 25394 9550 25508 9602
rect 25340 9548 25508 9550
rect 26124 11956 26180 11966
rect 25340 9044 25396 9548
rect 25340 8932 25396 8988
rect 26124 8932 26180 11900
rect 26236 10500 26292 10510
rect 26236 10406 26292 10444
rect 26348 9714 26404 13468
rect 26460 12066 26516 13692
rect 27132 13076 27188 13086
rect 27692 13076 27748 14254
rect 28428 14140 28692 14150
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28428 14074 28692 14084
rect 27132 13074 27748 13076
rect 27132 13022 27134 13074
rect 27186 13022 27748 13074
rect 27132 13020 27748 13022
rect 27132 13010 27188 13020
rect 26684 12738 26740 12750
rect 26684 12686 26686 12738
rect 26738 12686 26740 12738
rect 26684 12292 26740 12686
rect 28428 12572 28692 12582
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28428 12506 28692 12516
rect 26684 12226 26740 12236
rect 27356 12292 27412 12302
rect 27356 12198 27412 12236
rect 26460 12014 26462 12066
rect 26514 12014 26516 12066
rect 26460 12002 26516 12014
rect 27356 11394 27412 11406
rect 27356 11342 27358 11394
rect 27410 11342 27412 11394
rect 26908 11172 26964 11182
rect 26908 11078 26964 11116
rect 27244 10724 27300 10734
rect 27244 10630 27300 10668
rect 27356 10612 27412 11342
rect 28428 11004 28692 11014
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28428 10938 28692 10948
rect 26348 9662 26350 9714
rect 26402 9662 26404 9714
rect 26348 9650 26404 9662
rect 26684 9940 26740 9950
rect 26236 8932 26292 8942
rect 25340 8930 25508 8932
rect 25340 8878 25342 8930
rect 25394 8878 25508 8930
rect 25340 8876 25508 8878
rect 26124 8930 26292 8932
rect 26124 8878 26238 8930
rect 26290 8878 26292 8930
rect 26124 8876 26292 8878
rect 25340 8866 25396 8876
rect 25026 8652 25290 8662
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25026 8586 25290 8596
rect 25452 8484 25508 8876
rect 26236 8866 26292 8876
rect 25452 8418 25508 8428
rect 26460 8820 26516 8830
rect 24892 7522 24948 7532
rect 25788 8036 25844 8046
rect 24332 7422 24334 7474
rect 24386 7422 24388 7474
rect 24332 7410 24388 7422
rect 21084 6850 21140 6860
rect 22652 7364 22708 7374
rect 20300 6692 20356 6702
rect 20300 6018 20356 6636
rect 22652 6690 22708 7308
rect 23324 7364 23380 7374
rect 23324 7270 23380 7308
rect 22988 7250 23044 7262
rect 22988 7198 22990 7250
rect 23042 7198 23044 7250
rect 22988 6804 23044 7198
rect 22988 6738 23044 6748
rect 23100 7252 23156 7262
rect 22652 6638 22654 6690
rect 22706 6638 22708 6690
rect 21624 6300 21888 6310
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21624 6234 21888 6244
rect 20300 5966 20302 6018
rect 20354 5966 20356 6018
rect 20300 5954 20356 5966
rect 19964 5730 20020 5740
rect 22092 5796 22148 5806
rect 22092 5702 22148 5740
rect 11418 5516 11682 5526
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11418 5450 11682 5460
rect 18222 5516 18486 5526
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18222 5450 18486 5460
rect 9884 5292 10164 5348
rect 8540 5124 8596 5134
rect 8016 4732 8280 4742
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8016 4666 8280 4676
rect 4614 3948 4878 3958
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4614 3882 4878 3892
rect 8540 3556 8596 5068
rect 8652 4452 8708 4462
rect 9660 4452 9716 4462
rect 9884 4452 9940 5292
rect 9996 5122 10052 5134
rect 9996 5070 9998 5122
rect 10050 5070 10052 5122
rect 9996 4676 10052 5070
rect 10556 5124 10612 5134
rect 10556 5010 10612 5068
rect 12012 5124 12068 5134
rect 12684 5124 12740 5134
rect 12012 5122 12404 5124
rect 12012 5070 12014 5122
rect 12066 5070 12404 5122
rect 12012 5068 12404 5070
rect 12012 5058 12068 5068
rect 10556 4958 10558 5010
rect 10610 4958 10612 5010
rect 10556 4946 10612 4958
rect 10892 5010 10948 5022
rect 11228 5012 11284 5022
rect 10892 4958 10894 5010
rect 10946 4958 10948 5010
rect 10220 4900 10276 4910
rect 10220 4898 10500 4900
rect 10220 4846 10222 4898
rect 10274 4846 10500 4898
rect 10220 4844 10500 4846
rect 10220 4834 10276 4844
rect 9996 4620 10388 4676
rect 10332 4562 10388 4620
rect 10332 4510 10334 4562
rect 10386 4510 10388 4562
rect 10332 4498 10388 4510
rect 9996 4452 10052 4462
rect 8652 4450 9828 4452
rect 8652 4398 8654 4450
rect 8706 4398 9662 4450
rect 9714 4398 9828 4450
rect 8652 4396 9828 4398
rect 9884 4450 10052 4452
rect 9884 4398 9998 4450
rect 10050 4398 10052 4450
rect 9884 4396 10052 4398
rect 8652 4386 8708 4396
rect 9660 4386 9716 4396
rect 9100 4228 9156 4238
rect 9100 4134 9156 4172
rect 9772 4004 9828 4396
rect 9996 4386 10052 4396
rect 9772 3948 9940 4004
rect 8652 3556 8708 3566
rect 8540 3554 8708 3556
rect 8540 3502 8654 3554
rect 8706 3502 8708 3554
rect 8540 3500 8708 3502
rect 8652 3490 8708 3500
rect 6748 3330 6804 3342
rect 6748 3278 6750 3330
rect 6802 3278 6804 3330
rect 6748 800 6804 3278
rect 7196 3332 7252 3342
rect 7980 3332 8036 3342
rect 7196 3330 7476 3332
rect 7196 3278 7198 3330
rect 7250 3278 7476 3330
rect 7196 3276 7476 3278
rect 7196 3266 7252 3276
rect 7420 800 7476 3276
rect 7868 3330 8036 3332
rect 7868 3278 7982 3330
rect 8034 3278 8036 3330
rect 7868 3276 8036 3278
rect 7868 1988 7924 3276
rect 7980 3266 8036 3276
rect 9772 3330 9828 3342
rect 9772 3278 9774 3330
rect 9826 3278 9828 3330
rect 8016 3164 8280 3174
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8016 3098 8280 3108
rect 7868 1932 8148 1988
rect 8092 800 8148 1932
rect 9772 1652 9828 3278
rect 8764 1596 9828 1652
rect 8764 800 8820 1596
rect 9884 980 9940 3948
rect 10444 3554 10500 4844
rect 10444 3502 10446 3554
rect 10498 3502 10500 3554
rect 10444 3490 10500 3502
rect 10556 4338 10612 4350
rect 10556 4286 10558 4338
rect 10610 4286 10612 4338
rect 10556 4228 10612 4286
rect 10556 3388 10612 4172
rect 10332 3332 10612 3388
rect 10892 3442 10948 4958
rect 10892 3390 10894 3442
rect 10946 3390 10948 3442
rect 10892 3378 10948 3390
rect 11116 5010 11284 5012
rect 11116 4958 11230 5010
rect 11282 4958 11284 5010
rect 11116 4956 11284 4958
rect 11116 3332 11172 4956
rect 11228 4946 11284 4956
rect 11564 4898 11620 4910
rect 11564 4846 11566 4898
rect 11618 4846 11620 4898
rect 11564 4564 11620 4846
rect 12236 4898 12292 4910
rect 12236 4846 12238 4898
rect 12290 4846 12292 4898
rect 12124 4564 12180 4574
rect 11564 4562 12180 4564
rect 11564 4510 12126 4562
rect 12178 4510 12180 4562
rect 11564 4508 12180 4510
rect 12124 4498 12180 4508
rect 12236 4564 12292 4846
rect 12236 4498 12292 4508
rect 11340 4228 11396 4238
rect 10332 980 10388 3332
rect 11116 3266 11172 3276
rect 11228 4226 11396 4228
rect 11228 4174 11342 4226
rect 11394 4174 11396 4226
rect 11228 4172 11396 4174
rect 11228 3554 11284 4172
rect 11340 4162 11396 4172
rect 11788 4226 11844 4238
rect 11788 4174 11790 4226
rect 11842 4174 11844 4226
rect 11418 3948 11682 3958
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11418 3882 11682 3892
rect 11788 3556 11844 4174
rect 11228 3502 11230 3554
rect 11282 3502 11284 3554
rect 11228 1764 11284 3502
rect 9436 924 9940 980
rect 10108 924 10388 980
rect 10780 1708 11284 1764
rect 11452 3554 11844 3556
rect 11452 3502 11790 3554
rect 11842 3502 11844 3554
rect 11452 3500 11844 3502
rect 9436 800 9492 924
rect 10108 800 10164 924
rect 10780 800 10836 1708
rect 11452 800 11508 3500
rect 11788 3490 11844 3500
rect 12236 3444 12292 3454
rect 12348 3444 12404 5068
rect 12684 5030 12740 5068
rect 18060 5124 18116 5134
rect 13468 5010 13524 5022
rect 13468 4958 13470 5010
rect 13522 4958 13524 5010
rect 12908 4900 12964 4910
rect 12908 4806 12964 4844
rect 13468 4452 13524 4958
rect 14476 5012 14532 5022
rect 14476 4918 14532 4956
rect 15260 5012 15316 5022
rect 13468 4386 13524 4396
rect 13580 4900 13636 4910
rect 12796 4226 12852 4238
rect 12796 4174 12798 4226
rect 12850 4174 12852 4226
rect 12572 3444 12628 3482
rect 12684 3444 12740 3454
rect 12236 3442 12404 3444
rect 12236 3390 12238 3442
rect 12290 3390 12404 3442
rect 12236 3388 12404 3390
rect 12460 3442 12684 3444
rect 12460 3390 12574 3442
rect 12626 3390 12684 3442
rect 12460 3388 12684 3390
rect 12236 3378 12292 3388
rect 11564 3332 11620 3342
rect 11564 3238 11620 3276
rect 12460 1764 12516 3388
rect 12572 3378 12628 3388
rect 12684 3378 12740 3388
rect 12124 1708 12516 1764
rect 12124 800 12180 1708
rect 12796 800 12852 4174
rect 13580 3554 13636 4844
rect 13804 4900 13860 4910
rect 14812 4900 14868 4910
rect 13804 4806 13860 4844
rect 14700 4898 14868 4900
rect 14700 4846 14814 4898
rect 14866 4846 14868 4898
rect 14700 4844 14868 4846
rect 13692 4564 13748 4574
rect 13692 4470 13748 4508
rect 14140 4228 14196 4238
rect 13580 3502 13582 3554
rect 13634 3502 13636 3554
rect 13580 3490 13636 3502
rect 13916 4226 14196 4228
rect 13916 4174 14142 4226
rect 14194 4174 14196 4226
rect 13916 4172 14196 4174
rect 13244 3444 13300 3482
rect 13916 3388 13972 4172
rect 14140 4162 14196 4172
rect 14700 3556 14756 4844
rect 14812 4834 14868 4844
rect 15148 4900 15204 4910
rect 14820 4732 15084 4742
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 14820 4666 15084 4676
rect 14700 3490 14756 3500
rect 14924 4340 14980 4350
rect 14924 3388 14980 4284
rect 15148 3554 15204 4844
rect 15260 4562 15316 4956
rect 15260 4510 15262 4562
rect 15314 4510 15316 4562
rect 15260 4498 15316 4510
rect 17836 4898 17892 4910
rect 17836 4846 17838 4898
rect 17890 4846 17892 4898
rect 17388 4452 17444 4462
rect 17388 4358 17444 4396
rect 15596 4340 15652 4350
rect 15596 4246 15652 4284
rect 17612 4338 17668 4350
rect 17612 4286 17614 4338
rect 17666 4286 17668 4338
rect 16828 4228 16884 4238
rect 17612 4228 17668 4286
rect 16828 4226 17668 4228
rect 16828 4174 16830 4226
rect 16882 4174 17668 4226
rect 16828 4172 17668 4174
rect 15596 3668 15652 3678
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3490 15204 3502
rect 15484 3666 15652 3668
rect 15484 3614 15598 3666
rect 15650 3614 15652 3666
rect 15484 3612 15652 3614
rect 13244 3378 13300 3388
rect 13692 3332 13972 3388
rect 14364 3332 14420 3342
rect 13692 980 13748 3332
rect 13468 924 13748 980
rect 14140 3330 14420 3332
rect 14140 3278 14366 3330
rect 14418 3278 14420 3330
rect 14140 3276 14420 3278
rect 13468 800 13524 924
rect 14140 800 14196 3276
rect 14364 3266 14420 3276
rect 14700 3332 14980 3388
rect 14700 1092 14756 3332
rect 14820 3164 15084 3174
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 14820 3098 15084 3108
rect 14700 1036 14868 1092
rect 14812 800 14868 1036
rect 15484 800 15540 3612
rect 15596 3602 15652 3612
rect 16156 3668 16212 3678
rect 16156 800 16212 3612
rect 16828 800 16884 4172
rect 17836 4116 17892 4846
rect 18060 4562 18116 5068
rect 18284 5124 18340 5134
rect 21868 5124 21924 5134
rect 18284 5122 18452 5124
rect 18284 5070 18286 5122
rect 18338 5070 18452 5122
rect 18284 5068 18452 5070
rect 18284 5058 18340 5068
rect 18060 4510 18062 4562
rect 18114 4510 18116 4562
rect 18060 4498 18116 4510
rect 18396 4564 18452 5068
rect 21196 5122 21924 5124
rect 21196 5070 21870 5122
rect 21922 5070 21924 5122
rect 21196 5068 21924 5070
rect 18508 4900 18564 4910
rect 18508 4898 19012 4900
rect 18508 4846 18510 4898
rect 18562 4846 19012 4898
rect 18508 4844 19012 4846
rect 18508 4834 18564 4844
rect 18732 4564 18788 4574
rect 18396 4562 18788 4564
rect 18396 4510 18734 4562
rect 18786 4510 18788 4562
rect 18396 4508 18788 4510
rect 18732 4498 18788 4508
rect 18284 4338 18340 4350
rect 18284 4286 18286 4338
rect 18338 4286 18340 4338
rect 18284 4116 18340 4286
rect 17836 4060 18340 4116
rect 17388 3668 17444 3678
rect 17388 3574 17444 3612
rect 16940 3556 16996 3566
rect 16940 3462 16996 3500
rect 18060 3108 18116 4060
rect 18222 3948 18486 3958
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18222 3882 18486 3892
rect 18956 3554 19012 4844
rect 20748 4898 20804 4910
rect 20748 4846 20750 4898
rect 20802 4846 20804 4898
rect 20748 4676 20804 4846
rect 20300 4620 20804 4676
rect 18956 3502 18958 3554
rect 19010 3502 19012 3554
rect 18956 3490 19012 3502
rect 19068 4338 19124 4350
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 18396 3444 18452 3454
rect 18396 3332 18452 3388
rect 19068 3444 19124 4286
rect 20188 4340 20244 4350
rect 20300 4340 20356 4620
rect 20412 4452 20468 4462
rect 20748 4452 20804 4462
rect 20412 4450 20804 4452
rect 20412 4398 20414 4450
rect 20466 4398 20750 4450
rect 20802 4398 20804 4450
rect 20412 4396 20804 4398
rect 20412 4386 20468 4396
rect 20748 4386 20804 4396
rect 21084 4450 21140 4462
rect 21084 4398 21086 4450
rect 21138 4398 21140 4450
rect 20188 4338 20356 4340
rect 20188 4286 20190 4338
rect 20242 4286 20356 4338
rect 20188 4284 20356 4286
rect 19404 3668 19460 3678
rect 19068 3378 19124 3388
rect 19180 3666 19460 3668
rect 19180 3614 19406 3666
rect 19458 3614 19460 3666
rect 19180 3612 19460 3614
rect 17500 3052 18116 3108
rect 18172 3276 18452 3332
rect 17500 800 17556 3052
rect 18172 800 18228 3276
rect 19180 980 19236 3612
rect 19404 3602 19460 3612
rect 20188 2100 20244 4284
rect 21084 3780 21140 4398
rect 21084 3714 21140 3724
rect 20860 3554 20916 3566
rect 20860 3502 20862 3554
rect 20914 3502 20916 3554
rect 20300 3444 20356 3454
rect 20860 3444 20916 3502
rect 20300 3442 20916 3444
rect 20300 3390 20302 3442
rect 20354 3390 20916 3442
rect 20300 3388 20916 3390
rect 20300 3378 20356 3388
rect 20860 2772 20916 3388
rect 21084 3444 21140 3454
rect 21196 3444 21252 5068
rect 21868 5058 21924 5068
rect 22652 5122 22708 6638
rect 23100 6018 23156 7196
rect 24556 7250 24612 7262
rect 24556 7198 24558 7250
rect 24610 7198 24612 7250
rect 23324 6916 23380 6926
rect 23324 6690 23380 6860
rect 23324 6638 23326 6690
rect 23378 6638 23380 6690
rect 23324 6626 23380 6638
rect 23100 5966 23102 6018
rect 23154 5966 23156 6018
rect 23100 5954 23156 5966
rect 24220 6132 24276 6142
rect 22652 5070 22654 5122
rect 22706 5070 22708 5122
rect 22652 5058 22708 5070
rect 23100 5796 23156 5806
rect 23100 5122 23156 5740
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 23100 5058 23156 5070
rect 23212 5236 23268 5246
rect 21532 4900 21588 4910
rect 21420 4844 21532 4900
rect 21420 3780 21476 4844
rect 21532 4834 21588 4844
rect 22204 4898 22260 4910
rect 22204 4846 22206 4898
rect 22258 4846 22260 4898
rect 21624 4732 21888 4742
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21624 4666 21888 4676
rect 22204 4676 22260 4846
rect 22204 4610 22260 4620
rect 23100 4564 23156 4574
rect 21756 4450 21812 4462
rect 21756 4398 21758 4450
rect 21810 4398 21812 4450
rect 21532 4340 21588 4350
rect 21532 4338 21700 4340
rect 21532 4286 21534 4338
rect 21586 4286 21700 4338
rect 21532 4284 21700 4286
rect 21532 4274 21588 4284
rect 21644 3892 21700 4284
rect 21756 4116 21812 4398
rect 22428 4452 22484 4462
rect 22428 4358 22484 4396
rect 22764 4450 22820 4462
rect 22764 4398 22766 4450
rect 22818 4398 22820 4450
rect 22204 4338 22260 4350
rect 22204 4286 22206 4338
rect 22258 4286 22260 4338
rect 22204 4228 22260 4286
rect 22764 4228 22820 4398
rect 23100 4450 23156 4508
rect 23100 4398 23102 4450
rect 23154 4398 23156 4450
rect 23100 4386 23156 4398
rect 22204 4172 22820 4228
rect 21756 4050 21812 4060
rect 22876 4116 22932 4126
rect 21644 3836 22148 3892
rect 21420 3724 21812 3780
rect 21084 3442 21252 3444
rect 21084 3390 21086 3442
rect 21138 3390 21252 3442
rect 21084 3388 21252 3390
rect 21532 3554 21588 3566
rect 21532 3502 21534 3554
rect 21586 3502 21588 3554
rect 21532 3444 21588 3502
rect 21084 3378 21140 3388
rect 21532 3378 21588 3388
rect 21756 3442 21812 3724
rect 21756 3390 21758 3442
rect 21810 3390 21812 3442
rect 21756 3378 21812 3390
rect 22092 3442 22148 3836
rect 22428 3668 22484 3678
rect 22428 3554 22484 3612
rect 22428 3502 22430 3554
rect 22482 3502 22484 3554
rect 22428 3490 22484 3502
rect 22876 3554 22932 4060
rect 23212 3666 23268 5180
rect 24220 4562 24276 6076
rect 24332 5906 24388 5918
rect 24332 5854 24334 5906
rect 24386 5854 24388 5906
rect 24332 5124 24388 5854
rect 24556 5348 24612 7198
rect 25026 7084 25290 7094
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25026 7018 25290 7028
rect 25676 6692 25732 6702
rect 24668 6020 24724 6030
rect 24668 5926 24724 5964
rect 25026 5516 25290 5526
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25026 5450 25290 5460
rect 24556 5282 24612 5292
rect 25340 5348 25396 5358
rect 24332 5058 24388 5068
rect 25340 5010 25396 5292
rect 25340 4958 25342 5010
rect 25394 4958 25396 5010
rect 25340 4946 25396 4958
rect 24220 4510 24222 4562
rect 24274 4510 24276 4562
rect 24220 4498 24276 4510
rect 24780 4564 24836 4574
rect 24780 4470 24836 4508
rect 23436 4452 23492 4462
rect 23436 4358 23492 4396
rect 23212 3614 23214 3666
rect 23266 3614 23268 3666
rect 23212 3602 23268 3614
rect 24668 4116 24724 4126
rect 24668 3668 24724 4060
rect 25026 3948 25290 3958
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25026 3882 25290 3892
rect 24668 3574 24724 3612
rect 25004 3780 25060 3790
rect 22876 3502 22878 3554
rect 22930 3502 22932 3554
rect 22876 3490 22932 3502
rect 25004 3554 25060 3724
rect 25676 3666 25732 6636
rect 25788 6466 25844 7980
rect 26236 7362 26292 7374
rect 26236 7310 26238 7362
rect 26290 7310 26292 7362
rect 26236 6916 26292 7310
rect 26236 6850 26292 6860
rect 25788 6414 25790 6466
rect 25842 6414 25844 6466
rect 25788 6402 25844 6414
rect 26124 6468 26180 6478
rect 26124 5346 26180 6412
rect 26348 6466 26404 6478
rect 26348 6414 26350 6466
rect 26402 6414 26404 6466
rect 26236 5796 26292 5806
rect 26236 5702 26292 5740
rect 26124 5294 26126 5346
rect 26178 5294 26180 5346
rect 26124 5282 26180 5294
rect 26348 4452 26404 6414
rect 26348 4386 26404 4396
rect 26460 4226 26516 8764
rect 26684 8258 26740 9884
rect 27244 9156 27300 9166
rect 27244 9062 27300 9100
rect 26684 8206 26686 8258
rect 26738 8206 26740 8258
rect 26684 8194 26740 8206
rect 27132 8484 27188 8494
rect 27132 8258 27188 8428
rect 27132 8206 27134 8258
rect 27186 8206 27188 8258
rect 27132 8194 27188 8206
rect 27356 8260 27412 10556
rect 27468 9940 27524 9950
rect 27468 9846 27524 9884
rect 28428 9436 28692 9446
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28428 9370 28692 9380
rect 27692 8820 27748 8830
rect 27468 8260 27524 8270
rect 27356 8258 27524 8260
rect 27356 8206 27470 8258
rect 27522 8206 27524 8258
rect 27356 8204 27524 8206
rect 27468 8148 27524 8204
rect 27468 8082 27524 8092
rect 27580 8036 27636 8046
rect 27580 7942 27636 7980
rect 27244 7588 27300 7598
rect 27244 7494 27300 7532
rect 27356 7476 27412 7486
rect 27244 6804 27300 6814
rect 26908 6468 26964 6478
rect 26908 6374 26964 6412
rect 26908 6020 26964 6030
rect 26908 5122 26964 5964
rect 27244 6018 27300 6748
rect 27244 5966 27246 6018
rect 27298 5966 27300 6018
rect 27244 5954 27300 5966
rect 26908 5070 26910 5122
rect 26962 5070 26964 5122
rect 26908 5058 26964 5070
rect 26572 4900 26628 4910
rect 26572 4898 26740 4900
rect 26572 4846 26574 4898
rect 26626 4846 26740 4898
rect 26572 4844 26740 4846
rect 26572 4834 26628 4844
rect 26460 4174 26462 4226
rect 26514 4174 26516 4226
rect 26460 4162 26516 4174
rect 26572 4676 26628 4686
rect 25676 3614 25678 3666
rect 25730 3614 25732 3666
rect 25676 3602 25732 3614
rect 25004 3502 25006 3554
rect 25058 3502 25060 3554
rect 25004 3490 25060 3502
rect 26572 3554 26628 4620
rect 26572 3502 26574 3554
rect 26626 3502 26628 3554
rect 26572 3490 26628 3502
rect 22092 3390 22094 3442
rect 22146 3390 22148 3442
rect 22092 3378 22148 3390
rect 24108 3444 24164 3454
rect 24108 3350 24164 3388
rect 21624 3164 21888 3174
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21624 3098 21888 3108
rect 20860 2706 20916 2716
rect 20188 2034 20244 2044
rect 26684 1428 26740 4844
rect 27356 3778 27412 7420
rect 27692 6690 27748 8764
rect 28140 8484 28196 8494
rect 27692 6638 27694 6690
rect 27746 6638 27748 6690
rect 27692 6626 27748 6638
rect 27804 8148 27860 8158
rect 27692 5348 27748 5358
rect 27804 5348 27860 8092
rect 27692 5346 27860 5348
rect 27692 5294 27694 5346
rect 27746 5294 27860 5346
rect 27692 5292 27860 5294
rect 28140 7362 28196 8428
rect 28428 7868 28692 7878
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28428 7802 28692 7812
rect 28140 7310 28142 7362
rect 28194 7310 28196 7362
rect 28140 6466 28196 7310
rect 28140 6414 28142 6466
rect 28194 6414 28196 6466
rect 27692 5282 27748 5292
rect 28140 5234 28196 6414
rect 28428 6300 28692 6310
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28428 6234 28692 6244
rect 28140 5182 28142 5234
rect 28194 5182 28196 5234
rect 28140 5170 28196 5182
rect 28428 4732 28692 4742
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28428 4666 28692 4676
rect 27468 4452 27524 4462
rect 27468 4358 27524 4396
rect 27356 3726 27358 3778
rect 27410 3726 27412 3778
rect 27356 3714 27412 3726
rect 28428 3164 28692 3174
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28428 3098 28692 3108
rect 26684 1362 26740 1372
rect 18844 924 19236 980
rect 18844 800 18900 924
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
<< via2 >>
rect 24444 29596 24500 29652
rect 2156 25282 2212 25284
rect 2156 25230 2158 25282
rect 2158 25230 2210 25282
rect 2210 25230 2212 25282
rect 2156 25228 2212 25230
rect 3388 26290 3444 26292
rect 3388 26238 3390 26290
rect 3390 26238 3442 26290
rect 3442 26238 3444 26290
rect 3388 26236 3444 26238
rect 4284 26124 4340 26180
rect 3948 25676 4004 25732
rect 2940 25282 2996 25284
rect 2940 25230 2942 25282
rect 2942 25230 2994 25282
rect 2994 25230 2996 25282
rect 2940 25228 2996 25230
rect 2716 25116 2772 25172
rect 3500 25228 3556 25284
rect 4284 25116 4340 25172
rect 4614 25898 4670 25900
rect 4614 25846 4616 25898
rect 4616 25846 4668 25898
rect 4668 25846 4670 25898
rect 4614 25844 4670 25846
rect 4718 25898 4774 25900
rect 4718 25846 4720 25898
rect 4720 25846 4772 25898
rect 4772 25846 4774 25898
rect 4718 25844 4774 25846
rect 4822 25898 4878 25900
rect 4822 25846 4824 25898
rect 4824 25846 4876 25898
rect 4876 25846 4878 25898
rect 4822 25844 4878 25846
rect 6076 25618 6132 25620
rect 6076 25566 6078 25618
rect 6078 25566 6130 25618
rect 6130 25566 6132 25618
rect 6076 25564 6132 25566
rect 4620 25282 4676 25284
rect 4620 25230 4622 25282
rect 4622 25230 4674 25282
rect 4674 25230 4676 25282
rect 4620 25228 4676 25230
rect 2380 24220 2436 24276
rect 2044 24108 2100 24164
rect 2044 23826 2100 23828
rect 2044 23774 2046 23826
rect 2046 23774 2098 23826
rect 2098 23774 2100 23826
rect 2044 23772 2100 23774
rect 4614 24330 4670 24332
rect 4614 24278 4616 24330
rect 4616 24278 4668 24330
rect 4668 24278 4670 24330
rect 4614 24276 4670 24278
rect 4718 24330 4774 24332
rect 4718 24278 4720 24330
rect 4720 24278 4772 24330
rect 4772 24278 4774 24330
rect 4718 24276 4774 24278
rect 4822 24330 4878 24332
rect 4822 24278 4824 24330
rect 4824 24278 4876 24330
rect 4876 24278 4878 24330
rect 4822 24276 4878 24278
rect 3724 23772 3780 23828
rect 1708 23548 1764 23604
rect 2492 23548 2548 23604
rect 6636 25452 6692 25508
rect 6972 25564 7028 25620
rect 7308 25564 7364 25620
rect 8016 26682 8072 26684
rect 8016 26630 8018 26682
rect 8018 26630 8070 26682
rect 8070 26630 8072 26682
rect 8016 26628 8072 26630
rect 8120 26682 8176 26684
rect 8120 26630 8122 26682
rect 8122 26630 8174 26682
rect 8174 26630 8176 26682
rect 8120 26628 8176 26630
rect 8224 26682 8280 26684
rect 8224 26630 8226 26682
rect 8226 26630 8278 26682
rect 8278 26630 8280 26682
rect 8224 26628 8280 26630
rect 7980 25394 8036 25396
rect 7980 25342 7982 25394
rect 7982 25342 8034 25394
rect 8034 25342 8036 25394
rect 7980 25340 8036 25342
rect 8428 25228 8484 25284
rect 8016 25114 8072 25116
rect 8016 25062 8018 25114
rect 8018 25062 8070 25114
rect 8070 25062 8072 25114
rect 8016 25060 8072 25062
rect 8120 25114 8176 25116
rect 8120 25062 8122 25114
rect 8122 25062 8174 25114
rect 8174 25062 8176 25114
rect 8120 25060 8176 25062
rect 8224 25114 8280 25116
rect 8224 25062 8226 25114
rect 8226 25062 8278 25114
rect 8278 25062 8280 25114
rect 8224 25060 8280 25062
rect 6860 23772 6916 23828
rect 9212 25676 9268 25732
rect 8876 24780 8932 24836
rect 9324 25282 9380 25284
rect 9324 25230 9326 25282
rect 9326 25230 9378 25282
rect 9378 25230 9380 25282
rect 9324 25228 9380 25230
rect 9436 24892 9492 24948
rect 9548 26236 9604 26292
rect 8016 23546 8072 23548
rect 8016 23494 8018 23546
rect 8018 23494 8070 23546
rect 8070 23494 8072 23546
rect 8016 23492 8072 23494
rect 8120 23546 8176 23548
rect 8120 23494 8122 23546
rect 8122 23494 8174 23546
rect 8174 23494 8176 23546
rect 8120 23492 8176 23494
rect 8224 23546 8280 23548
rect 8224 23494 8226 23546
rect 8226 23494 8278 23546
rect 8278 23494 8280 23546
rect 8224 23492 8280 23494
rect 9772 25452 9828 25508
rect 9660 24834 9716 24836
rect 9660 24782 9662 24834
rect 9662 24782 9714 24834
rect 9714 24782 9716 24834
rect 9660 24780 9716 24782
rect 9660 24108 9716 24164
rect 4956 23212 5012 23268
rect 9996 25452 10052 25508
rect 10668 26124 10724 26180
rect 10444 24946 10500 24948
rect 10444 24894 10446 24946
rect 10446 24894 10498 24946
rect 10498 24894 10500 24946
rect 10444 24892 10500 24894
rect 10780 25564 10836 25620
rect 10556 23436 10612 23492
rect 10220 23266 10276 23268
rect 10220 23214 10222 23266
rect 10222 23214 10274 23266
rect 10274 23214 10276 23266
rect 10220 23212 10276 23214
rect 11004 25004 11060 25060
rect 10892 24444 10948 24500
rect 11452 26012 11508 26068
rect 12124 26012 12180 26068
rect 11418 25898 11474 25900
rect 11418 25846 11420 25898
rect 11420 25846 11472 25898
rect 11472 25846 11474 25898
rect 11418 25844 11474 25846
rect 11522 25898 11578 25900
rect 11522 25846 11524 25898
rect 11524 25846 11576 25898
rect 11576 25846 11578 25898
rect 11522 25844 11578 25846
rect 11626 25898 11682 25900
rect 11626 25846 11628 25898
rect 11628 25846 11680 25898
rect 11680 25846 11682 25898
rect 11626 25844 11682 25846
rect 12796 25676 12852 25732
rect 11788 25506 11844 25508
rect 11788 25454 11790 25506
rect 11790 25454 11842 25506
rect 11842 25454 11844 25506
rect 11788 25452 11844 25454
rect 11900 25340 11956 25396
rect 11340 24444 11396 24500
rect 11418 24330 11474 24332
rect 11418 24278 11420 24330
rect 11420 24278 11472 24330
rect 11472 24278 11474 24330
rect 11418 24276 11474 24278
rect 11522 24330 11578 24332
rect 11522 24278 11524 24330
rect 11524 24278 11576 24330
rect 11576 24278 11578 24330
rect 11522 24276 11578 24278
rect 11626 24330 11682 24332
rect 11626 24278 11628 24330
rect 11628 24278 11680 24330
rect 11680 24278 11682 24330
rect 11626 24276 11682 24278
rect 11676 23826 11732 23828
rect 11676 23774 11678 23826
rect 11678 23774 11730 23826
rect 11730 23774 11732 23826
rect 11676 23772 11732 23774
rect 13916 25676 13972 25732
rect 14820 26682 14876 26684
rect 14820 26630 14822 26682
rect 14822 26630 14874 26682
rect 14874 26630 14876 26682
rect 14820 26628 14876 26630
rect 14924 26682 14980 26684
rect 14924 26630 14926 26682
rect 14926 26630 14978 26682
rect 14978 26630 14980 26682
rect 14924 26628 14980 26630
rect 15028 26682 15084 26684
rect 15028 26630 15030 26682
rect 15030 26630 15082 26682
rect 15082 26630 15084 26682
rect 15028 26628 15084 26630
rect 16156 26460 16212 26516
rect 15932 25788 15988 25844
rect 14820 25114 14876 25116
rect 14820 25062 14822 25114
rect 14822 25062 14874 25114
rect 14874 25062 14876 25114
rect 14820 25060 14876 25062
rect 14924 25114 14980 25116
rect 14924 25062 14926 25114
rect 14926 25062 14978 25114
rect 14978 25062 14980 25114
rect 14924 25060 14980 25062
rect 15028 25114 15084 25116
rect 15028 25062 15030 25114
rect 15030 25062 15082 25114
rect 15082 25062 15084 25114
rect 15028 25060 15084 25062
rect 15260 25228 15316 25284
rect 17500 26796 17556 26852
rect 18956 26796 19012 26852
rect 18172 26572 18228 26628
rect 18844 26572 18900 26628
rect 17388 26460 17444 26516
rect 16940 25788 16996 25844
rect 18222 25898 18278 25900
rect 18222 25846 18224 25898
rect 18224 25846 18276 25898
rect 18276 25846 18278 25898
rect 18222 25844 18278 25846
rect 18326 25898 18382 25900
rect 18326 25846 18328 25898
rect 18328 25846 18380 25898
rect 18380 25846 18382 25898
rect 18326 25844 18382 25846
rect 18430 25898 18486 25900
rect 18430 25846 18432 25898
rect 18432 25846 18484 25898
rect 18484 25846 18486 25898
rect 18430 25844 18486 25846
rect 18508 25506 18564 25508
rect 18508 25454 18510 25506
rect 18510 25454 18562 25506
rect 18562 25454 18564 25506
rect 18508 25452 18564 25454
rect 16828 25340 16884 25396
rect 16492 25228 16548 25284
rect 19628 25618 19684 25620
rect 19628 25566 19630 25618
rect 19630 25566 19682 25618
rect 19682 25566 19684 25618
rect 19628 25564 19684 25566
rect 18620 25340 18676 25396
rect 17052 25282 17108 25284
rect 17052 25230 17054 25282
rect 17054 25230 17106 25282
rect 17106 25230 17108 25282
rect 17052 25228 17108 25230
rect 18222 24330 18278 24332
rect 18222 24278 18224 24330
rect 18224 24278 18276 24330
rect 18276 24278 18278 24330
rect 18222 24276 18278 24278
rect 18326 24330 18382 24332
rect 18326 24278 18328 24330
rect 18328 24278 18380 24330
rect 18380 24278 18382 24330
rect 18326 24276 18382 24278
rect 18430 24330 18486 24332
rect 18430 24278 18432 24330
rect 18432 24278 18484 24330
rect 18484 24278 18486 24330
rect 18430 24276 18486 24278
rect 20188 25564 20244 25620
rect 21532 26796 21588 26852
rect 22764 26796 22820 26852
rect 21624 26682 21680 26684
rect 21624 26630 21626 26682
rect 21626 26630 21678 26682
rect 21678 26630 21680 26682
rect 21624 26628 21680 26630
rect 21728 26682 21784 26684
rect 21728 26630 21730 26682
rect 21730 26630 21782 26682
rect 21782 26630 21784 26682
rect 21728 26628 21784 26630
rect 21832 26682 21888 26684
rect 21832 26630 21834 26682
rect 21834 26630 21886 26682
rect 21886 26630 21888 26682
rect 21832 26628 21888 26630
rect 20748 25340 20804 25396
rect 20524 25228 20580 25284
rect 20860 24668 20916 24724
rect 13356 23436 13412 23492
rect 14820 23546 14876 23548
rect 14820 23494 14822 23546
rect 14822 23494 14874 23546
rect 14874 23494 14876 23546
rect 14820 23492 14876 23494
rect 14924 23546 14980 23548
rect 14924 23494 14926 23546
rect 14926 23494 14978 23546
rect 14978 23494 14980 23546
rect 14924 23492 14980 23494
rect 15028 23546 15084 23548
rect 15028 23494 15030 23546
rect 15030 23494 15082 23546
rect 15082 23494 15084 23546
rect 15028 23492 15084 23494
rect 21624 25114 21680 25116
rect 21624 25062 21626 25114
rect 21626 25062 21678 25114
rect 21678 25062 21680 25114
rect 21624 25060 21680 25062
rect 21728 25114 21784 25116
rect 21728 25062 21730 25114
rect 21730 25062 21782 25114
rect 21782 25062 21784 25114
rect 21728 25060 21784 25062
rect 21832 25114 21888 25116
rect 21832 25062 21834 25114
rect 21834 25062 21886 25114
rect 21886 25062 21888 25114
rect 21832 25060 21888 25062
rect 22988 26796 23044 26852
rect 23996 25282 24052 25284
rect 23996 25230 23998 25282
rect 23998 25230 24050 25282
rect 24050 25230 24052 25282
rect 23996 25228 24052 25230
rect 22540 24668 22596 24724
rect 23100 25116 23156 25172
rect 23660 25116 23716 25172
rect 22764 24610 22820 24612
rect 22764 24558 22766 24610
rect 22766 24558 22818 24610
rect 22818 24558 22820 24610
rect 22764 24556 22820 24558
rect 27804 28924 27860 28980
rect 25116 28252 25172 28308
rect 24892 26460 24948 26516
rect 25004 26796 25060 26852
rect 27468 27580 27524 27636
rect 25900 26908 25956 26964
rect 25026 25898 25082 25900
rect 25026 25846 25028 25898
rect 25028 25846 25080 25898
rect 25080 25846 25082 25898
rect 25026 25844 25082 25846
rect 25130 25898 25186 25900
rect 25130 25846 25132 25898
rect 25132 25846 25184 25898
rect 25184 25846 25186 25898
rect 25130 25844 25186 25846
rect 25234 25898 25290 25900
rect 25234 25846 25236 25898
rect 25236 25846 25288 25898
rect 25288 25846 25290 25898
rect 25234 25844 25290 25846
rect 24556 25340 24612 25396
rect 24668 25282 24724 25284
rect 24668 25230 24670 25282
rect 24670 25230 24722 25282
rect 24722 25230 24724 25282
rect 24668 25228 24724 25230
rect 24444 25116 24500 25172
rect 23772 24892 23828 24948
rect 23996 24834 24052 24836
rect 23996 24782 23998 24834
rect 23998 24782 24050 24834
rect 24050 24782 24052 24834
rect 23996 24780 24052 24782
rect 23324 23884 23380 23940
rect 24668 24556 24724 24612
rect 24220 24108 24276 24164
rect 21624 23546 21680 23548
rect 21624 23494 21626 23546
rect 21626 23494 21678 23546
rect 21678 23494 21680 23546
rect 21624 23492 21680 23494
rect 21728 23546 21784 23548
rect 21728 23494 21730 23546
rect 21730 23494 21782 23546
rect 21782 23494 21784 23546
rect 21728 23492 21784 23494
rect 21832 23546 21888 23548
rect 21832 23494 21834 23546
rect 21834 23494 21886 23546
rect 21886 23494 21888 23546
rect 21832 23492 21888 23494
rect 20636 23212 20692 23268
rect 4614 22762 4670 22764
rect 4614 22710 4616 22762
rect 4616 22710 4668 22762
rect 4668 22710 4670 22762
rect 4614 22708 4670 22710
rect 4718 22762 4774 22764
rect 4718 22710 4720 22762
rect 4720 22710 4772 22762
rect 4772 22710 4774 22762
rect 4718 22708 4774 22710
rect 4822 22762 4878 22764
rect 4822 22710 4824 22762
rect 4824 22710 4876 22762
rect 4876 22710 4878 22762
rect 4822 22708 4878 22710
rect 11418 22762 11474 22764
rect 11418 22710 11420 22762
rect 11420 22710 11472 22762
rect 11472 22710 11474 22762
rect 11418 22708 11474 22710
rect 11522 22762 11578 22764
rect 11522 22710 11524 22762
rect 11524 22710 11576 22762
rect 11576 22710 11578 22762
rect 11522 22708 11578 22710
rect 11626 22762 11682 22764
rect 11626 22710 11628 22762
rect 11628 22710 11680 22762
rect 11680 22710 11682 22762
rect 11626 22708 11682 22710
rect 18222 22762 18278 22764
rect 18222 22710 18224 22762
rect 18224 22710 18276 22762
rect 18276 22710 18278 22762
rect 18222 22708 18278 22710
rect 18326 22762 18382 22764
rect 18326 22710 18328 22762
rect 18328 22710 18380 22762
rect 18380 22710 18382 22762
rect 18326 22708 18382 22710
rect 18430 22762 18486 22764
rect 18430 22710 18432 22762
rect 18432 22710 18484 22762
rect 18484 22710 18486 22762
rect 18430 22708 18486 22710
rect 8016 21978 8072 21980
rect 8016 21926 8018 21978
rect 8018 21926 8070 21978
rect 8070 21926 8072 21978
rect 8016 21924 8072 21926
rect 8120 21978 8176 21980
rect 8120 21926 8122 21978
rect 8122 21926 8174 21978
rect 8174 21926 8176 21978
rect 8120 21924 8176 21926
rect 8224 21978 8280 21980
rect 8224 21926 8226 21978
rect 8226 21926 8278 21978
rect 8278 21926 8280 21978
rect 8224 21924 8280 21926
rect 14820 21978 14876 21980
rect 14820 21926 14822 21978
rect 14822 21926 14874 21978
rect 14874 21926 14876 21978
rect 14820 21924 14876 21926
rect 14924 21978 14980 21980
rect 14924 21926 14926 21978
rect 14926 21926 14978 21978
rect 14978 21926 14980 21978
rect 14924 21924 14980 21926
rect 15028 21978 15084 21980
rect 15028 21926 15030 21978
rect 15030 21926 15082 21978
rect 15082 21926 15084 21978
rect 15028 21924 15084 21926
rect 21624 21978 21680 21980
rect 21624 21926 21626 21978
rect 21626 21926 21678 21978
rect 21678 21926 21680 21978
rect 21624 21924 21680 21926
rect 21728 21978 21784 21980
rect 21728 21926 21730 21978
rect 21730 21926 21782 21978
rect 21782 21926 21784 21978
rect 21728 21924 21784 21926
rect 21832 21978 21888 21980
rect 21832 21926 21834 21978
rect 21834 21926 21886 21978
rect 21886 21926 21888 21978
rect 21832 21924 21888 21926
rect 13020 21644 13076 21700
rect 12348 21420 12404 21476
rect 4614 21194 4670 21196
rect 4614 21142 4616 21194
rect 4616 21142 4668 21194
rect 4668 21142 4670 21194
rect 4614 21140 4670 21142
rect 4718 21194 4774 21196
rect 4718 21142 4720 21194
rect 4720 21142 4772 21194
rect 4772 21142 4774 21194
rect 4718 21140 4774 21142
rect 4822 21194 4878 21196
rect 4822 21142 4824 21194
rect 4824 21142 4876 21194
rect 4876 21142 4878 21194
rect 4822 21140 4878 21142
rect 11418 21194 11474 21196
rect 11418 21142 11420 21194
rect 11420 21142 11472 21194
rect 11472 21142 11474 21194
rect 11418 21140 11474 21142
rect 11522 21194 11578 21196
rect 11522 21142 11524 21194
rect 11524 21142 11576 21194
rect 11576 21142 11578 21194
rect 11522 21140 11578 21142
rect 11626 21194 11682 21196
rect 11626 21142 11628 21194
rect 11628 21142 11680 21194
rect 11680 21142 11682 21194
rect 11626 21140 11682 21142
rect 8016 20410 8072 20412
rect 8016 20358 8018 20410
rect 8018 20358 8070 20410
rect 8070 20358 8072 20410
rect 8016 20356 8072 20358
rect 8120 20410 8176 20412
rect 8120 20358 8122 20410
rect 8122 20358 8174 20410
rect 8174 20358 8176 20410
rect 8120 20356 8176 20358
rect 8224 20410 8280 20412
rect 8224 20358 8226 20410
rect 8226 20358 8278 20410
rect 8278 20358 8280 20410
rect 8224 20356 8280 20358
rect 8540 19740 8596 19796
rect 4614 19626 4670 19628
rect 4284 19516 4340 19572
rect 4614 19574 4616 19626
rect 4616 19574 4668 19626
rect 4668 19574 4670 19626
rect 4614 19572 4670 19574
rect 4718 19626 4774 19628
rect 4718 19574 4720 19626
rect 4720 19574 4772 19626
rect 4772 19574 4774 19626
rect 4718 19572 4774 19574
rect 4822 19626 4878 19628
rect 4822 19574 4824 19626
rect 4824 19574 4876 19626
rect 4876 19574 4878 19626
rect 4822 19572 4878 19574
rect 1596 16658 1652 16660
rect 1596 16606 1598 16658
rect 1598 16606 1650 16658
rect 1650 16606 1652 16658
rect 1596 16604 1652 16606
rect 3612 16828 3668 16884
rect 2716 16604 2772 16660
rect 2044 14252 2100 14308
rect 3948 16604 4004 16660
rect 3052 14418 3108 14420
rect 3052 14366 3054 14418
rect 3054 14366 3106 14418
rect 3106 14366 3108 14418
rect 3052 14364 3108 14366
rect 2716 14252 2772 14308
rect 3388 14252 3444 14308
rect 1596 11228 1652 11284
rect 1820 10834 1876 10836
rect 1820 10782 1822 10834
rect 1822 10782 1874 10834
rect 1874 10782 1876 10834
rect 1820 10780 1876 10782
rect 4060 13692 4116 13748
rect 6076 19292 6132 19348
rect 4614 18058 4670 18060
rect 4614 18006 4616 18058
rect 4616 18006 4668 18058
rect 4668 18006 4670 18058
rect 4614 18004 4670 18006
rect 4718 18058 4774 18060
rect 4718 18006 4720 18058
rect 4720 18006 4772 18058
rect 4772 18006 4774 18058
rect 4718 18004 4774 18006
rect 4822 18058 4878 18060
rect 4822 18006 4824 18058
rect 4824 18006 4876 18058
rect 4876 18006 4878 18058
rect 4822 18004 4878 18006
rect 7644 19346 7700 19348
rect 7644 19294 7646 19346
rect 7646 19294 7698 19346
rect 7698 19294 7700 19346
rect 7644 19292 7700 19294
rect 8016 18842 8072 18844
rect 8016 18790 8018 18842
rect 8018 18790 8070 18842
rect 8070 18790 8072 18842
rect 8016 18788 8072 18790
rect 8120 18842 8176 18844
rect 8120 18790 8122 18842
rect 8122 18790 8174 18842
rect 8174 18790 8176 18842
rect 8120 18788 8176 18790
rect 8224 18842 8280 18844
rect 8224 18790 8226 18842
rect 8226 18790 8278 18842
rect 8278 18790 8280 18842
rect 8224 18788 8280 18790
rect 9548 19794 9604 19796
rect 9548 19742 9550 19794
rect 9550 19742 9602 19794
rect 9602 19742 9604 19794
rect 9548 19740 9604 19742
rect 5516 17612 5572 17668
rect 4956 17442 5012 17444
rect 4956 17390 4958 17442
rect 4958 17390 5010 17442
rect 5010 17390 5012 17442
rect 4956 17388 5012 17390
rect 4284 12908 4340 12964
rect 4614 16490 4670 16492
rect 4614 16438 4616 16490
rect 4616 16438 4668 16490
rect 4668 16438 4670 16490
rect 4614 16436 4670 16438
rect 4718 16490 4774 16492
rect 4718 16438 4720 16490
rect 4720 16438 4772 16490
rect 4772 16438 4774 16490
rect 4718 16436 4774 16438
rect 4822 16490 4878 16492
rect 4822 16438 4824 16490
rect 4824 16438 4876 16490
rect 4876 16438 4878 16490
rect 4822 16436 4878 16438
rect 4614 14922 4670 14924
rect 4614 14870 4616 14922
rect 4616 14870 4668 14922
rect 4668 14870 4670 14922
rect 4614 14868 4670 14870
rect 4718 14922 4774 14924
rect 4718 14870 4720 14922
rect 4720 14870 4772 14922
rect 4772 14870 4774 14922
rect 4718 14868 4774 14870
rect 4822 14922 4878 14924
rect 4822 14870 4824 14922
rect 4824 14870 4876 14922
rect 4876 14870 4878 14922
rect 4822 14868 4878 14870
rect 5068 16882 5124 16884
rect 5068 16830 5070 16882
rect 5070 16830 5122 16882
rect 5122 16830 5124 16882
rect 5068 16828 5124 16830
rect 7532 17666 7588 17668
rect 7532 17614 7534 17666
rect 7534 17614 7586 17666
rect 7586 17614 7588 17666
rect 7532 17612 7588 17614
rect 5628 17388 5684 17444
rect 5516 16882 5572 16884
rect 5516 16830 5518 16882
rect 5518 16830 5570 16882
rect 5570 16830 5572 16882
rect 5516 16828 5572 16830
rect 5852 16604 5908 16660
rect 6076 16156 6132 16212
rect 6636 17442 6692 17444
rect 6636 17390 6638 17442
rect 6638 17390 6690 17442
rect 6690 17390 6692 17442
rect 6636 17388 6692 17390
rect 8016 17274 8072 17276
rect 8016 17222 8018 17274
rect 8018 17222 8070 17274
rect 8070 17222 8072 17274
rect 8016 17220 8072 17222
rect 8120 17274 8176 17276
rect 8120 17222 8122 17274
rect 8122 17222 8174 17274
rect 8174 17222 8176 17274
rect 8120 17220 8176 17222
rect 8224 17274 8280 17276
rect 8224 17222 8226 17274
rect 8226 17222 8278 17274
rect 8278 17222 8280 17274
rect 8224 17220 8280 17222
rect 6972 16210 7028 16212
rect 6972 16158 6974 16210
rect 6974 16158 7026 16210
rect 7026 16158 7028 16210
rect 6972 16156 7028 16158
rect 9548 18396 9604 18452
rect 8428 16716 8484 16772
rect 8016 15706 8072 15708
rect 8016 15654 8018 15706
rect 8018 15654 8070 15706
rect 8070 15654 8072 15706
rect 8016 15652 8072 15654
rect 8120 15706 8176 15708
rect 8120 15654 8122 15706
rect 8122 15654 8174 15706
rect 8174 15654 8176 15706
rect 8120 15652 8176 15654
rect 8224 15706 8280 15708
rect 8224 15654 8226 15706
rect 8226 15654 8278 15706
rect 8278 15654 8280 15706
rect 8224 15652 8280 15654
rect 9212 15932 9268 15988
rect 9548 17612 9604 17668
rect 11418 19626 11474 19628
rect 11418 19574 11420 19626
rect 11420 19574 11472 19626
rect 11472 19574 11474 19626
rect 11418 19572 11474 19574
rect 11522 19626 11578 19628
rect 11522 19574 11524 19626
rect 11524 19574 11576 19626
rect 11576 19574 11578 19626
rect 11522 19572 11578 19574
rect 11626 19626 11682 19628
rect 11626 19574 11628 19626
rect 11628 19574 11680 19626
rect 11680 19574 11682 19626
rect 11626 19572 11682 19574
rect 9996 18284 10052 18340
rect 11228 18508 11284 18564
rect 9996 17612 10052 17668
rect 14812 21698 14868 21700
rect 14812 21646 14814 21698
rect 14814 21646 14866 21698
rect 14866 21646 14868 21698
rect 14812 21644 14868 21646
rect 24444 21644 24500 21700
rect 13804 21474 13860 21476
rect 13804 21422 13806 21474
rect 13806 21422 13858 21474
rect 13858 21422 13860 21474
rect 13804 21420 13860 21422
rect 18222 21194 18278 21196
rect 18222 21142 18224 21194
rect 18224 21142 18276 21194
rect 18276 21142 18278 21194
rect 18222 21140 18278 21142
rect 18326 21194 18382 21196
rect 18326 21142 18328 21194
rect 18328 21142 18380 21194
rect 18380 21142 18382 21194
rect 18326 21140 18382 21142
rect 18430 21194 18486 21196
rect 18430 21142 18432 21194
rect 18432 21142 18484 21194
rect 18484 21142 18486 21194
rect 18430 21140 18486 21142
rect 15372 20636 15428 20692
rect 14820 20410 14876 20412
rect 14820 20358 14822 20410
rect 14822 20358 14874 20410
rect 14874 20358 14876 20410
rect 14820 20356 14876 20358
rect 14924 20410 14980 20412
rect 14924 20358 14926 20410
rect 14926 20358 14978 20410
rect 14978 20358 14980 20410
rect 14924 20356 14980 20358
rect 15028 20410 15084 20412
rect 15028 20358 15030 20410
rect 15030 20358 15082 20410
rect 15082 20358 15084 20410
rect 15028 20356 15084 20358
rect 14924 20188 14980 20244
rect 11900 18396 11956 18452
rect 11564 18338 11620 18340
rect 11564 18286 11566 18338
rect 11566 18286 11618 18338
rect 11618 18286 11620 18338
rect 11564 18284 11620 18286
rect 11418 18058 11474 18060
rect 11418 18006 11420 18058
rect 11420 18006 11472 18058
rect 11472 18006 11474 18058
rect 11418 18004 11474 18006
rect 11522 18058 11578 18060
rect 11522 18006 11524 18058
rect 11524 18006 11576 18058
rect 11576 18006 11578 18058
rect 11522 18004 11578 18006
rect 11626 18058 11682 18060
rect 11626 18006 11628 18058
rect 11628 18006 11680 18058
rect 11680 18006 11682 18058
rect 11626 18004 11682 18006
rect 12572 18562 12628 18564
rect 12572 18510 12574 18562
rect 12574 18510 12626 18562
rect 12626 18510 12628 18562
rect 12572 18508 12628 18510
rect 12460 18396 12516 18452
rect 11676 17666 11732 17668
rect 11676 17614 11678 17666
rect 11678 17614 11730 17666
rect 11730 17614 11732 17666
rect 11676 17612 11732 17614
rect 8988 15314 9044 15316
rect 8988 15262 8990 15314
rect 8990 15262 9042 15314
rect 9042 15262 9044 15314
rect 8988 15260 9044 15262
rect 5516 14418 5572 14420
rect 5516 14366 5518 14418
rect 5518 14366 5570 14418
rect 5570 14366 5572 14418
rect 5516 14364 5572 14366
rect 4508 14306 4564 14308
rect 4508 14254 4510 14306
rect 4510 14254 4562 14306
rect 4562 14254 4564 14306
rect 4508 14252 4564 14254
rect 8652 14588 8708 14644
rect 9772 16716 9828 16772
rect 11418 16490 11474 16492
rect 11418 16438 11420 16490
rect 11420 16438 11472 16490
rect 11472 16438 11474 16490
rect 11418 16436 11474 16438
rect 11522 16490 11578 16492
rect 11522 16438 11524 16490
rect 11524 16438 11576 16490
rect 11576 16438 11578 16490
rect 11522 16436 11578 16438
rect 11626 16490 11682 16492
rect 11626 16438 11628 16490
rect 11628 16438 11680 16490
rect 11680 16438 11682 16490
rect 11626 16436 11682 16438
rect 10780 15986 10836 15988
rect 10780 15934 10782 15986
rect 10782 15934 10834 15986
rect 10834 15934 10836 15986
rect 10780 15932 10836 15934
rect 11452 15314 11508 15316
rect 11452 15262 11454 15314
rect 11454 15262 11506 15314
rect 11506 15262 11508 15314
rect 11452 15260 11508 15262
rect 12012 15932 12068 15988
rect 13244 18450 13300 18452
rect 13244 18398 13246 18450
rect 13246 18398 13298 18450
rect 13298 18398 13300 18450
rect 13244 18396 13300 18398
rect 22876 20860 22932 20916
rect 17276 20690 17332 20692
rect 17276 20638 17278 20690
rect 17278 20638 17330 20690
rect 17330 20638 17332 20690
rect 17276 20636 17332 20638
rect 21624 20410 21680 20412
rect 21624 20358 21626 20410
rect 21626 20358 21678 20410
rect 21678 20358 21680 20410
rect 21624 20356 21680 20358
rect 21728 20410 21784 20412
rect 21728 20358 21730 20410
rect 21730 20358 21782 20410
rect 21782 20358 21784 20410
rect 21728 20356 21784 20358
rect 21832 20410 21888 20412
rect 21832 20358 21834 20410
rect 21834 20358 21886 20410
rect 21886 20358 21888 20410
rect 21832 20356 21888 20358
rect 16268 20188 16324 20244
rect 14820 18842 14876 18844
rect 14820 18790 14822 18842
rect 14822 18790 14874 18842
rect 14874 18790 14876 18842
rect 14820 18788 14876 18790
rect 14924 18842 14980 18844
rect 14924 18790 14926 18842
rect 14926 18790 14978 18842
rect 14978 18790 14980 18842
rect 14924 18788 14980 18790
rect 15028 18842 15084 18844
rect 15028 18790 15030 18842
rect 15030 18790 15082 18842
rect 15082 18790 15084 18842
rect 15028 18788 15084 18790
rect 14252 18508 14308 18564
rect 13468 17612 13524 17668
rect 12796 17388 12852 17444
rect 13804 17442 13860 17444
rect 13804 17390 13806 17442
rect 13806 17390 13858 17442
rect 13858 17390 13860 17442
rect 13804 17388 13860 17390
rect 16380 19068 16436 19124
rect 17164 19122 17220 19124
rect 17164 19070 17166 19122
rect 17166 19070 17218 19122
rect 17218 19070 17220 19122
rect 17164 19068 17220 19070
rect 16940 18508 16996 18564
rect 16940 18172 16996 18228
rect 15708 17666 15764 17668
rect 15708 17614 15710 17666
rect 15710 17614 15762 17666
rect 15762 17614 15764 17666
rect 15708 17612 15764 17614
rect 13580 15986 13636 15988
rect 13580 15934 13582 15986
rect 13582 15934 13634 15986
rect 13634 15934 13636 15986
rect 13580 15932 13636 15934
rect 8016 14138 8072 14140
rect 8016 14086 8018 14138
rect 8018 14086 8070 14138
rect 8070 14086 8072 14138
rect 8016 14084 8072 14086
rect 8120 14138 8176 14140
rect 8120 14086 8122 14138
rect 8122 14086 8174 14138
rect 8174 14086 8176 14138
rect 8120 14084 8176 14086
rect 8224 14138 8280 14140
rect 8224 14086 8226 14138
rect 8226 14086 8278 14138
rect 8278 14086 8280 14138
rect 8224 14084 8280 14086
rect 7980 13916 8036 13972
rect 5068 13746 5124 13748
rect 5068 13694 5070 13746
rect 5070 13694 5122 13746
rect 5122 13694 5124 13746
rect 5068 13692 5124 13694
rect 4614 13354 4670 13356
rect 4614 13302 4616 13354
rect 4616 13302 4668 13354
rect 4668 13302 4670 13354
rect 4614 13300 4670 13302
rect 4718 13354 4774 13356
rect 4718 13302 4720 13354
rect 4720 13302 4772 13354
rect 4772 13302 4774 13354
rect 4718 13300 4774 13302
rect 4822 13354 4878 13356
rect 4822 13302 4824 13354
rect 4824 13302 4876 13354
rect 4876 13302 4878 13354
rect 4822 13300 4878 13302
rect 5628 12348 5684 12404
rect 3388 11340 3444 11396
rect 2716 11282 2772 11284
rect 2716 11230 2718 11282
rect 2718 11230 2770 11282
rect 2770 11230 2772 11282
rect 2716 11228 2772 11230
rect 2380 10332 2436 10388
rect 2716 10556 2772 10612
rect 3276 10444 3332 10500
rect 3388 10444 3444 10500
rect 5292 12012 5348 12068
rect 4614 11786 4670 11788
rect 4614 11734 4616 11786
rect 4616 11734 4668 11786
rect 4668 11734 4670 11786
rect 4614 11732 4670 11734
rect 4718 11786 4774 11788
rect 4718 11734 4720 11786
rect 4720 11734 4772 11786
rect 4772 11734 4774 11786
rect 4718 11732 4774 11734
rect 4822 11786 4878 11788
rect 4822 11734 4824 11786
rect 4824 11734 4876 11786
rect 4876 11734 4878 11786
rect 4822 11732 4878 11734
rect 4284 10610 4340 10612
rect 4284 10558 4286 10610
rect 4286 10558 4338 10610
rect 4338 10558 4340 10610
rect 4284 10556 4340 10558
rect 9884 13916 9940 13972
rect 9884 13468 9940 13524
rect 6972 13132 7028 13188
rect 9100 13186 9156 13188
rect 9100 13134 9102 13186
rect 9102 13134 9154 13186
rect 9154 13134 9156 13186
rect 9100 13132 9156 13134
rect 6524 12348 6580 12404
rect 5740 12012 5796 12068
rect 7756 12012 7812 12068
rect 6188 10780 6244 10836
rect 6300 11394 6356 11396
rect 6300 11342 6302 11394
rect 6302 11342 6354 11394
rect 6354 11342 6356 11394
rect 6300 11340 6356 11342
rect 4396 10332 4452 10388
rect 4614 10218 4670 10220
rect 4614 10166 4616 10218
rect 4616 10166 4668 10218
rect 4668 10166 4670 10218
rect 4614 10164 4670 10166
rect 4718 10218 4774 10220
rect 4718 10166 4720 10218
rect 4720 10166 4772 10218
rect 4772 10166 4774 10218
rect 4718 10164 4774 10166
rect 4822 10218 4878 10220
rect 4822 10166 4824 10218
rect 4824 10166 4876 10218
rect 4876 10166 4878 10218
rect 4822 10164 4878 10166
rect 5292 10556 5348 10612
rect 7308 11394 7364 11396
rect 7308 11342 7310 11394
rect 7310 11342 7362 11394
rect 7362 11342 7364 11394
rect 7308 11340 7364 11342
rect 8016 12570 8072 12572
rect 8016 12518 8018 12570
rect 8018 12518 8070 12570
rect 8070 12518 8072 12570
rect 8016 12516 8072 12518
rect 8120 12570 8176 12572
rect 8120 12518 8122 12570
rect 8122 12518 8174 12570
rect 8174 12518 8176 12570
rect 8120 12516 8176 12518
rect 8224 12570 8280 12572
rect 8224 12518 8226 12570
rect 8226 12518 8278 12570
rect 8278 12518 8280 12570
rect 8224 12516 8280 12518
rect 8016 11002 8072 11004
rect 8016 10950 8018 11002
rect 8018 10950 8070 11002
rect 8070 10950 8072 11002
rect 8016 10948 8072 10950
rect 8120 11002 8176 11004
rect 8120 10950 8122 11002
rect 8122 10950 8174 11002
rect 8174 10950 8176 11002
rect 8120 10948 8176 10950
rect 8224 11002 8280 11004
rect 8224 10950 8226 11002
rect 8226 10950 8278 11002
rect 8278 10950 8280 11002
rect 8224 10948 8280 10950
rect 8092 10834 8148 10836
rect 8092 10782 8094 10834
rect 8094 10782 8146 10834
rect 8146 10782 8148 10834
rect 8092 10780 8148 10782
rect 4844 9324 4900 9380
rect 4614 8650 4670 8652
rect 4614 8598 4616 8650
rect 4616 8598 4668 8650
rect 4668 8598 4670 8650
rect 4614 8596 4670 8598
rect 4718 8650 4774 8652
rect 4718 8598 4720 8650
rect 4720 8598 4772 8650
rect 4772 8598 4774 8650
rect 4718 8596 4774 8598
rect 4822 8650 4878 8652
rect 4822 8598 4824 8650
rect 4824 8598 4876 8650
rect 4876 8598 4878 8650
rect 4822 8596 4878 8598
rect 4844 8316 4900 8372
rect 9100 12012 9156 12068
rect 8540 11340 8596 11396
rect 8988 10444 9044 10500
rect 11418 14922 11474 14924
rect 11418 14870 11420 14922
rect 11420 14870 11472 14922
rect 11472 14870 11474 14922
rect 11418 14868 11474 14870
rect 11522 14922 11578 14924
rect 11522 14870 11524 14922
rect 11524 14870 11576 14922
rect 11576 14870 11578 14922
rect 11522 14868 11578 14870
rect 11626 14922 11682 14924
rect 11626 14870 11628 14922
rect 11628 14870 11680 14922
rect 11680 14870 11682 14922
rect 11626 14868 11682 14870
rect 11228 13468 11284 13524
rect 11418 13354 11474 13356
rect 11418 13302 11420 13354
rect 11420 13302 11472 13354
rect 11472 13302 11474 13354
rect 11418 13300 11474 13302
rect 11522 13354 11578 13356
rect 11522 13302 11524 13354
rect 11524 13302 11576 13354
rect 11576 13302 11578 13354
rect 11522 13300 11578 13302
rect 11626 13354 11682 13356
rect 11626 13302 11628 13354
rect 11628 13302 11680 13354
rect 11680 13302 11682 13354
rect 11788 13356 11844 13412
rect 11626 13300 11682 13302
rect 12460 13132 12516 13188
rect 10780 12066 10836 12068
rect 10780 12014 10782 12066
rect 10782 12014 10834 12066
rect 10834 12014 10836 12066
rect 10780 12012 10836 12014
rect 9884 10498 9940 10500
rect 9884 10446 9886 10498
rect 9886 10446 9938 10498
rect 9938 10446 9940 10498
rect 9884 10444 9940 10446
rect 8016 9434 8072 9436
rect 6636 9324 6692 9380
rect 8016 9382 8018 9434
rect 8018 9382 8070 9434
rect 8070 9382 8072 9434
rect 8016 9380 8072 9382
rect 8120 9434 8176 9436
rect 8120 9382 8122 9434
rect 8122 9382 8174 9434
rect 8174 9382 8176 9434
rect 8120 9380 8176 9382
rect 8224 9434 8280 9436
rect 8224 9382 8226 9434
rect 8226 9382 8278 9434
rect 8278 9382 8280 9434
rect 8224 9380 8280 9382
rect 5852 8370 5908 8372
rect 5852 8318 5854 8370
rect 5854 8318 5906 8370
rect 5906 8318 5908 8370
rect 5852 8316 5908 8318
rect 6412 8092 6468 8148
rect 7756 8146 7812 8148
rect 7756 8094 7758 8146
rect 7758 8094 7810 8146
rect 7810 8094 7812 8146
rect 7756 8092 7812 8094
rect 8016 7866 8072 7868
rect 8016 7814 8018 7866
rect 8018 7814 8070 7866
rect 8070 7814 8072 7866
rect 8016 7812 8072 7814
rect 8120 7866 8176 7868
rect 8120 7814 8122 7866
rect 8122 7814 8174 7866
rect 8174 7814 8176 7866
rect 8120 7812 8176 7814
rect 8224 7866 8280 7868
rect 8224 7814 8226 7866
rect 8226 7814 8278 7866
rect 8278 7814 8280 7866
rect 8224 7812 8280 7814
rect 4614 7082 4670 7084
rect 4614 7030 4616 7082
rect 4616 7030 4668 7082
rect 4668 7030 4670 7082
rect 4614 7028 4670 7030
rect 4718 7082 4774 7084
rect 4718 7030 4720 7082
rect 4720 7030 4772 7082
rect 4772 7030 4774 7082
rect 4718 7028 4774 7030
rect 4822 7082 4878 7084
rect 4822 7030 4824 7082
rect 4824 7030 4876 7082
rect 4876 7030 4878 7082
rect 4822 7028 4878 7030
rect 8016 6298 8072 6300
rect 8016 6246 8018 6298
rect 8018 6246 8070 6298
rect 8070 6246 8072 6298
rect 8016 6244 8072 6246
rect 8120 6298 8176 6300
rect 8120 6246 8122 6298
rect 8122 6246 8174 6298
rect 8174 6246 8176 6298
rect 8120 6244 8176 6246
rect 8224 6298 8280 6300
rect 8224 6246 8226 6298
rect 8226 6246 8278 6298
rect 8278 6246 8280 6298
rect 8224 6244 8280 6246
rect 1708 6076 1764 6132
rect 4614 5514 4670 5516
rect 4614 5462 4616 5514
rect 4616 5462 4668 5514
rect 4668 5462 4670 5514
rect 4614 5460 4670 5462
rect 4718 5514 4774 5516
rect 4718 5462 4720 5514
rect 4720 5462 4772 5514
rect 4772 5462 4774 5514
rect 4718 5460 4774 5462
rect 4822 5514 4878 5516
rect 4822 5462 4824 5514
rect 4824 5462 4876 5514
rect 4876 5462 4878 5514
rect 4822 5460 4878 5462
rect 11418 11786 11474 11788
rect 11418 11734 11420 11786
rect 11420 11734 11472 11786
rect 11472 11734 11474 11786
rect 11418 11732 11474 11734
rect 11522 11786 11578 11788
rect 11522 11734 11524 11786
rect 11524 11734 11576 11786
rect 11576 11734 11578 11786
rect 11522 11732 11578 11734
rect 11626 11786 11682 11788
rect 11626 11734 11628 11786
rect 11628 11734 11680 11786
rect 11680 11734 11682 11786
rect 11626 11732 11682 11734
rect 11228 11170 11284 11172
rect 11228 11118 11230 11170
rect 11230 11118 11282 11170
rect 11282 11118 11284 11170
rect 11228 11116 11284 11118
rect 14476 14642 14532 14644
rect 14476 14590 14478 14642
rect 14478 14590 14530 14642
rect 14530 14590 14532 14642
rect 14476 14588 14532 14590
rect 13020 14418 13076 14420
rect 13020 14366 13022 14418
rect 13022 14366 13074 14418
rect 13074 14366 13076 14418
rect 13020 14364 13076 14366
rect 13916 13356 13972 13412
rect 13468 13186 13524 13188
rect 13468 13134 13470 13186
rect 13470 13134 13522 13186
rect 13522 13134 13524 13186
rect 13468 13132 13524 13134
rect 14820 17274 14876 17276
rect 14820 17222 14822 17274
rect 14822 17222 14874 17274
rect 14874 17222 14876 17274
rect 14820 17220 14876 17222
rect 14924 17274 14980 17276
rect 14924 17222 14926 17274
rect 14926 17222 14978 17274
rect 14978 17222 14980 17274
rect 14924 17220 14980 17222
rect 15028 17274 15084 17276
rect 15028 17222 15030 17274
rect 15030 17222 15082 17274
rect 15082 17222 15084 17274
rect 15028 17220 15084 17222
rect 16044 16828 16100 16884
rect 14820 15706 14876 15708
rect 14820 15654 14822 15706
rect 14822 15654 14874 15706
rect 14874 15654 14876 15706
rect 14820 15652 14876 15654
rect 14924 15706 14980 15708
rect 14924 15654 14926 15706
rect 14926 15654 14978 15706
rect 14978 15654 14980 15706
rect 14924 15652 14980 15654
rect 15028 15706 15084 15708
rect 15028 15654 15030 15706
rect 15030 15654 15082 15706
rect 15082 15654 15084 15706
rect 15028 15652 15084 15654
rect 15036 15314 15092 15316
rect 15036 15262 15038 15314
rect 15038 15262 15090 15314
rect 15090 15262 15092 15314
rect 15036 15260 15092 15262
rect 21084 20018 21140 20020
rect 21084 19966 21086 20018
rect 21086 19966 21138 20018
rect 21138 19966 21140 20018
rect 21084 19964 21140 19966
rect 20748 19852 20804 19908
rect 18222 19626 18278 19628
rect 18222 19574 18224 19626
rect 18224 19574 18276 19626
rect 18276 19574 18278 19626
rect 18222 19572 18278 19574
rect 18326 19626 18382 19628
rect 18326 19574 18328 19626
rect 18328 19574 18380 19626
rect 18380 19574 18382 19626
rect 18326 19572 18382 19574
rect 18430 19626 18486 19628
rect 18430 19574 18432 19626
rect 18432 19574 18484 19626
rect 18484 19574 18486 19626
rect 18430 19572 18486 19574
rect 18060 19292 18116 19348
rect 19180 19346 19236 19348
rect 19180 19294 19182 19346
rect 19182 19294 19234 19346
rect 19234 19294 19236 19346
rect 19180 19292 19236 19294
rect 17948 19122 18004 19124
rect 17948 19070 17950 19122
rect 17950 19070 18002 19122
rect 18002 19070 18004 19122
rect 17948 19068 18004 19070
rect 20188 19122 20244 19124
rect 20188 19070 20190 19122
rect 20190 19070 20242 19122
rect 20242 19070 20244 19122
rect 20188 19068 20244 19070
rect 19404 18562 19460 18564
rect 19404 18510 19406 18562
rect 19406 18510 19458 18562
rect 19458 18510 19460 18562
rect 19404 18508 19460 18510
rect 18396 18172 18452 18228
rect 18222 18058 18278 18060
rect 18222 18006 18224 18058
rect 18224 18006 18276 18058
rect 18276 18006 18278 18058
rect 18222 18004 18278 18006
rect 18326 18058 18382 18060
rect 18326 18006 18328 18058
rect 18328 18006 18380 18058
rect 18380 18006 18382 18058
rect 18326 18004 18382 18006
rect 18430 18058 18486 18060
rect 18430 18006 18432 18058
rect 18432 18006 18484 18058
rect 18484 18006 18486 18058
rect 18430 18004 18486 18006
rect 19292 17442 19348 17444
rect 19292 17390 19294 17442
rect 19294 17390 19346 17442
rect 19346 17390 19348 17442
rect 19292 17388 19348 17390
rect 17612 16828 17668 16884
rect 17948 16882 18004 16884
rect 17948 16830 17950 16882
rect 17950 16830 18002 16882
rect 18002 16830 18004 16882
rect 17948 16828 18004 16830
rect 18222 16490 18278 16492
rect 18222 16438 18224 16490
rect 18224 16438 18276 16490
rect 18276 16438 18278 16490
rect 18222 16436 18278 16438
rect 18326 16490 18382 16492
rect 18326 16438 18328 16490
rect 18328 16438 18380 16490
rect 18380 16438 18382 16490
rect 18326 16436 18382 16438
rect 18430 16490 18486 16492
rect 18430 16438 18432 16490
rect 18432 16438 18484 16490
rect 18484 16438 18486 16490
rect 18430 16436 18486 16438
rect 20076 17442 20132 17444
rect 20076 17390 20078 17442
rect 20078 17390 20130 17442
rect 20130 17390 20132 17442
rect 20076 17388 20132 17390
rect 19852 15932 19908 15988
rect 22316 19906 22372 19908
rect 22316 19854 22318 19906
rect 22318 19854 22370 19906
rect 22370 19854 22372 19906
rect 22316 19852 22372 19854
rect 21624 18842 21680 18844
rect 21624 18790 21626 18842
rect 21626 18790 21678 18842
rect 21678 18790 21680 18842
rect 21624 18788 21680 18790
rect 21728 18842 21784 18844
rect 21728 18790 21730 18842
rect 21730 18790 21782 18842
rect 21782 18790 21784 18842
rect 21728 18788 21784 18790
rect 21832 18842 21888 18844
rect 21832 18790 21834 18842
rect 21834 18790 21886 18842
rect 21886 18790 21888 18842
rect 21832 18788 21888 18790
rect 21420 18284 21476 18340
rect 20076 16828 20132 16884
rect 20636 17666 20692 17668
rect 20636 17614 20638 17666
rect 20638 17614 20690 17666
rect 20690 17614 20692 17666
rect 20636 17612 20692 17614
rect 20300 15986 20356 15988
rect 20300 15934 20302 15986
rect 20302 15934 20354 15986
rect 20354 15934 20356 15986
rect 20300 15932 20356 15934
rect 20524 15314 20580 15316
rect 20524 15262 20526 15314
rect 20526 15262 20578 15314
rect 20578 15262 20580 15314
rect 20524 15260 20580 15262
rect 18222 14922 18278 14924
rect 18222 14870 18224 14922
rect 18224 14870 18276 14922
rect 18276 14870 18278 14922
rect 18222 14868 18278 14870
rect 18326 14922 18382 14924
rect 18326 14870 18328 14922
rect 18328 14870 18380 14922
rect 18380 14870 18382 14922
rect 18326 14868 18382 14870
rect 18430 14922 18486 14924
rect 18430 14870 18432 14922
rect 18432 14870 18484 14922
rect 18484 14870 18486 14922
rect 18430 14868 18486 14870
rect 21420 17612 21476 17668
rect 21624 17274 21680 17276
rect 21624 17222 21626 17274
rect 21626 17222 21678 17274
rect 21678 17222 21680 17274
rect 21624 17220 21680 17222
rect 21728 17274 21784 17276
rect 21728 17222 21730 17274
rect 21730 17222 21782 17274
rect 21782 17222 21784 17274
rect 21728 17220 21784 17222
rect 21832 17274 21888 17276
rect 21832 17222 21834 17274
rect 21834 17222 21886 17274
rect 21886 17222 21888 17274
rect 21832 17220 21888 17222
rect 21644 17106 21700 17108
rect 21644 17054 21646 17106
rect 21646 17054 21698 17106
rect 21698 17054 21700 17106
rect 21644 17052 21700 17054
rect 24444 20914 24500 20916
rect 24444 20862 24446 20914
rect 24446 20862 24498 20914
rect 24498 20862 24500 20914
rect 24444 20860 24500 20862
rect 23548 19964 23604 20020
rect 23772 19964 23828 20020
rect 23212 19740 23268 19796
rect 26124 26514 26180 26516
rect 26124 26462 26126 26514
rect 26126 26462 26178 26514
rect 26178 26462 26180 26514
rect 26124 26460 26180 26462
rect 26124 26236 26180 26292
rect 25452 24946 25508 24948
rect 25452 24894 25454 24946
rect 25454 24894 25506 24946
rect 25506 24894 25508 24946
rect 25452 24892 25508 24894
rect 25564 25228 25620 25284
rect 24668 23772 24724 23828
rect 25026 24330 25082 24332
rect 25026 24278 25028 24330
rect 25028 24278 25080 24330
rect 25080 24278 25082 24330
rect 25026 24276 25082 24278
rect 25130 24330 25186 24332
rect 25130 24278 25132 24330
rect 25132 24278 25184 24330
rect 25184 24278 25186 24330
rect 25130 24276 25186 24278
rect 25234 24330 25290 24332
rect 25234 24278 25236 24330
rect 25236 24278 25288 24330
rect 25288 24278 25290 24330
rect 25234 24276 25290 24278
rect 25228 23938 25284 23940
rect 25228 23886 25230 23938
rect 25230 23886 25282 23938
rect 25282 23886 25284 23938
rect 25228 23884 25284 23886
rect 25900 24780 25956 24836
rect 26908 25282 26964 25284
rect 26908 25230 26910 25282
rect 26910 25230 26962 25282
rect 26962 25230 26964 25282
rect 26908 25228 26964 25230
rect 25788 23660 25844 23716
rect 24668 23266 24724 23268
rect 24668 23214 24670 23266
rect 24670 23214 24722 23266
rect 24722 23214 24724 23266
rect 24668 23212 24724 23214
rect 25026 22762 25082 22764
rect 25026 22710 25028 22762
rect 25028 22710 25080 22762
rect 25080 22710 25082 22762
rect 25026 22708 25082 22710
rect 25130 22762 25186 22764
rect 25130 22710 25132 22762
rect 25132 22710 25184 22762
rect 25184 22710 25186 22762
rect 25130 22708 25186 22710
rect 25234 22762 25290 22764
rect 25234 22710 25236 22762
rect 25236 22710 25288 22762
rect 25288 22710 25290 22762
rect 25234 22708 25290 22710
rect 26236 22764 26292 22820
rect 25026 21194 25082 21196
rect 25026 21142 25028 21194
rect 25028 21142 25080 21194
rect 25080 21142 25082 21194
rect 25026 21140 25082 21142
rect 25130 21194 25186 21196
rect 25130 21142 25132 21194
rect 25132 21142 25184 21194
rect 25184 21142 25186 21194
rect 25130 21140 25186 21142
rect 25234 21194 25290 21196
rect 25234 21142 25236 21194
rect 25236 21142 25288 21194
rect 25288 21142 25290 21194
rect 25234 21140 25290 21142
rect 24556 20076 24612 20132
rect 23996 19852 24052 19908
rect 24108 19794 24164 19796
rect 24108 19742 24110 19794
rect 24110 19742 24162 19794
rect 24162 19742 24164 19794
rect 24108 19740 24164 19742
rect 23884 18956 23940 19012
rect 23100 18284 23156 18340
rect 21980 16882 22036 16884
rect 21980 16830 21982 16882
rect 21982 16830 22034 16882
rect 22034 16830 22036 16882
rect 21980 16828 22036 16830
rect 21624 15706 21680 15708
rect 21624 15654 21626 15706
rect 21626 15654 21678 15706
rect 21678 15654 21680 15706
rect 21624 15652 21680 15654
rect 21728 15706 21784 15708
rect 21728 15654 21730 15706
rect 21730 15654 21782 15706
rect 21782 15654 21784 15706
rect 21728 15652 21784 15654
rect 21832 15706 21888 15708
rect 21832 15654 21834 15706
rect 21834 15654 21886 15706
rect 21886 15654 21888 15706
rect 21832 15652 21888 15654
rect 15484 14418 15540 14420
rect 15484 14366 15486 14418
rect 15486 14366 15538 14418
rect 15538 14366 15540 14418
rect 15484 14364 15540 14366
rect 18060 14252 18116 14308
rect 14820 14138 14876 14140
rect 14820 14086 14822 14138
rect 14822 14086 14874 14138
rect 14874 14086 14876 14138
rect 14820 14084 14876 14086
rect 14924 14138 14980 14140
rect 14924 14086 14926 14138
rect 14926 14086 14978 14138
rect 14978 14086 14980 14138
rect 14924 14084 14980 14086
rect 15028 14138 15084 14140
rect 15028 14086 15030 14138
rect 15030 14086 15082 14138
rect 15082 14086 15084 14138
rect 15028 14084 15084 14086
rect 14588 13020 14644 13076
rect 16828 13074 16884 13076
rect 16828 13022 16830 13074
rect 16830 13022 16882 13074
rect 16882 13022 16884 13074
rect 16828 13020 16884 13022
rect 15148 12962 15204 12964
rect 15148 12910 15150 12962
rect 15150 12910 15202 12962
rect 15202 12910 15204 12962
rect 15148 12908 15204 12910
rect 14820 12570 14876 12572
rect 14820 12518 14822 12570
rect 14822 12518 14874 12570
rect 14874 12518 14876 12570
rect 14820 12516 14876 12518
rect 14924 12570 14980 12572
rect 14924 12518 14926 12570
rect 14926 12518 14978 12570
rect 14978 12518 14980 12570
rect 14924 12516 14980 12518
rect 15028 12570 15084 12572
rect 15028 12518 15030 12570
rect 15030 12518 15082 12570
rect 15082 12518 15084 12570
rect 15028 12516 15084 12518
rect 19852 14306 19908 14308
rect 19852 14254 19854 14306
rect 19854 14254 19906 14306
rect 19906 14254 19908 14306
rect 19852 14252 19908 14254
rect 21624 14138 21680 14140
rect 21624 14086 21626 14138
rect 21626 14086 21678 14138
rect 21678 14086 21680 14138
rect 21624 14084 21680 14086
rect 21728 14138 21784 14140
rect 21728 14086 21730 14138
rect 21730 14086 21782 14138
rect 21782 14086 21784 14138
rect 21728 14084 21784 14086
rect 21832 14138 21888 14140
rect 21832 14086 21834 14138
rect 21834 14086 21886 14138
rect 21886 14086 21888 14138
rect 21832 14084 21888 14086
rect 18222 13354 18278 13356
rect 18222 13302 18224 13354
rect 18224 13302 18276 13354
rect 18276 13302 18278 13354
rect 18222 13300 18278 13302
rect 18326 13354 18382 13356
rect 18326 13302 18328 13354
rect 18328 13302 18380 13354
rect 18380 13302 18382 13354
rect 18326 13300 18382 13302
rect 18430 13354 18486 13356
rect 18430 13302 18432 13354
rect 18432 13302 18484 13354
rect 18484 13302 18486 13354
rect 18430 13300 18486 13302
rect 18222 11786 18278 11788
rect 18222 11734 18224 11786
rect 18224 11734 18276 11786
rect 18276 11734 18278 11786
rect 18222 11732 18278 11734
rect 18326 11786 18382 11788
rect 18326 11734 18328 11786
rect 18328 11734 18380 11786
rect 18380 11734 18382 11786
rect 18326 11732 18382 11734
rect 18430 11786 18486 11788
rect 18430 11734 18432 11786
rect 18432 11734 18484 11786
rect 18484 11734 18486 11786
rect 18430 11732 18486 11734
rect 19628 11788 19684 11844
rect 12236 10444 12292 10500
rect 12684 10556 12740 10612
rect 11418 10218 11474 10220
rect 11418 10166 11420 10218
rect 11420 10166 11472 10218
rect 11472 10166 11474 10218
rect 11418 10164 11474 10166
rect 11522 10218 11578 10220
rect 11522 10166 11524 10218
rect 11524 10166 11576 10218
rect 11576 10166 11578 10218
rect 11522 10164 11578 10166
rect 11626 10218 11682 10220
rect 11626 10166 11628 10218
rect 11628 10166 11680 10218
rect 11680 10166 11682 10218
rect 11626 10164 11682 10166
rect 13468 10610 13524 10612
rect 13468 10558 13470 10610
rect 13470 10558 13522 10610
rect 13522 10558 13524 10610
rect 13468 10556 13524 10558
rect 10780 8988 10836 9044
rect 12236 9042 12292 9044
rect 12236 8990 12238 9042
rect 12238 8990 12290 9042
rect 12290 8990 12292 9042
rect 12236 8988 12292 8990
rect 11418 8650 11474 8652
rect 11418 8598 11420 8650
rect 11420 8598 11472 8650
rect 11472 8598 11474 8650
rect 11418 8596 11474 8598
rect 11522 8650 11578 8652
rect 11522 8598 11524 8650
rect 11524 8598 11576 8650
rect 11576 8598 11578 8650
rect 11522 8596 11578 8598
rect 11626 8650 11682 8652
rect 11626 8598 11628 8650
rect 11628 8598 11680 8650
rect 11680 8598 11682 8650
rect 11626 8596 11682 8598
rect 12908 7868 12964 7924
rect 15820 11116 15876 11172
rect 14820 11002 14876 11004
rect 14820 10950 14822 11002
rect 14822 10950 14874 11002
rect 14874 10950 14876 11002
rect 14820 10948 14876 10950
rect 14924 11002 14980 11004
rect 14924 10950 14926 11002
rect 14926 10950 14978 11002
rect 14978 10950 14980 11002
rect 14924 10948 14980 10950
rect 15028 11002 15084 11004
rect 15028 10950 15030 11002
rect 15030 10950 15082 11002
rect 15082 10950 15084 11002
rect 15028 10948 15084 10950
rect 14140 10556 14196 10612
rect 17500 10556 17556 10612
rect 14812 10498 14868 10500
rect 14812 10446 14814 10498
rect 14814 10446 14866 10498
rect 14866 10446 14868 10498
rect 14812 10444 14868 10446
rect 18284 10610 18340 10612
rect 18284 10558 18286 10610
rect 18286 10558 18338 10610
rect 18338 10558 18340 10610
rect 18284 10556 18340 10558
rect 21756 13746 21812 13748
rect 21756 13694 21758 13746
rect 21758 13694 21810 13746
rect 21810 13694 21812 13746
rect 21756 13692 21812 13694
rect 25340 19964 25396 20020
rect 25026 19626 25082 19628
rect 25026 19574 25028 19626
rect 25028 19574 25080 19626
rect 25080 19574 25082 19626
rect 25026 19572 25082 19574
rect 25130 19626 25186 19628
rect 25130 19574 25132 19626
rect 25132 19574 25184 19626
rect 25184 19574 25186 19626
rect 25130 19572 25186 19574
rect 25234 19626 25290 19628
rect 25234 19574 25236 19626
rect 25236 19574 25288 19626
rect 25288 19574 25290 19626
rect 25234 19572 25290 19574
rect 24444 18284 24500 18340
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 25026 18058 25082 18060
rect 25026 18006 25028 18058
rect 25028 18006 25080 18058
rect 25080 18006 25082 18058
rect 25026 18004 25082 18006
rect 25130 18058 25186 18060
rect 25130 18006 25132 18058
rect 25132 18006 25184 18058
rect 25184 18006 25186 18058
rect 25130 18004 25186 18006
rect 25234 18058 25290 18060
rect 25234 18006 25236 18058
rect 25236 18006 25288 18058
rect 25288 18006 25290 18058
rect 25234 18004 25290 18006
rect 23324 16940 23380 16996
rect 23996 16994 24052 16996
rect 23996 16942 23998 16994
rect 23998 16942 24050 16994
rect 24050 16942 24052 16994
rect 23996 16940 24052 16942
rect 25026 16490 25082 16492
rect 25026 16438 25028 16490
rect 25028 16438 25080 16490
rect 25080 16438 25082 16490
rect 25026 16436 25082 16438
rect 25130 16490 25186 16492
rect 25130 16438 25132 16490
rect 25132 16438 25184 16490
rect 25184 16438 25186 16490
rect 25130 16436 25186 16438
rect 25234 16490 25290 16492
rect 25234 16438 25236 16490
rect 25236 16438 25288 16490
rect 25288 16438 25290 16490
rect 25234 16436 25290 16438
rect 22876 15484 22932 15540
rect 24556 15372 24612 15428
rect 25340 15372 25396 15428
rect 22428 15148 22484 15204
rect 23212 15148 23268 15204
rect 22540 13580 22596 13636
rect 21980 13020 22036 13076
rect 21624 12570 21680 12572
rect 21624 12518 21626 12570
rect 21626 12518 21678 12570
rect 21678 12518 21680 12570
rect 21624 12516 21680 12518
rect 21728 12570 21784 12572
rect 21728 12518 21730 12570
rect 21730 12518 21782 12570
rect 21782 12518 21784 12570
rect 21728 12516 21784 12518
rect 21832 12570 21888 12572
rect 21832 12518 21834 12570
rect 21834 12518 21886 12570
rect 21886 12518 21888 12570
rect 21832 12516 21888 12518
rect 21308 11788 21364 11844
rect 20524 11452 20580 11508
rect 25788 21196 25844 21252
rect 26236 21756 26292 21812
rect 26908 24108 26964 24164
rect 26908 23714 26964 23716
rect 26908 23662 26910 23714
rect 26910 23662 26962 23714
rect 26962 23662 26964 23714
rect 26908 23660 26964 23662
rect 26908 23266 26964 23268
rect 26908 23214 26910 23266
rect 26910 23214 26962 23266
rect 26962 23214 26964 23266
rect 26908 23212 26964 23214
rect 27692 25564 27748 25620
rect 27692 24892 27748 24948
rect 28428 26682 28484 26684
rect 28428 26630 28430 26682
rect 28430 26630 28482 26682
rect 28482 26630 28484 26682
rect 28428 26628 28484 26630
rect 28532 26682 28588 26684
rect 28532 26630 28534 26682
rect 28534 26630 28586 26682
rect 28586 26630 28588 26682
rect 28532 26628 28588 26630
rect 28636 26682 28692 26684
rect 28636 26630 28638 26682
rect 28638 26630 28690 26682
rect 28690 26630 28692 26682
rect 28636 26628 28692 26630
rect 28428 25114 28484 25116
rect 28428 25062 28430 25114
rect 28430 25062 28482 25114
rect 28482 25062 28484 25114
rect 28428 25060 28484 25062
rect 28532 25114 28588 25116
rect 28532 25062 28534 25114
rect 28534 25062 28586 25114
rect 28586 25062 28588 25114
rect 28532 25060 28588 25062
rect 28636 25114 28692 25116
rect 28636 25062 28638 25114
rect 28638 25062 28690 25114
rect 28690 25062 28692 25114
rect 28636 25060 28692 25062
rect 28028 24220 28084 24276
rect 28428 23546 28484 23548
rect 28428 23494 28430 23546
rect 28430 23494 28482 23546
rect 28482 23494 28484 23546
rect 28428 23492 28484 23494
rect 28532 23546 28588 23548
rect 28532 23494 28534 23546
rect 28534 23494 28586 23546
rect 28586 23494 28588 23546
rect 28532 23492 28588 23494
rect 28636 23546 28692 23548
rect 28636 23494 28638 23546
rect 28638 23494 28690 23546
rect 28690 23494 28692 23546
rect 28636 23492 28692 23494
rect 26796 22876 26852 22932
rect 26908 22764 26964 22820
rect 28028 22258 28084 22260
rect 28028 22206 28030 22258
rect 28030 22206 28082 22258
rect 28082 22206 28084 22258
rect 28028 22204 28084 22206
rect 27804 21810 27860 21812
rect 27804 21758 27806 21810
rect 27806 21758 27858 21810
rect 27858 21758 27860 21810
rect 27804 21756 27860 21758
rect 26684 21532 26740 21588
rect 26236 21474 26292 21476
rect 26236 21422 26238 21474
rect 26238 21422 26290 21474
rect 26290 21422 26292 21474
rect 26236 21420 26292 21422
rect 27132 21698 27188 21700
rect 27132 21646 27134 21698
rect 27134 21646 27186 21698
rect 27186 21646 27188 21698
rect 27132 21644 27188 21646
rect 27468 21586 27524 21588
rect 27468 21534 27470 21586
rect 27470 21534 27522 21586
rect 27522 21534 27524 21586
rect 27468 21532 27524 21534
rect 28428 21978 28484 21980
rect 28428 21926 28430 21978
rect 28430 21926 28482 21978
rect 28482 21926 28484 21978
rect 28428 21924 28484 21926
rect 28532 21978 28588 21980
rect 28532 21926 28534 21978
rect 28534 21926 28586 21978
rect 28586 21926 28588 21978
rect 28532 21924 28588 21926
rect 28636 21978 28692 21980
rect 28636 21926 28638 21978
rect 28638 21926 28690 21978
rect 28690 21926 28692 21978
rect 28636 21924 28692 21926
rect 26796 21420 26852 21476
rect 27468 21196 27524 21252
rect 25900 20748 25956 20804
rect 26908 20802 26964 20804
rect 26908 20750 26910 20802
rect 26910 20750 26962 20802
rect 26962 20750 26964 20802
rect 26908 20748 26964 20750
rect 26236 19906 26292 19908
rect 26236 19854 26238 19906
rect 26238 19854 26290 19906
rect 26290 19854 26292 19906
rect 26236 19852 26292 19854
rect 26124 19010 26180 19012
rect 26124 18958 26126 19010
rect 26126 18958 26178 19010
rect 26178 18958 26180 19010
rect 26124 18956 26180 18958
rect 28140 20860 28196 20916
rect 28428 20410 28484 20412
rect 28428 20358 28430 20410
rect 28430 20358 28482 20410
rect 28482 20358 28484 20410
rect 28428 20356 28484 20358
rect 28532 20410 28588 20412
rect 28532 20358 28534 20410
rect 28534 20358 28586 20410
rect 28586 20358 28588 20410
rect 28532 20356 28588 20358
rect 28636 20410 28692 20412
rect 28636 20358 28638 20410
rect 28638 20358 28690 20410
rect 28690 20358 28692 20410
rect 28636 20356 28692 20358
rect 28028 20188 28084 20244
rect 27804 20130 27860 20132
rect 27804 20078 27806 20130
rect 27806 20078 27858 20130
rect 27858 20078 27860 20130
rect 27804 20076 27860 20078
rect 28140 19516 28196 19572
rect 27580 19010 27636 19012
rect 27580 18958 27582 19010
rect 27582 18958 27634 19010
rect 27634 18958 27636 19010
rect 27580 18956 27636 18958
rect 28140 18956 28196 19012
rect 28428 18842 28484 18844
rect 28428 18790 28430 18842
rect 28430 18790 28482 18842
rect 28482 18790 28484 18842
rect 28428 18788 28484 18790
rect 28532 18842 28588 18844
rect 28532 18790 28534 18842
rect 28534 18790 28586 18842
rect 28586 18790 28588 18842
rect 28532 18788 28588 18790
rect 28636 18842 28692 18844
rect 28636 18790 28638 18842
rect 28638 18790 28690 18842
rect 28690 18790 28692 18842
rect 28636 18788 28692 18790
rect 26348 18284 26404 18340
rect 26348 17666 26404 17668
rect 26348 17614 26350 17666
rect 26350 17614 26402 17666
rect 26402 17614 26404 17666
rect 26348 17612 26404 17614
rect 25564 17500 25620 17556
rect 27692 18172 27748 18228
rect 28140 18172 28196 18228
rect 27132 17612 27188 17668
rect 27804 17554 27860 17556
rect 27804 17502 27806 17554
rect 27806 17502 27858 17554
rect 27858 17502 27860 17554
rect 27804 17500 27860 17502
rect 27244 17052 27300 17108
rect 23548 15090 23604 15092
rect 23548 15038 23550 15090
rect 23550 15038 23602 15090
rect 23602 15038 23604 15090
rect 23548 15036 23604 15038
rect 23660 14700 23716 14756
rect 25026 14922 25082 14924
rect 25026 14870 25028 14922
rect 25028 14870 25080 14922
rect 25080 14870 25082 14922
rect 25026 14868 25082 14870
rect 25130 14922 25186 14924
rect 25130 14870 25132 14922
rect 25132 14870 25184 14922
rect 25184 14870 25186 14922
rect 25130 14868 25186 14870
rect 25234 14922 25290 14924
rect 25234 14870 25236 14922
rect 25236 14870 25288 14922
rect 25288 14870 25290 14922
rect 25234 14868 25290 14870
rect 25564 15596 25620 15652
rect 25788 15202 25844 15204
rect 25788 15150 25790 15202
rect 25790 15150 25842 15202
rect 25842 15150 25844 15202
rect 25788 15148 25844 15150
rect 26236 15260 26292 15316
rect 28428 17274 28484 17276
rect 28428 17222 28430 17274
rect 28430 17222 28482 17274
rect 28482 17222 28484 17274
rect 28428 17220 28484 17222
rect 28532 17274 28588 17276
rect 28532 17222 28534 17274
rect 28534 17222 28586 17274
rect 28586 17222 28588 17274
rect 28532 17220 28588 17222
rect 28636 17274 28692 17276
rect 28636 17222 28638 17274
rect 28638 17222 28690 17274
rect 28690 17222 28692 17274
rect 28636 17220 28692 17222
rect 27692 15596 27748 15652
rect 28428 15706 28484 15708
rect 28428 15654 28430 15706
rect 28430 15654 28482 15706
rect 28482 15654 28484 15706
rect 28428 15652 28484 15654
rect 28532 15706 28588 15708
rect 28532 15654 28534 15706
rect 28534 15654 28586 15706
rect 28586 15654 28588 15706
rect 28532 15652 28588 15654
rect 28636 15706 28692 15708
rect 28636 15654 28638 15706
rect 28638 15654 28690 15706
rect 28690 15654 28692 15706
rect 28636 15652 28692 15654
rect 27356 15148 27412 15204
rect 27692 15148 27748 15204
rect 26684 14700 26740 14756
rect 27244 15036 27300 15092
rect 25452 14476 25508 14532
rect 24220 14252 24276 14308
rect 24780 13522 24836 13524
rect 24780 13470 24782 13522
rect 24782 13470 24834 13522
rect 24834 13470 24836 13522
rect 24780 13468 24836 13470
rect 25026 13354 25082 13356
rect 25026 13302 25028 13354
rect 25028 13302 25080 13354
rect 25080 13302 25082 13354
rect 25026 13300 25082 13302
rect 25130 13354 25186 13356
rect 25130 13302 25132 13354
rect 25132 13302 25184 13354
rect 25184 13302 25186 13354
rect 25130 13300 25186 13302
rect 25234 13354 25290 13356
rect 25234 13302 25236 13354
rect 25236 13302 25288 13354
rect 25288 13302 25290 13354
rect 25234 13300 25290 13302
rect 26348 14530 26404 14532
rect 26348 14478 26350 14530
rect 26350 14478 26402 14530
rect 26402 14478 26404 14530
rect 26348 14476 26404 14478
rect 27132 14530 27188 14532
rect 27132 14478 27134 14530
rect 27134 14478 27186 14530
rect 27186 14478 27188 14530
rect 27132 14476 27188 14478
rect 26684 14306 26740 14308
rect 26684 14254 26686 14306
rect 26686 14254 26738 14306
rect 26738 14254 26740 14306
rect 26684 14252 26740 14254
rect 28140 14530 28196 14532
rect 28140 14478 28142 14530
rect 28142 14478 28194 14530
rect 28194 14478 28196 14530
rect 28140 14476 28196 14478
rect 26460 13692 26516 13748
rect 22876 11900 22932 11956
rect 23436 11676 23492 11732
rect 23660 11452 23716 11508
rect 23436 11228 23492 11284
rect 20748 11170 20804 11172
rect 20748 11118 20750 11170
rect 20750 11118 20802 11170
rect 20802 11118 20804 11170
rect 20748 11116 20804 11118
rect 22316 11116 22372 11172
rect 21624 11002 21680 11004
rect 21624 10950 21626 11002
rect 21626 10950 21678 11002
rect 21678 10950 21680 11002
rect 21624 10948 21680 10950
rect 21728 11002 21784 11004
rect 21728 10950 21730 11002
rect 21730 10950 21782 11002
rect 21782 10950 21784 11002
rect 21728 10948 21784 10950
rect 21832 11002 21888 11004
rect 21832 10950 21834 11002
rect 21834 10950 21886 11002
rect 21886 10950 21888 11002
rect 21832 10948 21888 10950
rect 23100 10722 23156 10724
rect 23100 10670 23102 10722
rect 23102 10670 23154 10722
rect 23154 10670 23156 10722
rect 23100 10668 23156 10670
rect 20300 10556 20356 10612
rect 23884 10610 23940 10612
rect 23884 10558 23886 10610
rect 23886 10558 23938 10610
rect 23938 10558 23940 10610
rect 23884 10556 23940 10558
rect 21980 10444 22036 10500
rect 14820 9434 14876 9436
rect 14820 9382 14822 9434
rect 14822 9382 14874 9434
rect 14874 9382 14876 9434
rect 14820 9380 14876 9382
rect 14924 9434 14980 9436
rect 14924 9382 14926 9434
rect 14926 9382 14978 9434
rect 14978 9382 14980 9434
rect 14924 9380 14980 9382
rect 15028 9434 15084 9436
rect 15028 9382 15030 9434
rect 15030 9382 15082 9434
rect 15082 9382 15084 9434
rect 15028 9380 15084 9382
rect 15932 9042 15988 9044
rect 15932 8990 15934 9042
rect 15934 8990 15986 9042
rect 15986 8990 15988 9042
rect 15932 8988 15988 8990
rect 14140 8764 14196 8820
rect 15372 8876 15428 8932
rect 14924 8258 14980 8260
rect 14924 8206 14926 8258
rect 14926 8206 14978 8258
rect 14978 8206 14980 8258
rect 14924 8204 14980 8206
rect 16156 8764 16212 8820
rect 17948 8316 18004 8372
rect 17276 8204 17332 8260
rect 18222 10218 18278 10220
rect 18222 10166 18224 10218
rect 18224 10166 18276 10218
rect 18276 10166 18278 10218
rect 18222 10164 18278 10166
rect 18326 10218 18382 10220
rect 18326 10166 18328 10218
rect 18328 10166 18380 10218
rect 18380 10166 18382 10218
rect 18326 10164 18382 10166
rect 18430 10218 18486 10220
rect 18430 10166 18432 10218
rect 18432 10166 18484 10218
rect 18484 10166 18486 10218
rect 18430 10164 18486 10166
rect 20748 9772 20804 9828
rect 19068 8876 19124 8932
rect 19292 9100 19348 9156
rect 18222 8650 18278 8652
rect 18222 8598 18224 8650
rect 18224 8598 18276 8650
rect 18276 8598 18278 8650
rect 18222 8596 18278 8598
rect 18326 8650 18382 8652
rect 18326 8598 18328 8650
rect 18328 8598 18380 8650
rect 18380 8598 18382 8650
rect 18326 8596 18382 8598
rect 18430 8650 18486 8652
rect 18430 8598 18432 8650
rect 18432 8598 18484 8650
rect 18484 8598 18486 8650
rect 18430 8596 18486 8598
rect 20188 9154 20244 9156
rect 20188 9102 20190 9154
rect 20190 9102 20242 9154
rect 20242 9102 20244 9154
rect 20188 9100 20244 9102
rect 20412 8988 20468 9044
rect 19516 8316 19572 8372
rect 18508 8204 18564 8260
rect 14476 7868 14532 7924
rect 11418 7082 11474 7084
rect 11418 7030 11420 7082
rect 11420 7030 11472 7082
rect 11472 7030 11474 7082
rect 11418 7028 11474 7030
rect 11522 7082 11578 7084
rect 11522 7030 11524 7082
rect 11524 7030 11576 7082
rect 11576 7030 11578 7082
rect 11522 7028 11578 7030
rect 11626 7082 11682 7084
rect 11626 7030 11628 7082
rect 11628 7030 11680 7082
rect 11680 7030 11682 7082
rect 11626 7028 11682 7030
rect 11228 6748 11284 6804
rect 14820 7866 14876 7868
rect 14820 7814 14822 7866
rect 14822 7814 14874 7866
rect 14874 7814 14876 7866
rect 14820 7812 14876 7814
rect 14924 7866 14980 7868
rect 14924 7814 14926 7866
rect 14926 7814 14978 7866
rect 14978 7814 14980 7866
rect 14924 7812 14980 7814
rect 15028 7866 15084 7868
rect 15028 7814 15030 7866
rect 15030 7814 15082 7866
rect 15082 7814 15084 7866
rect 15028 7812 15084 7814
rect 19068 8092 19124 8148
rect 18508 7698 18564 7700
rect 18508 7646 18510 7698
rect 18510 7646 18562 7698
rect 18562 7646 18564 7698
rect 18508 7644 18564 7646
rect 19292 7644 19348 7700
rect 17276 6802 17332 6804
rect 17276 6750 17278 6802
rect 17278 6750 17330 6802
rect 17330 6750 17332 6802
rect 17276 6748 17332 6750
rect 18222 7082 18278 7084
rect 18222 7030 18224 7082
rect 18224 7030 18276 7082
rect 18276 7030 18278 7082
rect 18222 7028 18278 7030
rect 18326 7082 18382 7084
rect 18326 7030 18328 7082
rect 18328 7030 18380 7082
rect 18380 7030 18382 7082
rect 18326 7028 18382 7030
rect 18430 7082 18486 7084
rect 18430 7030 18432 7082
rect 18432 7030 18484 7082
rect 18484 7030 18486 7082
rect 18430 7028 18486 7030
rect 18060 6636 18116 6692
rect 18620 6860 18676 6916
rect 14252 6524 14308 6580
rect 15484 6578 15540 6580
rect 15484 6526 15486 6578
rect 15486 6526 15538 6578
rect 15538 6526 15540 6578
rect 15484 6524 15540 6526
rect 14820 6298 14876 6300
rect 14820 6246 14822 6298
rect 14822 6246 14874 6298
rect 14874 6246 14876 6298
rect 14820 6244 14876 6246
rect 14924 6298 14980 6300
rect 14924 6246 14926 6298
rect 14926 6246 14978 6298
rect 14978 6246 14980 6298
rect 14924 6244 14980 6246
rect 15028 6298 15084 6300
rect 15028 6246 15030 6298
rect 15030 6246 15082 6298
rect 15082 6246 15084 6298
rect 15028 6244 15084 6246
rect 21532 9826 21588 9828
rect 21532 9774 21534 9826
rect 21534 9774 21586 9826
rect 21586 9774 21588 9826
rect 21532 9772 21588 9774
rect 21624 9434 21680 9436
rect 21624 9382 21626 9434
rect 21626 9382 21678 9434
rect 21678 9382 21680 9434
rect 21624 9380 21680 9382
rect 21728 9434 21784 9436
rect 21728 9382 21730 9434
rect 21730 9382 21782 9434
rect 21782 9382 21784 9434
rect 21728 9380 21784 9382
rect 21832 9434 21888 9436
rect 21832 9382 21834 9434
rect 21834 9382 21886 9434
rect 21886 9382 21888 9434
rect 21832 9380 21888 9382
rect 24332 11282 24388 11284
rect 24332 11230 24334 11282
rect 24334 11230 24386 11282
rect 24386 11230 24388 11282
rect 24332 11228 24388 11230
rect 24332 9772 24388 9828
rect 20748 7644 20804 7700
rect 20748 7308 20804 7364
rect 20972 7196 21028 7252
rect 23548 9100 23604 9156
rect 24108 8764 24164 8820
rect 21420 8092 21476 8148
rect 22988 8092 23044 8148
rect 21624 7866 21680 7868
rect 21624 7814 21626 7866
rect 21626 7814 21678 7866
rect 21678 7814 21680 7866
rect 21624 7812 21680 7814
rect 21728 7866 21784 7868
rect 21728 7814 21730 7866
rect 21730 7814 21782 7866
rect 21782 7814 21784 7866
rect 21728 7812 21784 7814
rect 21832 7866 21888 7868
rect 21832 7814 21834 7866
rect 21834 7814 21886 7866
rect 21886 7814 21888 7866
rect 21832 7812 21888 7814
rect 24444 11116 24500 11172
rect 26236 13634 26292 13636
rect 26236 13582 26238 13634
rect 26238 13582 26290 13634
rect 26290 13582 26292 13634
rect 26236 13580 26292 13582
rect 26348 13468 26404 13524
rect 25026 11786 25082 11788
rect 25026 11734 25028 11786
rect 25028 11734 25080 11786
rect 25080 11734 25082 11786
rect 25026 11732 25082 11734
rect 25130 11786 25186 11788
rect 25130 11734 25132 11786
rect 25132 11734 25184 11786
rect 25184 11734 25186 11786
rect 25130 11732 25186 11734
rect 25234 11786 25290 11788
rect 25234 11734 25236 11786
rect 25236 11734 25288 11786
rect 25288 11734 25290 11786
rect 25234 11732 25290 11734
rect 24556 10556 24612 10612
rect 25026 10218 25082 10220
rect 25026 10166 25028 10218
rect 25028 10166 25080 10218
rect 25080 10166 25082 10218
rect 25026 10164 25082 10166
rect 25130 10218 25186 10220
rect 25130 10166 25132 10218
rect 25132 10166 25184 10218
rect 25184 10166 25186 10218
rect 25130 10164 25186 10166
rect 25234 10218 25290 10220
rect 25234 10166 25236 10218
rect 25236 10166 25288 10218
rect 25288 10166 25290 10218
rect 25234 10164 25290 10166
rect 24668 9042 24724 9044
rect 24668 8990 24670 9042
rect 24670 8990 24722 9042
rect 24722 8990 24724 9042
rect 24668 8988 24724 8990
rect 24332 8092 24388 8148
rect 26124 11900 26180 11956
rect 25340 8988 25396 9044
rect 26236 10498 26292 10500
rect 26236 10446 26238 10498
rect 26238 10446 26290 10498
rect 26290 10446 26292 10498
rect 26236 10444 26292 10446
rect 28428 14138 28484 14140
rect 28428 14086 28430 14138
rect 28430 14086 28482 14138
rect 28482 14086 28484 14138
rect 28428 14084 28484 14086
rect 28532 14138 28588 14140
rect 28532 14086 28534 14138
rect 28534 14086 28586 14138
rect 28586 14086 28588 14138
rect 28532 14084 28588 14086
rect 28636 14138 28692 14140
rect 28636 14086 28638 14138
rect 28638 14086 28690 14138
rect 28690 14086 28692 14138
rect 28636 14084 28692 14086
rect 28428 12570 28484 12572
rect 28428 12518 28430 12570
rect 28430 12518 28482 12570
rect 28482 12518 28484 12570
rect 28428 12516 28484 12518
rect 28532 12570 28588 12572
rect 28532 12518 28534 12570
rect 28534 12518 28586 12570
rect 28586 12518 28588 12570
rect 28532 12516 28588 12518
rect 28636 12570 28692 12572
rect 28636 12518 28638 12570
rect 28638 12518 28690 12570
rect 28690 12518 28692 12570
rect 28636 12516 28692 12518
rect 26684 12236 26740 12292
rect 27356 12290 27412 12292
rect 27356 12238 27358 12290
rect 27358 12238 27410 12290
rect 27410 12238 27412 12290
rect 27356 12236 27412 12238
rect 26908 11170 26964 11172
rect 26908 11118 26910 11170
rect 26910 11118 26962 11170
rect 26962 11118 26964 11170
rect 26908 11116 26964 11118
rect 27244 10722 27300 10724
rect 27244 10670 27246 10722
rect 27246 10670 27298 10722
rect 27298 10670 27300 10722
rect 27244 10668 27300 10670
rect 28428 11002 28484 11004
rect 28428 10950 28430 11002
rect 28430 10950 28482 11002
rect 28482 10950 28484 11002
rect 28428 10948 28484 10950
rect 28532 11002 28588 11004
rect 28532 10950 28534 11002
rect 28534 10950 28586 11002
rect 28586 10950 28588 11002
rect 28532 10948 28588 10950
rect 28636 11002 28692 11004
rect 28636 10950 28638 11002
rect 28638 10950 28690 11002
rect 28690 10950 28692 11002
rect 28636 10948 28692 10950
rect 27356 10556 27412 10612
rect 26684 9884 26740 9940
rect 25026 8650 25082 8652
rect 25026 8598 25028 8650
rect 25028 8598 25080 8650
rect 25080 8598 25082 8650
rect 25026 8596 25082 8598
rect 25130 8650 25186 8652
rect 25130 8598 25132 8650
rect 25132 8598 25184 8650
rect 25184 8598 25186 8650
rect 25130 8596 25186 8598
rect 25234 8650 25290 8652
rect 25234 8598 25236 8650
rect 25236 8598 25288 8650
rect 25288 8598 25290 8650
rect 25234 8596 25290 8598
rect 25452 8428 25508 8484
rect 26460 8764 26516 8820
rect 24892 7532 24948 7588
rect 25788 7980 25844 8036
rect 21084 6860 21140 6916
rect 22652 7308 22708 7364
rect 20300 6636 20356 6692
rect 23324 7362 23380 7364
rect 23324 7310 23326 7362
rect 23326 7310 23378 7362
rect 23378 7310 23380 7362
rect 23324 7308 23380 7310
rect 22988 6748 23044 6804
rect 23100 7196 23156 7252
rect 21624 6298 21680 6300
rect 21624 6246 21626 6298
rect 21626 6246 21678 6298
rect 21678 6246 21680 6298
rect 21624 6244 21680 6246
rect 21728 6298 21784 6300
rect 21728 6246 21730 6298
rect 21730 6246 21782 6298
rect 21782 6246 21784 6298
rect 21728 6244 21784 6246
rect 21832 6298 21888 6300
rect 21832 6246 21834 6298
rect 21834 6246 21886 6298
rect 21886 6246 21888 6298
rect 21832 6244 21888 6246
rect 19964 5740 20020 5796
rect 22092 5794 22148 5796
rect 22092 5742 22094 5794
rect 22094 5742 22146 5794
rect 22146 5742 22148 5794
rect 22092 5740 22148 5742
rect 11418 5514 11474 5516
rect 11418 5462 11420 5514
rect 11420 5462 11472 5514
rect 11472 5462 11474 5514
rect 11418 5460 11474 5462
rect 11522 5514 11578 5516
rect 11522 5462 11524 5514
rect 11524 5462 11576 5514
rect 11576 5462 11578 5514
rect 11522 5460 11578 5462
rect 11626 5514 11682 5516
rect 11626 5462 11628 5514
rect 11628 5462 11680 5514
rect 11680 5462 11682 5514
rect 11626 5460 11682 5462
rect 18222 5514 18278 5516
rect 18222 5462 18224 5514
rect 18224 5462 18276 5514
rect 18276 5462 18278 5514
rect 18222 5460 18278 5462
rect 18326 5514 18382 5516
rect 18326 5462 18328 5514
rect 18328 5462 18380 5514
rect 18380 5462 18382 5514
rect 18326 5460 18382 5462
rect 18430 5514 18486 5516
rect 18430 5462 18432 5514
rect 18432 5462 18484 5514
rect 18484 5462 18486 5514
rect 18430 5460 18486 5462
rect 8540 5068 8596 5124
rect 8016 4730 8072 4732
rect 8016 4678 8018 4730
rect 8018 4678 8070 4730
rect 8070 4678 8072 4730
rect 8016 4676 8072 4678
rect 8120 4730 8176 4732
rect 8120 4678 8122 4730
rect 8122 4678 8174 4730
rect 8174 4678 8176 4730
rect 8120 4676 8176 4678
rect 8224 4730 8280 4732
rect 8224 4678 8226 4730
rect 8226 4678 8278 4730
rect 8278 4678 8280 4730
rect 8224 4676 8280 4678
rect 4614 3946 4670 3948
rect 4614 3894 4616 3946
rect 4616 3894 4668 3946
rect 4668 3894 4670 3946
rect 4614 3892 4670 3894
rect 4718 3946 4774 3948
rect 4718 3894 4720 3946
rect 4720 3894 4772 3946
rect 4772 3894 4774 3946
rect 4718 3892 4774 3894
rect 4822 3946 4878 3948
rect 4822 3894 4824 3946
rect 4824 3894 4876 3946
rect 4876 3894 4878 3946
rect 4822 3892 4878 3894
rect 10556 5068 10612 5124
rect 9100 4226 9156 4228
rect 9100 4174 9102 4226
rect 9102 4174 9154 4226
rect 9154 4174 9156 4226
rect 9100 4172 9156 4174
rect 8016 3162 8072 3164
rect 8016 3110 8018 3162
rect 8018 3110 8070 3162
rect 8070 3110 8072 3162
rect 8016 3108 8072 3110
rect 8120 3162 8176 3164
rect 8120 3110 8122 3162
rect 8122 3110 8174 3162
rect 8174 3110 8176 3162
rect 8120 3108 8176 3110
rect 8224 3162 8280 3164
rect 8224 3110 8226 3162
rect 8226 3110 8278 3162
rect 8278 3110 8280 3162
rect 8224 3108 8280 3110
rect 10556 4172 10612 4228
rect 12236 4508 12292 4564
rect 11116 3276 11172 3332
rect 11418 3946 11474 3948
rect 11418 3894 11420 3946
rect 11420 3894 11472 3946
rect 11472 3894 11474 3946
rect 11418 3892 11474 3894
rect 11522 3946 11578 3948
rect 11522 3894 11524 3946
rect 11524 3894 11576 3946
rect 11576 3894 11578 3946
rect 11522 3892 11578 3894
rect 11626 3946 11682 3948
rect 11626 3894 11628 3946
rect 11628 3894 11680 3946
rect 11680 3894 11682 3946
rect 11626 3892 11682 3894
rect 12684 5122 12740 5124
rect 12684 5070 12686 5122
rect 12686 5070 12738 5122
rect 12738 5070 12740 5122
rect 12684 5068 12740 5070
rect 18060 5068 18116 5124
rect 12908 4898 12964 4900
rect 12908 4846 12910 4898
rect 12910 4846 12962 4898
rect 12962 4846 12964 4898
rect 12908 4844 12964 4846
rect 14476 5010 14532 5012
rect 14476 4958 14478 5010
rect 14478 4958 14530 5010
rect 14530 4958 14532 5010
rect 14476 4956 14532 4958
rect 15260 4956 15316 5012
rect 13468 4396 13524 4452
rect 13580 4844 13636 4900
rect 12684 3388 12740 3444
rect 11564 3330 11620 3332
rect 11564 3278 11566 3330
rect 11566 3278 11618 3330
rect 11618 3278 11620 3330
rect 11564 3276 11620 3278
rect 13804 4898 13860 4900
rect 13804 4846 13806 4898
rect 13806 4846 13858 4898
rect 13858 4846 13860 4898
rect 13804 4844 13860 4846
rect 13692 4562 13748 4564
rect 13692 4510 13694 4562
rect 13694 4510 13746 4562
rect 13746 4510 13748 4562
rect 13692 4508 13748 4510
rect 13244 3442 13300 3444
rect 13244 3390 13246 3442
rect 13246 3390 13298 3442
rect 13298 3390 13300 3442
rect 13244 3388 13300 3390
rect 15148 4844 15204 4900
rect 14820 4730 14876 4732
rect 14820 4678 14822 4730
rect 14822 4678 14874 4730
rect 14874 4678 14876 4730
rect 14820 4676 14876 4678
rect 14924 4730 14980 4732
rect 14924 4678 14926 4730
rect 14926 4678 14978 4730
rect 14978 4678 14980 4730
rect 14924 4676 14980 4678
rect 15028 4730 15084 4732
rect 15028 4678 15030 4730
rect 15030 4678 15082 4730
rect 15082 4678 15084 4730
rect 15028 4676 15084 4678
rect 14700 3500 14756 3556
rect 14924 4338 14980 4340
rect 14924 4286 14926 4338
rect 14926 4286 14978 4338
rect 14978 4286 14980 4338
rect 14924 4284 14980 4286
rect 17388 4450 17444 4452
rect 17388 4398 17390 4450
rect 17390 4398 17442 4450
rect 17442 4398 17444 4450
rect 17388 4396 17444 4398
rect 15596 4338 15652 4340
rect 15596 4286 15598 4338
rect 15598 4286 15650 4338
rect 15650 4286 15652 4338
rect 15596 4284 15652 4286
rect 14820 3162 14876 3164
rect 14820 3110 14822 3162
rect 14822 3110 14874 3162
rect 14874 3110 14876 3162
rect 14820 3108 14876 3110
rect 14924 3162 14980 3164
rect 14924 3110 14926 3162
rect 14926 3110 14978 3162
rect 14978 3110 14980 3162
rect 14924 3108 14980 3110
rect 15028 3162 15084 3164
rect 15028 3110 15030 3162
rect 15030 3110 15082 3162
rect 15082 3110 15084 3162
rect 15028 3108 15084 3110
rect 16156 3612 16212 3668
rect 17388 3666 17444 3668
rect 17388 3614 17390 3666
rect 17390 3614 17442 3666
rect 17442 3614 17444 3666
rect 17388 3612 17444 3614
rect 16940 3554 16996 3556
rect 16940 3502 16942 3554
rect 16942 3502 16994 3554
rect 16994 3502 16996 3554
rect 16940 3500 16996 3502
rect 18222 3946 18278 3948
rect 18222 3894 18224 3946
rect 18224 3894 18276 3946
rect 18276 3894 18278 3946
rect 18222 3892 18278 3894
rect 18326 3946 18382 3948
rect 18326 3894 18328 3946
rect 18328 3894 18380 3946
rect 18380 3894 18382 3946
rect 18326 3892 18382 3894
rect 18430 3946 18486 3948
rect 18430 3894 18432 3946
rect 18432 3894 18484 3946
rect 18484 3894 18486 3946
rect 18430 3892 18486 3894
rect 18396 3442 18452 3444
rect 18396 3390 18398 3442
rect 18398 3390 18450 3442
rect 18450 3390 18452 3442
rect 18396 3388 18452 3390
rect 19068 3388 19124 3444
rect 21084 3724 21140 3780
rect 23324 6860 23380 6916
rect 24220 6076 24276 6132
rect 23100 5740 23156 5796
rect 23212 5180 23268 5236
rect 21532 4844 21588 4900
rect 21624 4730 21680 4732
rect 21624 4678 21626 4730
rect 21626 4678 21678 4730
rect 21678 4678 21680 4730
rect 21624 4676 21680 4678
rect 21728 4730 21784 4732
rect 21728 4678 21730 4730
rect 21730 4678 21782 4730
rect 21782 4678 21784 4730
rect 21728 4676 21784 4678
rect 21832 4730 21888 4732
rect 21832 4678 21834 4730
rect 21834 4678 21886 4730
rect 21886 4678 21888 4730
rect 21832 4676 21888 4678
rect 22204 4620 22260 4676
rect 23100 4508 23156 4564
rect 22428 4450 22484 4452
rect 22428 4398 22430 4450
rect 22430 4398 22482 4450
rect 22482 4398 22484 4450
rect 22428 4396 22484 4398
rect 21756 4060 21812 4116
rect 22876 4060 22932 4116
rect 21532 3388 21588 3444
rect 22428 3612 22484 3668
rect 25026 7082 25082 7084
rect 25026 7030 25028 7082
rect 25028 7030 25080 7082
rect 25080 7030 25082 7082
rect 25026 7028 25082 7030
rect 25130 7082 25186 7084
rect 25130 7030 25132 7082
rect 25132 7030 25184 7082
rect 25184 7030 25186 7082
rect 25130 7028 25186 7030
rect 25234 7082 25290 7084
rect 25234 7030 25236 7082
rect 25236 7030 25288 7082
rect 25288 7030 25290 7082
rect 25234 7028 25290 7030
rect 25676 6636 25732 6692
rect 24668 6018 24724 6020
rect 24668 5966 24670 6018
rect 24670 5966 24722 6018
rect 24722 5966 24724 6018
rect 24668 5964 24724 5966
rect 25026 5514 25082 5516
rect 25026 5462 25028 5514
rect 25028 5462 25080 5514
rect 25080 5462 25082 5514
rect 25026 5460 25082 5462
rect 25130 5514 25186 5516
rect 25130 5462 25132 5514
rect 25132 5462 25184 5514
rect 25184 5462 25186 5514
rect 25130 5460 25186 5462
rect 25234 5514 25290 5516
rect 25234 5462 25236 5514
rect 25236 5462 25288 5514
rect 25288 5462 25290 5514
rect 25234 5460 25290 5462
rect 24556 5292 24612 5348
rect 25340 5292 25396 5348
rect 24332 5068 24388 5124
rect 24780 4562 24836 4564
rect 24780 4510 24782 4562
rect 24782 4510 24834 4562
rect 24834 4510 24836 4562
rect 24780 4508 24836 4510
rect 23436 4450 23492 4452
rect 23436 4398 23438 4450
rect 23438 4398 23490 4450
rect 23490 4398 23492 4450
rect 23436 4396 23492 4398
rect 24668 4060 24724 4116
rect 25026 3946 25082 3948
rect 25026 3894 25028 3946
rect 25028 3894 25080 3946
rect 25080 3894 25082 3946
rect 25026 3892 25082 3894
rect 25130 3946 25186 3948
rect 25130 3894 25132 3946
rect 25132 3894 25184 3946
rect 25184 3894 25186 3946
rect 25130 3892 25186 3894
rect 25234 3946 25290 3948
rect 25234 3894 25236 3946
rect 25236 3894 25288 3946
rect 25288 3894 25290 3946
rect 25234 3892 25290 3894
rect 24668 3666 24724 3668
rect 24668 3614 24670 3666
rect 24670 3614 24722 3666
rect 24722 3614 24724 3666
rect 24668 3612 24724 3614
rect 25004 3724 25060 3780
rect 26236 6860 26292 6916
rect 26124 6412 26180 6468
rect 26236 5794 26292 5796
rect 26236 5742 26238 5794
rect 26238 5742 26290 5794
rect 26290 5742 26292 5794
rect 26236 5740 26292 5742
rect 26348 4396 26404 4452
rect 27244 9154 27300 9156
rect 27244 9102 27246 9154
rect 27246 9102 27298 9154
rect 27298 9102 27300 9154
rect 27244 9100 27300 9102
rect 27132 8428 27188 8484
rect 27468 9938 27524 9940
rect 27468 9886 27470 9938
rect 27470 9886 27522 9938
rect 27522 9886 27524 9938
rect 27468 9884 27524 9886
rect 28428 9434 28484 9436
rect 28428 9382 28430 9434
rect 28430 9382 28482 9434
rect 28482 9382 28484 9434
rect 28428 9380 28484 9382
rect 28532 9434 28588 9436
rect 28532 9382 28534 9434
rect 28534 9382 28586 9434
rect 28586 9382 28588 9434
rect 28532 9380 28588 9382
rect 28636 9434 28692 9436
rect 28636 9382 28638 9434
rect 28638 9382 28690 9434
rect 28690 9382 28692 9434
rect 28636 9380 28692 9382
rect 27692 8764 27748 8820
rect 27468 8092 27524 8148
rect 27580 8034 27636 8036
rect 27580 7982 27582 8034
rect 27582 7982 27634 8034
rect 27634 7982 27636 8034
rect 27580 7980 27636 7982
rect 27244 7586 27300 7588
rect 27244 7534 27246 7586
rect 27246 7534 27298 7586
rect 27298 7534 27300 7586
rect 27244 7532 27300 7534
rect 27356 7420 27412 7476
rect 27244 6748 27300 6804
rect 26908 6466 26964 6468
rect 26908 6414 26910 6466
rect 26910 6414 26962 6466
rect 26962 6414 26964 6466
rect 26908 6412 26964 6414
rect 26908 5964 26964 6020
rect 26572 4620 26628 4676
rect 24108 3442 24164 3444
rect 24108 3390 24110 3442
rect 24110 3390 24162 3442
rect 24162 3390 24164 3442
rect 24108 3388 24164 3390
rect 21624 3162 21680 3164
rect 21624 3110 21626 3162
rect 21626 3110 21678 3162
rect 21678 3110 21680 3162
rect 21624 3108 21680 3110
rect 21728 3162 21784 3164
rect 21728 3110 21730 3162
rect 21730 3110 21782 3162
rect 21782 3110 21784 3162
rect 21728 3108 21784 3110
rect 21832 3162 21888 3164
rect 21832 3110 21834 3162
rect 21834 3110 21886 3162
rect 21886 3110 21888 3162
rect 21832 3108 21888 3110
rect 20860 2716 20916 2772
rect 20188 2044 20244 2100
rect 28140 8428 28196 8484
rect 27804 8092 27860 8148
rect 28428 7866 28484 7868
rect 28428 7814 28430 7866
rect 28430 7814 28482 7866
rect 28482 7814 28484 7866
rect 28428 7812 28484 7814
rect 28532 7866 28588 7868
rect 28532 7814 28534 7866
rect 28534 7814 28586 7866
rect 28586 7814 28588 7866
rect 28532 7812 28588 7814
rect 28636 7866 28692 7868
rect 28636 7814 28638 7866
rect 28638 7814 28690 7866
rect 28690 7814 28692 7866
rect 28636 7812 28692 7814
rect 28428 6298 28484 6300
rect 28428 6246 28430 6298
rect 28430 6246 28482 6298
rect 28482 6246 28484 6298
rect 28428 6244 28484 6246
rect 28532 6298 28588 6300
rect 28532 6246 28534 6298
rect 28534 6246 28586 6298
rect 28586 6246 28588 6298
rect 28532 6244 28588 6246
rect 28636 6298 28692 6300
rect 28636 6246 28638 6298
rect 28638 6246 28690 6298
rect 28690 6246 28692 6298
rect 28636 6244 28692 6246
rect 28428 4730 28484 4732
rect 28428 4678 28430 4730
rect 28430 4678 28482 4730
rect 28482 4678 28484 4730
rect 28428 4676 28484 4678
rect 28532 4730 28588 4732
rect 28532 4678 28534 4730
rect 28534 4678 28586 4730
rect 28586 4678 28588 4730
rect 28532 4676 28588 4678
rect 28636 4730 28692 4732
rect 28636 4678 28638 4730
rect 28638 4678 28690 4730
rect 28690 4678 28692 4730
rect 28636 4676 28692 4678
rect 27468 4450 27524 4452
rect 27468 4398 27470 4450
rect 27470 4398 27522 4450
rect 27522 4398 27524 4450
rect 27468 4396 27524 4398
rect 28428 3162 28484 3164
rect 28428 3110 28430 3162
rect 28430 3110 28482 3162
rect 28482 3110 28484 3162
rect 28428 3108 28484 3110
rect 28532 3162 28588 3164
rect 28532 3110 28534 3162
rect 28534 3110 28586 3162
rect 28586 3110 28588 3162
rect 28532 3108 28588 3110
rect 28636 3162 28692 3164
rect 28636 3110 28638 3162
rect 28638 3110 28690 3162
rect 28690 3110 28692 3162
rect 28636 3108 28692 3110
rect 26684 1372 26740 1428
<< metal3 >>
rect 29200 29652 30000 29680
rect 24434 29596 24444 29652
rect 24500 29596 30000 29652
rect 29200 29568 30000 29596
rect 29200 28980 30000 29008
rect 27794 28924 27804 28980
rect 27860 28924 30000 28980
rect 29200 28896 30000 28924
rect 29200 28308 30000 28336
rect 25106 28252 25116 28308
rect 25172 28252 30000 28308
rect 29200 28224 30000 28252
rect 29200 27636 30000 27664
rect 27458 27580 27468 27636
rect 27524 27580 30000 27636
rect 29200 27552 30000 27580
rect 29200 26964 30000 26992
rect 25890 26908 25900 26964
rect 25956 26908 30000 26964
rect 29200 26880 30000 26908
rect 17490 26796 17500 26852
rect 17556 26796 18956 26852
rect 19012 26796 19022 26852
rect 21522 26796 21532 26852
rect 21588 26796 22764 26852
rect 22820 26796 22830 26852
rect 22978 26796 22988 26852
rect 23044 26796 25004 26852
rect 25060 26796 25070 26852
rect 8006 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8290 26684
rect 14810 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15094 26684
rect 21614 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21898 26684
rect 28418 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28702 26684
rect 18162 26572 18172 26628
rect 18228 26572 18844 26628
rect 18900 26572 18910 26628
rect 16146 26460 16156 26516
rect 16212 26460 17388 26516
rect 17444 26460 17454 26516
rect 24882 26460 24892 26516
rect 24948 26460 26124 26516
rect 26180 26460 26190 26516
rect 29200 26292 30000 26320
rect 3378 26236 3388 26292
rect 3444 26236 9548 26292
rect 9604 26236 9614 26292
rect 26114 26236 26124 26292
rect 26180 26236 30000 26292
rect 29200 26208 30000 26236
rect 4274 26124 4284 26180
rect 4340 26124 10668 26180
rect 10724 26124 10734 26180
rect 11442 26012 11452 26068
rect 11508 26012 12124 26068
rect 12180 26012 12190 26068
rect 4604 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4888 25900
rect 11408 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11692 25900
rect 18212 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18496 25900
rect 25016 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25300 25900
rect 15922 25788 15932 25844
rect 15988 25788 16940 25844
rect 16996 25788 17006 25844
rect 3938 25676 3948 25732
rect 4004 25676 9212 25732
rect 9268 25676 9278 25732
rect 12786 25676 12796 25732
rect 12852 25676 13916 25732
rect 13972 25676 13982 25732
rect 29200 25620 30000 25648
rect 6066 25564 6076 25620
rect 6132 25564 6972 25620
rect 7028 25564 7038 25620
rect 7298 25564 7308 25620
rect 7364 25564 10780 25620
rect 10836 25564 10846 25620
rect 19618 25564 19628 25620
rect 19684 25564 20188 25620
rect 20244 25564 20254 25620
rect 27682 25564 27692 25620
rect 27748 25564 30000 25620
rect 29200 25536 30000 25564
rect 6626 25452 6636 25508
rect 6692 25452 9772 25508
rect 9828 25452 9838 25508
rect 9986 25452 9996 25508
rect 10052 25452 11788 25508
rect 11844 25452 11854 25508
rect 15260 25452 18508 25508
rect 18564 25452 18574 25508
rect 7970 25340 7980 25396
rect 8036 25340 11900 25396
rect 11956 25340 11966 25396
rect 15260 25284 15316 25452
rect 16818 25340 16828 25396
rect 16884 25340 18620 25396
rect 18676 25340 18686 25396
rect 20738 25340 20748 25396
rect 20804 25340 24556 25396
rect 24612 25340 24622 25396
rect 2146 25228 2156 25284
rect 2212 25228 2222 25284
rect 2930 25228 2940 25284
rect 2996 25228 3500 25284
rect 3556 25228 3566 25284
rect 4610 25228 4620 25284
rect 4676 25228 8428 25284
rect 8484 25228 8494 25284
rect 9314 25228 9324 25284
rect 9380 25228 11060 25284
rect 15250 25228 15260 25284
rect 15316 25228 15326 25284
rect 16482 25228 16492 25284
rect 16548 25228 17052 25284
rect 17108 25228 17118 25284
rect 20514 25228 20524 25284
rect 20580 25228 23996 25284
rect 24052 25228 24062 25284
rect 24210 25228 24220 25284
rect 24276 25228 24668 25284
rect 24724 25228 24734 25284
rect 25554 25228 25564 25284
rect 25620 25228 26908 25284
rect 26964 25228 26974 25284
rect 0 24948 800 24976
rect 2156 24948 2212 25228
rect 2706 25116 2716 25172
rect 2772 25116 4284 25172
rect 4340 25116 4350 25172
rect 8006 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8290 25116
rect 11004 25060 11060 25228
rect 23090 25116 23100 25172
rect 23156 25116 23660 25172
rect 23716 25116 24444 25172
rect 24500 25116 24510 25172
rect 14810 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15094 25116
rect 21614 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21898 25116
rect 28418 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28702 25116
rect 10994 25004 11004 25060
rect 11060 25004 11070 25060
rect 29200 24948 30000 24976
rect 0 24892 2212 24948
rect 9426 24892 9436 24948
rect 9492 24892 10444 24948
rect 10500 24892 10510 24948
rect 23762 24892 23772 24948
rect 23828 24892 25452 24948
rect 25508 24892 25518 24948
rect 27682 24892 27692 24948
rect 27748 24892 30000 24948
rect 0 24864 800 24892
rect 29200 24864 30000 24892
rect 8866 24780 8876 24836
rect 8932 24780 9660 24836
rect 9716 24780 9726 24836
rect 23986 24780 23996 24836
rect 24052 24780 25900 24836
rect 25956 24780 25966 24836
rect 20850 24668 20860 24724
rect 20916 24668 22540 24724
rect 22596 24668 22606 24724
rect 22754 24556 22764 24612
rect 22820 24556 24668 24612
rect 24724 24556 24734 24612
rect 10882 24444 10892 24500
rect 10948 24444 11340 24500
rect 11396 24444 11406 24500
rect 0 24276 800 24304
rect 4604 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4888 24332
rect 11408 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11692 24332
rect 18212 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18496 24332
rect 25016 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25300 24332
rect 29200 24276 30000 24304
rect 0 24220 2380 24276
rect 2436 24220 2446 24276
rect 28018 24220 28028 24276
rect 28084 24220 30000 24276
rect 0 24192 800 24220
rect 29200 24192 30000 24220
rect 2034 24108 2044 24164
rect 2100 24108 9660 24164
rect 9716 24108 9726 24164
rect 24210 24108 24220 24164
rect 24276 24108 26908 24164
rect 26964 24108 26974 24164
rect 23314 23884 23324 23940
rect 23380 23884 25228 23940
rect 25284 23884 25294 23940
rect 2034 23772 2044 23828
rect 2100 23772 3724 23828
rect 3780 23772 3790 23828
rect 6850 23772 6860 23828
rect 6916 23772 11676 23828
rect 11732 23772 11742 23828
rect 24658 23772 24668 23828
rect 24724 23772 28868 23828
rect 25778 23660 25788 23716
rect 25844 23660 26908 23716
rect 26964 23660 26974 23716
rect 0 23604 800 23632
rect 28812 23604 28868 23772
rect 29200 23604 30000 23632
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 28812 23548 30000 23604
rect 0 23520 800 23548
rect 8006 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8290 23548
rect 14810 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15094 23548
rect 21614 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21898 23548
rect 28418 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28702 23548
rect 29200 23520 30000 23548
rect 10546 23436 10556 23492
rect 10612 23436 13356 23492
rect 13412 23436 13422 23492
rect 4946 23212 4956 23268
rect 5012 23212 10220 23268
rect 10276 23212 10286 23268
rect 20626 23212 20636 23268
rect 20692 23212 24220 23268
rect 24276 23212 24286 23268
rect 24658 23212 24668 23268
rect 24724 23212 26908 23268
rect 26964 23212 26974 23268
rect 29200 22932 30000 22960
rect 26786 22876 26796 22932
rect 26852 22876 30000 22932
rect 29200 22848 30000 22876
rect 26226 22764 26236 22820
rect 26292 22764 26908 22820
rect 26964 22764 26974 22820
rect 4604 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4888 22764
rect 11408 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11692 22764
rect 18212 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18496 22764
rect 25016 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25300 22764
rect 29200 22260 30000 22288
rect 28018 22204 28028 22260
rect 28084 22204 30000 22260
rect 29200 22176 30000 22204
rect 8006 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8290 21980
rect 14810 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15094 21980
rect 21614 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21898 21980
rect 28418 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28702 21980
rect 26226 21756 26236 21812
rect 26292 21756 27804 21812
rect 27860 21756 27870 21812
rect 13010 21644 13020 21700
rect 13076 21644 14812 21700
rect 14868 21644 14878 21700
rect 24434 21644 24444 21700
rect 24500 21644 27132 21700
rect 27188 21644 27198 21700
rect 29200 21588 30000 21616
rect 26674 21532 26684 21588
rect 26740 21532 27468 21588
rect 27524 21532 30000 21588
rect 29200 21504 30000 21532
rect 12338 21420 12348 21476
rect 12404 21420 13804 21476
rect 13860 21420 13870 21476
rect 26226 21420 26236 21476
rect 26292 21420 26796 21476
rect 26852 21420 26862 21476
rect 25778 21196 25788 21252
rect 25844 21196 27468 21252
rect 27524 21196 27534 21252
rect 4604 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4888 21196
rect 11408 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11692 21196
rect 18212 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18496 21196
rect 25016 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25300 21196
rect 29200 20916 30000 20944
rect 22866 20860 22876 20916
rect 22932 20860 24444 20916
rect 24500 20860 24510 20916
rect 28130 20860 28140 20916
rect 28196 20860 30000 20916
rect 29200 20832 30000 20860
rect 25890 20748 25900 20804
rect 25956 20748 26908 20804
rect 26964 20748 26974 20804
rect 15362 20636 15372 20692
rect 15428 20636 17276 20692
rect 17332 20636 17342 20692
rect 8006 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8290 20412
rect 14810 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15094 20412
rect 21614 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21898 20412
rect 28418 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28702 20412
rect 29200 20244 30000 20272
rect 14914 20188 14924 20244
rect 14980 20188 16268 20244
rect 16324 20188 16334 20244
rect 28018 20188 28028 20244
rect 28084 20188 30000 20244
rect 29200 20160 30000 20188
rect 24546 20076 24556 20132
rect 24612 20076 27804 20132
rect 27860 20076 27870 20132
rect 21074 19964 21084 20020
rect 21140 19964 23548 20020
rect 23604 19964 23614 20020
rect 23762 19964 23772 20020
rect 23828 19964 25340 20020
rect 25396 19964 25406 20020
rect 20738 19852 20748 19908
rect 20804 19852 22316 19908
rect 22372 19852 22382 19908
rect 23986 19852 23996 19908
rect 24052 19852 26236 19908
rect 26292 19852 26302 19908
rect 8530 19740 8540 19796
rect 8596 19740 9548 19796
rect 9604 19740 9614 19796
rect 23202 19740 23212 19796
rect 23268 19740 24108 19796
rect 24164 19740 24174 19796
rect 0 19572 800 19600
rect 4604 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4888 19628
rect 11408 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11692 19628
rect 18212 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18496 19628
rect 25016 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25300 19628
rect 29200 19572 30000 19600
rect 0 19516 4284 19572
rect 4340 19516 4350 19572
rect 28130 19516 28140 19572
rect 28196 19516 30000 19572
rect 0 19488 800 19516
rect 29200 19488 30000 19516
rect 6066 19292 6076 19348
rect 6132 19292 7644 19348
rect 7700 19292 7710 19348
rect 18050 19292 18060 19348
rect 18116 19292 19180 19348
rect 19236 19292 19246 19348
rect 16370 19068 16380 19124
rect 16436 19068 17164 19124
rect 17220 19068 17230 19124
rect 17938 19068 17948 19124
rect 18004 19068 20188 19124
rect 20244 19068 20254 19124
rect 23874 18956 23884 19012
rect 23940 18956 26124 19012
rect 26180 18956 26190 19012
rect 27570 18956 27580 19012
rect 27636 18956 28140 19012
rect 28196 18956 28868 19012
rect 28812 18900 28868 18956
rect 29200 18900 30000 18928
rect 28812 18844 30000 18900
rect 8006 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8290 18844
rect 14810 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15094 18844
rect 21614 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21898 18844
rect 28418 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28702 18844
rect 29200 18816 30000 18844
rect 11218 18508 11228 18564
rect 11284 18508 12572 18564
rect 12628 18508 12638 18564
rect 13244 18508 14252 18564
rect 14308 18508 14318 18564
rect 16930 18508 16940 18564
rect 16996 18508 19404 18564
rect 19460 18508 19470 18564
rect 13244 18452 13300 18508
rect 9538 18396 9548 18452
rect 9604 18396 11900 18452
rect 11956 18396 12460 18452
rect 12516 18396 13244 18452
rect 13300 18396 13310 18452
rect 9986 18284 9996 18340
rect 10052 18284 11564 18340
rect 11620 18284 11630 18340
rect 21410 18284 21420 18340
rect 21476 18284 23100 18340
rect 23156 18284 24444 18340
rect 24500 18284 25340 18340
rect 25396 18284 26348 18340
rect 26404 18284 26414 18340
rect 29200 18228 30000 18256
rect 16930 18172 16940 18228
rect 16996 18172 18396 18228
rect 18452 18172 18462 18228
rect 27682 18172 27692 18228
rect 27748 18172 28140 18228
rect 28196 18172 30000 18228
rect 29200 18144 30000 18172
rect 4604 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4888 18060
rect 11408 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11692 18060
rect 18212 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18496 18060
rect 25016 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25300 18060
rect 5506 17612 5516 17668
rect 5572 17612 7532 17668
rect 7588 17612 9548 17668
rect 9604 17612 9614 17668
rect 9986 17612 9996 17668
rect 10052 17612 11676 17668
rect 11732 17612 13468 17668
rect 13524 17612 15708 17668
rect 15764 17612 15774 17668
rect 20626 17612 20636 17668
rect 20692 17612 21420 17668
rect 21476 17612 21486 17668
rect 26338 17612 26348 17668
rect 26404 17612 27132 17668
rect 27188 17612 27198 17668
rect 25554 17500 25564 17556
rect 25620 17500 27804 17556
rect 27860 17500 27870 17556
rect 4946 17388 4956 17444
rect 5012 17388 5628 17444
rect 5684 17388 6636 17444
rect 6692 17388 6702 17444
rect 12786 17388 12796 17444
rect 12852 17388 13804 17444
rect 13860 17388 13870 17444
rect 19282 17388 19292 17444
rect 19348 17388 20076 17444
rect 20132 17388 20142 17444
rect 8006 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8290 17276
rect 14810 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15094 17276
rect 21614 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21898 17276
rect 28418 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28702 17276
rect 21634 17052 21644 17108
rect 21700 17052 27244 17108
rect 27300 17052 27310 17108
rect 23314 16940 23324 16996
rect 23380 16940 23996 16996
rect 24052 16940 24062 16996
rect 3602 16828 3612 16884
rect 3668 16828 5068 16884
rect 5124 16828 5516 16884
rect 5572 16828 5582 16884
rect 16034 16828 16044 16884
rect 16100 16828 17612 16884
rect 17668 16828 17948 16884
rect 18004 16828 20076 16884
rect 20132 16828 21980 16884
rect 22036 16828 22046 16884
rect 8418 16716 8428 16772
rect 8484 16716 9772 16772
rect 9828 16716 9838 16772
rect 1586 16604 1596 16660
rect 1652 16604 2716 16660
rect 2772 16604 2782 16660
rect 3938 16604 3948 16660
rect 4004 16604 5852 16660
rect 5908 16604 5918 16660
rect 4604 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4888 16492
rect 11408 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11692 16492
rect 18212 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18496 16492
rect 25016 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25300 16492
rect 6066 16156 6076 16212
rect 6132 16156 6972 16212
rect 7028 16156 7038 16212
rect 9202 15932 9212 15988
rect 9268 15932 10780 15988
rect 10836 15932 10846 15988
rect 12002 15932 12012 15988
rect 12068 15932 13580 15988
rect 13636 15932 13646 15988
rect 19842 15932 19852 15988
rect 19908 15932 20300 15988
rect 20356 15932 20366 15988
rect 8006 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8290 15708
rect 14810 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15094 15708
rect 21614 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21898 15708
rect 28418 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28702 15708
rect 25554 15596 25564 15652
rect 25620 15596 27692 15652
rect 27748 15596 27758 15652
rect 20132 15484 22876 15540
rect 22932 15484 22942 15540
rect 20132 15316 20188 15484
rect 24546 15372 24556 15428
rect 24612 15372 25340 15428
rect 25396 15372 25406 15428
rect 8978 15260 8988 15316
rect 9044 15260 11452 15316
rect 11508 15260 11518 15316
rect 15026 15260 15036 15316
rect 15092 15260 20188 15316
rect 20514 15260 20524 15316
rect 20580 15260 26236 15316
rect 26292 15260 26302 15316
rect 22418 15148 22428 15204
rect 22484 15148 23212 15204
rect 23268 15148 25788 15204
rect 25844 15148 27356 15204
rect 27412 15148 27692 15204
rect 27748 15148 27758 15204
rect 23538 15036 23548 15092
rect 23604 15036 27244 15092
rect 27300 15036 27310 15092
rect 4604 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4888 14924
rect 11408 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11692 14924
rect 18212 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18496 14924
rect 25016 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25300 14924
rect 23650 14700 23660 14756
rect 23716 14700 26684 14756
rect 26740 14700 26750 14756
rect 8642 14588 8652 14644
rect 8708 14588 14476 14644
rect 14532 14588 14542 14644
rect 25442 14476 25452 14532
rect 25508 14476 26348 14532
rect 26404 14476 27132 14532
rect 27188 14476 28140 14532
rect 28196 14476 28206 14532
rect 3042 14364 3052 14420
rect 3108 14364 5516 14420
rect 5572 14364 5582 14420
rect 13010 14364 13020 14420
rect 13076 14364 15484 14420
rect 15540 14364 15550 14420
rect 2034 14252 2044 14308
rect 2100 14252 2716 14308
rect 2772 14252 3388 14308
rect 3444 14252 4508 14308
rect 4564 14252 4574 14308
rect 18050 14252 18060 14308
rect 18116 14252 19852 14308
rect 19908 14252 19918 14308
rect 24210 14252 24220 14308
rect 24276 14252 26684 14308
rect 26740 14252 26750 14308
rect 8006 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8290 14140
rect 14810 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15094 14140
rect 21614 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21898 14140
rect 28418 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28702 14140
rect 7970 13916 7980 13972
rect 8036 13916 9884 13972
rect 9940 13916 9950 13972
rect 4050 13692 4060 13748
rect 4116 13692 5068 13748
rect 5124 13692 5134 13748
rect 21746 13692 21756 13748
rect 21812 13692 26460 13748
rect 26516 13692 26526 13748
rect 22530 13580 22540 13636
rect 22596 13580 26236 13636
rect 26292 13580 26302 13636
rect 9874 13468 9884 13524
rect 9940 13468 11228 13524
rect 11284 13468 11294 13524
rect 24770 13468 24780 13524
rect 24836 13468 26348 13524
rect 26404 13468 26414 13524
rect 11778 13356 11788 13412
rect 11844 13356 13916 13412
rect 13972 13356 13982 13412
rect 4604 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4888 13356
rect 11408 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11692 13356
rect 18212 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18496 13356
rect 25016 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25300 13356
rect 6962 13132 6972 13188
rect 7028 13132 9100 13188
rect 9156 13132 9166 13188
rect 12450 13132 12460 13188
rect 12516 13132 13468 13188
rect 13524 13132 13534 13188
rect 14578 13020 14588 13076
rect 14644 13020 16828 13076
rect 16884 13020 21980 13076
rect 22036 13020 22046 13076
rect 4274 12908 4284 12964
rect 4340 12908 15148 12964
rect 15204 12908 15214 12964
rect 8006 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8290 12572
rect 14810 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15094 12572
rect 21614 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21898 12572
rect 28418 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28702 12572
rect 5618 12348 5628 12404
rect 5684 12348 6524 12404
rect 6580 12348 6590 12404
rect 26674 12236 26684 12292
rect 26740 12236 27356 12292
rect 27412 12236 27422 12292
rect 5282 12012 5292 12068
rect 5348 12012 5740 12068
rect 5796 12012 7756 12068
rect 7812 12012 9100 12068
rect 9156 12012 10780 12068
rect 10836 12012 10846 12068
rect 22866 11900 22876 11956
rect 22932 11900 26124 11956
rect 26180 11900 26190 11956
rect 19618 11788 19628 11844
rect 19684 11788 21308 11844
rect 21364 11788 21812 11844
rect 4604 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4888 11788
rect 11408 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11692 11788
rect 18212 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18496 11788
rect 21756 11732 21812 11788
rect 25016 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25300 11788
rect 21756 11676 23436 11732
rect 23492 11676 23502 11732
rect 20514 11452 20524 11508
rect 20580 11452 23660 11508
rect 23716 11452 23726 11508
rect 3378 11340 3388 11396
rect 3444 11340 6300 11396
rect 6356 11340 7308 11396
rect 7364 11340 8540 11396
rect 8596 11340 8606 11396
rect 1586 11228 1596 11284
rect 1652 11228 2716 11284
rect 2772 11228 2782 11284
rect 23426 11228 23436 11284
rect 23492 11228 24332 11284
rect 24388 11228 24398 11284
rect 11218 11116 11228 11172
rect 11284 11116 15820 11172
rect 15876 11116 15886 11172
rect 20738 11116 20748 11172
rect 20804 11116 22316 11172
rect 22372 11116 22382 11172
rect 24434 11116 24444 11172
rect 24500 11116 26908 11172
rect 26964 11116 26974 11172
rect 8006 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8290 11004
rect 14810 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15094 11004
rect 21614 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21898 11004
rect 28418 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28702 11004
rect 0 10836 800 10864
rect 0 10780 1820 10836
rect 1876 10780 1886 10836
rect 6178 10780 6188 10836
rect 6244 10780 8092 10836
rect 8148 10780 8158 10836
rect 0 10752 800 10780
rect 23090 10668 23100 10724
rect 23156 10668 27244 10724
rect 27300 10668 27310 10724
rect 2706 10556 2716 10612
rect 2772 10556 4284 10612
rect 4340 10556 5292 10612
rect 5348 10556 5358 10612
rect 12674 10556 12684 10612
rect 12740 10556 13468 10612
rect 13524 10556 14140 10612
rect 14196 10556 14206 10612
rect 17490 10556 17500 10612
rect 17556 10556 18284 10612
rect 18340 10556 20300 10612
rect 20356 10556 23884 10612
rect 23940 10556 24556 10612
rect 24612 10556 27356 10612
rect 27412 10556 27422 10612
rect 3266 10444 3276 10500
rect 3332 10444 3388 10500
rect 3444 10444 3454 10500
rect 8978 10444 8988 10500
rect 9044 10444 9884 10500
rect 9940 10444 9950 10500
rect 12226 10444 12236 10500
rect 12292 10444 14812 10500
rect 14868 10444 14878 10500
rect 21970 10444 21980 10500
rect 22036 10444 26236 10500
rect 26292 10444 26302 10500
rect 2370 10332 2380 10388
rect 2436 10332 4396 10388
rect 4452 10332 4462 10388
rect 4604 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4888 10220
rect 11408 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11692 10220
rect 18212 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18496 10220
rect 25016 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25300 10220
rect 26674 9884 26684 9940
rect 26740 9884 27468 9940
rect 27524 9884 27534 9940
rect 20738 9772 20748 9828
rect 20804 9772 21532 9828
rect 21588 9772 24332 9828
rect 24388 9772 24398 9828
rect 8006 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8290 9436
rect 14810 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15094 9436
rect 21614 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21898 9436
rect 28418 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28702 9436
rect 4834 9324 4844 9380
rect 4900 9324 6636 9380
rect 6692 9324 6702 9380
rect 19282 9100 19292 9156
rect 19348 9100 20188 9156
rect 20244 9100 20254 9156
rect 23538 9100 23548 9156
rect 23604 9100 27244 9156
rect 27300 9100 27310 9156
rect 10770 8988 10780 9044
rect 10836 8988 12236 9044
rect 12292 8988 12302 9044
rect 15922 8988 15932 9044
rect 15988 8988 20412 9044
rect 20468 8988 20478 9044
rect 24658 8988 24668 9044
rect 24724 8988 25340 9044
rect 25396 8988 25406 9044
rect 15362 8876 15372 8932
rect 15428 8876 19068 8932
rect 19124 8876 19134 8932
rect 29200 8820 30000 8848
rect 14130 8764 14140 8820
rect 14196 8764 16156 8820
rect 16212 8764 16222 8820
rect 24098 8764 24108 8820
rect 24164 8764 26460 8820
rect 26516 8764 26526 8820
rect 27682 8764 27692 8820
rect 27748 8764 30000 8820
rect 29200 8736 30000 8764
rect 4604 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4888 8652
rect 11408 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11692 8652
rect 18212 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18496 8652
rect 25016 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25300 8652
rect 25442 8428 25452 8484
rect 25508 8428 27132 8484
rect 27188 8428 28140 8484
rect 28196 8428 28206 8484
rect 4834 8316 4844 8372
rect 4900 8316 5852 8372
rect 5908 8316 5918 8372
rect 17938 8316 17948 8372
rect 18004 8316 19516 8372
rect 19572 8316 19582 8372
rect 14914 8204 14924 8260
rect 14980 8204 17276 8260
rect 17332 8204 18508 8260
rect 18564 8204 18574 8260
rect 29200 8148 30000 8176
rect 6402 8092 6412 8148
rect 6468 8092 7756 8148
rect 7812 8092 7822 8148
rect 19058 8092 19068 8148
rect 19124 8092 21420 8148
rect 21476 8092 22988 8148
rect 23044 8092 24332 8148
rect 24388 8092 27468 8148
rect 27524 8092 27534 8148
rect 27794 8092 27804 8148
rect 27860 8092 30000 8148
rect 29200 8064 30000 8092
rect 25778 7980 25788 8036
rect 25844 7980 27580 8036
rect 27636 7980 27646 8036
rect 12898 7868 12908 7924
rect 12964 7868 14476 7924
rect 14532 7868 14542 7924
rect 8006 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8290 7868
rect 14810 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15094 7868
rect 21614 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21898 7868
rect 28418 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28702 7868
rect 18498 7644 18508 7700
rect 18564 7644 19292 7700
rect 19348 7644 20748 7700
rect 20804 7644 20814 7700
rect 24882 7532 24892 7588
rect 24948 7532 27244 7588
rect 27300 7532 27310 7588
rect 29200 7476 30000 7504
rect 27346 7420 27356 7476
rect 27412 7420 30000 7476
rect 29200 7392 30000 7420
rect 20738 7308 20748 7364
rect 20804 7308 22652 7364
rect 22708 7308 23324 7364
rect 23380 7308 23390 7364
rect 20962 7196 20972 7252
rect 21028 7196 23100 7252
rect 23156 7196 23166 7252
rect 4604 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4888 7084
rect 11408 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11692 7084
rect 18212 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18496 7084
rect 25016 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25300 7084
rect 18610 6860 18620 6916
rect 18676 6860 21084 6916
rect 21140 6860 21150 6916
rect 23314 6860 23324 6916
rect 23380 6860 26236 6916
rect 26292 6860 26302 6916
rect 29200 6804 30000 6832
rect 11218 6748 11228 6804
rect 11284 6748 17276 6804
rect 17332 6748 17342 6804
rect 22978 6748 22988 6804
rect 23044 6748 27244 6804
rect 27300 6748 27310 6804
rect 27468 6748 30000 6804
rect 27468 6692 27524 6748
rect 29200 6720 30000 6748
rect 18050 6636 18060 6692
rect 18116 6636 20300 6692
rect 20356 6636 20366 6692
rect 25666 6636 25676 6692
rect 25732 6636 27524 6692
rect 14242 6524 14252 6580
rect 14308 6524 15484 6580
rect 15540 6524 15550 6580
rect 26114 6412 26124 6468
rect 26180 6412 26908 6468
rect 26964 6412 26974 6468
rect 8006 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8290 6300
rect 14810 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15094 6300
rect 21614 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21898 6300
rect 28418 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28702 6300
rect 0 6132 800 6160
rect 29200 6132 30000 6160
rect 0 6076 1708 6132
rect 1764 6076 1774 6132
rect 24210 6076 24220 6132
rect 24276 6076 30000 6132
rect 0 6048 800 6076
rect 29200 6048 30000 6076
rect 24658 5964 24668 6020
rect 24724 5964 26908 6020
rect 26964 5964 26974 6020
rect 19954 5740 19964 5796
rect 20020 5740 22092 5796
rect 22148 5740 22158 5796
rect 23090 5740 23100 5796
rect 23156 5740 26236 5796
rect 26292 5740 26302 5796
rect 4604 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4888 5516
rect 11408 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11692 5516
rect 18212 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18496 5516
rect 25016 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25300 5516
rect 29200 5460 30000 5488
rect 25564 5404 30000 5460
rect 24546 5292 24556 5348
rect 24612 5292 25340 5348
rect 25396 5292 25406 5348
rect 25564 5236 25620 5404
rect 29200 5376 30000 5404
rect 23202 5180 23212 5236
rect 23268 5180 25620 5236
rect 8530 5068 8540 5124
rect 8596 5068 10556 5124
rect 10612 5068 10622 5124
rect 12674 5068 12684 5124
rect 12740 5068 18060 5124
rect 18116 5068 18126 5124
rect 21532 5068 24332 5124
rect 24388 5068 24398 5124
rect 14466 4956 14476 5012
rect 14532 4956 15260 5012
rect 15316 4956 15326 5012
rect 21532 4900 21588 5068
rect 12898 4844 12908 4900
rect 12964 4844 13580 4900
rect 13636 4844 13646 4900
rect 13794 4844 13804 4900
rect 13860 4844 15148 4900
rect 15204 4844 15214 4900
rect 21522 4844 21532 4900
rect 21588 4844 21598 4900
rect 29200 4788 30000 4816
rect 28812 4732 30000 4788
rect 8006 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8290 4732
rect 14810 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15094 4732
rect 21614 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21898 4732
rect 28418 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28702 4732
rect 22194 4620 22204 4676
rect 22260 4620 26572 4676
rect 26628 4620 26638 4676
rect 28812 4564 28868 4732
rect 29200 4704 30000 4732
rect 12226 4508 12236 4564
rect 12292 4508 13692 4564
rect 13748 4508 13758 4564
rect 23090 4508 23100 4564
rect 23156 4508 24780 4564
rect 24836 4508 28868 4564
rect 13458 4396 13468 4452
rect 13524 4396 17388 4452
rect 17444 4396 17454 4452
rect 22418 4396 22428 4452
rect 22484 4396 23436 4452
rect 23492 4396 23502 4452
rect 26338 4396 26348 4452
rect 26404 4396 27468 4452
rect 27524 4396 27534 4452
rect 14914 4284 14924 4340
rect 14980 4284 15596 4340
rect 15652 4284 15662 4340
rect 9090 4172 9100 4228
rect 9156 4172 10556 4228
rect 10612 4172 10622 4228
rect 29200 4116 30000 4144
rect 21746 4060 21756 4116
rect 21812 4060 22876 4116
rect 22932 4060 22942 4116
rect 24658 4060 24668 4116
rect 24724 4060 30000 4116
rect 29200 4032 30000 4060
rect 4604 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4888 3948
rect 11408 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11692 3948
rect 18212 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18496 3948
rect 25016 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25300 3948
rect 21074 3724 21084 3780
rect 21140 3724 25004 3780
rect 25060 3724 25070 3780
rect 16146 3612 16156 3668
rect 16212 3612 17388 3668
rect 17444 3612 17454 3668
rect 22418 3612 22428 3668
rect 22484 3612 24668 3668
rect 24724 3612 24734 3668
rect 14690 3500 14700 3556
rect 14756 3500 16940 3556
rect 16996 3500 17006 3556
rect 29200 3444 30000 3472
rect 12674 3388 12684 3444
rect 12740 3388 13244 3444
rect 13300 3388 13310 3444
rect 18386 3388 18396 3444
rect 18452 3388 19068 3444
rect 19124 3388 19134 3444
rect 21522 3388 21532 3444
rect 21588 3388 24108 3444
rect 24164 3388 30000 3444
rect 29200 3360 30000 3388
rect 11106 3276 11116 3332
rect 11172 3276 11564 3332
rect 11620 3276 11630 3332
rect 8006 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8290 3164
rect 14810 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15094 3164
rect 21614 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21898 3164
rect 28418 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28702 3164
rect 29200 2772 30000 2800
rect 20850 2716 20860 2772
rect 20916 2716 30000 2772
rect 29200 2688 30000 2716
rect 29200 2100 30000 2128
rect 20178 2044 20188 2100
rect 20244 2044 30000 2100
rect 29200 2016 30000 2044
rect 29200 1428 30000 1456
rect 26674 1372 26684 1428
rect 26740 1372 30000 1428
rect 29200 1344 30000 1372
<< via3 >>
rect 8016 26628 8072 26684
rect 8120 26628 8176 26684
rect 8224 26628 8280 26684
rect 14820 26628 14876 26684
rect 14924 26628 14980 26684
rect 15028 26628 15084 26684
rect 21624 26628 21680 26684
rect 21728 26628 21784 26684
rect 21832 26628 21888 26684
rect 28428 26628 28484 26684
rect 28532 26628 28588 26684
rect 28636 26628 28692 26684
rect 4614 25844 4670 25900
rect 4718 25844 4774 25900
rect 4822 25844 4878 25900
rect 11418 25844 11474 25900
rect 11522 25844 11578 25900
rect 11626 25844 11682 25900
rect 18222 25844 18278 25900
rect 18326 25844 18382 25900
rect 18430 25844 18486 25900
rect 25026 25844 25082 25900
rect 25130 25844 25186 25900
rect 25234 25844 25290 25900
rect 24220 25228 24276 25284
rect 8016 25060 8072 25116
rect 8120 25060 8176 25116
rect 8224 25060 8280 25116
rect 14820 25060 14876 25116
rect 14924 25060 14980 25116
rect 15028 25060 15084 25116
rect 21624 25060 21680 25116
rect 21728 25060 21784 25116
rect 21832 25060 21888 25116
rect 28428 25060 28484 25116
rect 28532 25060 28588 25116
rect 28636 25060 28692 25116
rect 4614 24276 4670 24332
rect 4718 24276 4774 24332
rect 4822 24276 4878 24332
rect 11418 24276 11474 24332
rect 11522 24276 11578 24332
rect 11626 24276 11682 24332
rect 18222 24276 18278 24332
rect 18326 24276 18382 24332
rect 18430 24276 18486 24332
rect 25026 24276 25082 24332
rect 25130 24276 25186 24332
rect 25234 24276 25290 24332
rect 8016 23492 8072 23548
rect 8120 23492 8176 23548
rect 8224 23492 8280 23548
rect 14820 23492 14876 23548
rect 14924 23492 14980 23548
rect 15028 23492 15084 23548
rect 21624 23492 21680 23548
rect 21728 23492 21784 23548
rect 21832 23492 21888 23548
rect 28428 23492 28484 23548
rect 28532 23492 28588 23548
rect 28636 23492 28692 23548
rect 24220 23212 24276 23268
rect 4614 22708 4670 22764
rect 4718 22708 4774 22764
rect 4822 22708 4878 22764
rect 11418 22708 11474 22764
rect 11522 22708 11578 22764
rect 11626 22708 11682 22764
rect 18222 22708 18278 22764
rect 18326 22708 18382 22764
rect 18430 22708 18486 22764
rect 25026 22708 25082 22764
rect 25130 22708 25186 22764
rect 25234 22708 25290 22764
rect 8016 21924 8072 21980
rect 8120 21924 8176 21980
rect 8224 21924 8280 21980
rect 14820 21924 14876 21980
rect 14924 21924 14980 21980
rect 15028 21924 15084 21980
rect 21624 21924 21680 21980
rect 21728 21924 21784 21980
rect 21832 21924 21888 21980
rect 28428 21924 28484 21980
rect 28532 21924 28588 21980
rect 28636 21924 28692 21980
rect 4614 21140 4670 21196
rect 4718 21140 4774 21196
rect 4822 21140 4878 21196
rect 11418 21140 11474 21196
rect 11522 21140 11578 21196
rect 11626 21140 11682 21196
rect 18222 21140 18278 21196
rect 18326 21140 18382 21196
rect 18430 21140 18486 21196
rect 25026 21140 25082 21196
rect 25130 21140 25186 21196
rect 25234 21140 25290 21196
rect 8016 20356 8072 20412
rect 8120 20356 8176 20412
rect 8224 20356 8280 20412
rect 14820 20356 14876 20412
rect 14924 20356 14980 20412
rect 15028 20356 15084 20412
rect 21624 20356 21680 20412
rect 21728 20356 21784 20412
rect 21832 20356 21888 20412
rect 28428 20356 28484 20412
rect 28532 20356 28588 20412
rect 28636 20356 28692 20412
rect 4614 19572 4670 19628
rect 4718 19572 4774 19628
rect 4822 19572 4878 19628
rect 11418 19572 11474 19628
rect 11522 19572 11578 19628
rect 11626 19572 11682 19628
rect 18222 19572 18278 19628
rect 18326 19572 18382 19628
rect 18430 19572 18486 19628
rect 25026 19572 25082 19628
rect 25130 19572 25186 19628
rect 25234 19572 25290 19628
rect 8016 18788 8072 18844
rect 8120 18788 8176 18844
rect 8224 18788 8280 18844
rect 14820 18788 14876 18844
rect 14924 18788 14980 18844
rect 15028 18788 15084 18844
rect 21624 18788 21680 18844
rect 21728 18788 21784 18844
rect 21832 18788 21888 18844
rect 28428 18788 28484 18844
rect 28532 18788 28588 18844
rect 28636 18788 28692 18844
rect 4614 18004 4670 18060
rect 4718 18004 4774 18060
rect 4822 18004 4878 18060
rect 11418 18004 11474 18060
rect 11522 18004 11578 18060
rect 11626 18004 11682 18060
rect 18222 18004 18278 18060
rect 18326 18004 18382 18060
rect 18430 18004 18486 18060
rect 25026 18004 25082 18060
rect 25130 18004 25186 18060
rect 25234 18004 25290 18060
rect 8016 17220 8072 17276
rect 8120 17220 8176 17276
rect 8224 17220 8280 17276
rect 14820 17220 14876 17276
rect 14924 17220 14980 17276
rect 15028 17220 15084 17276
rect 21624 17220 21680 17276
rect 21728 17220 21784 17276
rect 21832 17220 21888 17276
rect 28428 17220 28484 17276
rect 28532 17220 28588 17276
rect 28636 17220 28692 17276
rect 4614 16436 4670 16492
rect 4718 16436 4774 16492
rect 4822 16436 4878 16492
rect 11418 16436 11474 16492
rect 11522 16436 11578 16492
rect 11626 16436 11682 16492
rect 18222 16436 18278 16492
rect 18326 16436 18382 16492
rect 18430 16436 18486 16492
rect 25026 16436 25082 16492
rect 25130 16436 25186 16492
rect 25234 16436 25290 16492
rect 8016 15652 8072 15708
rect 8120 15652 8176 15708
rect 8224 15652 8280 15708
rect 14820 15652 14876 15708
rect 14924 15652 14980 15708
rect 15028 15652 15084 15708
rect 21624 15652 21680 15708
rect 21728 15652 21784 15708
rect 21832 15652 21888 15708
rect 28428 15652 28484 15708
rect 28532 15652 28588 15708
rect 28636 15652 28692 15708
rect 4614 14868 4670 14924
rect 4718 14868 4774 14924
rect 4822 14868 4878 14924
rect 11418 14868 11474 14924
rect 11522 14868 11578 14924
rect 11626 14868 11682 14924
rect 18222 14868 18278 14924
rect 18326 14868 18382 14924
rect 18430 14868 18486 14924
rect 25026 14868 25082 14924
rect 25130 14868 25186 14924
rect 25234 14868 25290 14924
rect 8016 14084 8072 14140
rect 8120 14084 8176 14140
rect 8224 14084 8280 14140
rect 14820 14084 14876 14140
rect 14924 14084 14980 14140
rect 15028 14084 15084 14140
rect 21624 14084 21680 14140
rect 21728 14084 21784 14140
rect 21832 14084 21888 14140
rect 28428 14084 28484 14140
rect 28532 14084 28588 14140
rect 28636 14084 28692 14140
rect 4614 13300 4670 13356
rect 4718 13300 4774 13356
rect 4822 13300 4878 13356
rect 11418 13300 11474 13356
rect 11522 13300 11578 13356
rect 11626 13300 11682 13356
rect 18222 13300 18278 13356
rect 18326 13300 18382 13356
rect 18430 13300 18486 13356
rect 25026 13300 25082 13356
rect 25130 13300 25186 13356
rect 25234 13300 25290 13356
rect 8016 12516 8072 12572
rect 8120 12516 8176 12572
rect 8224 12516 8280 12572
rect 14820 12516 14876 12572
rect 14924 12516 14980 12572
rect 15028 12516 15084 12572
rect 21624 12516 21680 12572
rect 21728 12516 21784 12572
rect 21832 12516 21888 12572
rect 28428 12516 28484 12572
rect 28532 12516 28588 12572
rect 28636 12516 28692 12572
rect 4614 11732 4670 11788
rect 4718 11732 4774 11788
rect 4822 11732 4878 11788
rect 11418 11732 11474 11788
rect 11522 11732 11578 11788
rect 11626 11732 11682 11788
rect 18222 11732 18278 11788
rect 18326 11732 18382 11788
rect 18430 11732 18486 11788
rect 25026 11732 25082 11788
rect 25130 11732 25186 11788
rect 25234 11732 25290 11788
rect 8016 10948 8072 11004
rect 8120 10948 8176 11004
rect 8224 10948 8280 11004
rect 14820 10948 14876 11004
rect 14924 10948 14980 11004
rect 15028 10948 15084 11004
rect 21624 10948 21680 11004
rect 21728 10948 21784 11004
rect 21832 10948 21888 11004
rect 28428 10948 28484 11004
rect 28532 10948 28588 11004
rect 28636 10948 28692 11004
rect 4614 10164 4670 10220
rect 4718 10164 4774 10220
rect 4822 10164 4878 10220
rect 11418 10164 11474 10220
rect 11522 10164 11578 10220
rect 11626 10164 11682 10220
rect 18222 10164 18278 10220
rect 18326 10164 18382 10220
rect 18430 10164 18486 10220
rect 25026 10164 25082 10220
rect 25130 10164 25186 10220
rect 25234 10164 25290 10220
rect 8016 9380 8072 9436
rect 8120 9380 8176 9436
rect 8224 9380 8280 9436
rect 14820 9380 14876 9436
rect 14924 9380 14980 9436
rect 15028 9380 15084 9436
rect 21624 9380 21680 9436
rect 21728 9380 21784 9436
rect 21832 9380 21888 9436
rect 28428 9380 28484 9436
rect 28532 9380 28588 9436
rect 28636 9380 28692 9436
rect 4614 8596 4670 8652
rect 4718 8596 4774 8652
rect 4822 8596 4878 8652
rect 11418 8596 11474 8652
rect 11522 8596 11578 8652
rect 11626 8596 11682 8652
rect 18222 8596 18278 8652
rect 18326 8596 18382 8652
rect 18430 8596 18486 8652
rect 25026 8596 25082 8652
rect 25130 8596 25186 8652
rect 25234 8596 25290 8652
rect 8016 7812 8072 7868
rect 8120 7812 8176 7868
rect 8224 7812 8280 7868
rect 14820 7812 14876 7868
rect 14924 7812 14980 7868
rect 15028 7812 15084 7868
rect 21624 7812 21680 7868
rect 21728 7812 21784 7868
rect 21832 7812 21888 7868
rect 28428 7812 28484 7868
rect 28532 7812 28588 7868
rect 28636 7812 28692 7868
rect 4614 7028 4670 7084
rect 4718 7028 4774 7084
rect 4822 7028 4878 7084
rect 11418 7028 11474 7084
rect 11522 7028 11578 7084
rect 11626 7028 11682 7084
rect 18222 7028 18278 7084
rect 18326 7028 18382 7084
rect 18430 7028 18486 7084
rect 25026 7028 25082 7084
rect 25130 7028 25186 7084
rect 25234 7028 25290 7084
rect 8016 6244 8072 6300
rect 8120 6244 8176 6300
rect 8224 6244 8280 6300
rect 14820 6244 14876 6300
rect 14924 6244 14980 6300
rect 15028 6244 15084 6300
rect 21624 6244 21680 6300
rect 21728 6244 21784 6300
rect 21832 6244 21888 6300
rect 28428 6244 28484 6300
rect 28532 6244 28588 6300
rect 28636 6244 28692 6300
rect 4614 5460 4670 5516
rect 4718 5460 4774 5516
rect 4822 5460 4878 5516
rect 11418 5460 11474 5516
rect 11522 5460 11578 5516
rect 11626 5460 11682 5516
rect 18222 5460 18278 5516
rect 18326 5460 18382 5516
rect 18430 5460 18486 5516
rect 25026 5460 25082 5516
rect 25130 5460 25186 5516
rect 25234 5460 25290 5516
rect 8016 4676 8072 4732
rect 8120 4676 8176 4732
rect 8224 4676 8280 4732
rect 14820 4676 14876 4732
rect 14924 4676 14980 4732
rect 15028 4676 15084 4732
rect 21624 4676 21680 4732
rect 21728 4676 21784 4732
rect 21832 4676 21888 4732
rect 28428 4676 28484 4732
rect 28532 4676 28588 4732
rect 28636 4676 28692 4732
rect 4614 3892 4670 3948
rect 4718 3892 4774 3948
rect 4822 3892 4878 3948
rect 11418 3892 11474 3948
rect 11522 3892 11578 3948
rect 11626 3892 11682 3948
rect 18222 3892 18278 3948
rect 18326 3892 18382 3948
rect 18430 3892 18486 3948
rect 25026 3892 25082 3948
rect 25130 3892 25186 3948
rect 25234 3892 25290 3948
rect 8016 3108 8072 3164
rect 8120 3108 8176 3164
rect 8224 3108 8280 3164
rect 14820 3108 14876 3164
rect 14924 3108 14980 3164
rect 15028 3108 15084 3164
rect 21624 3108 21680 3164
rect 21728 3108 21784 3164
rect 21832 3108 21888 3164
rect 28428 3108 28484 3164
rect 28532 3108 28588 3164
rect 28636 3108 28692 3164
<< metal4 >>
rect 4586 25900 4906 26716
rect 4586 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4906 25900
rect 4586 24332 4906 25844
rect 4586 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4906 24332
rect 4586 22764 4906 24276
rect 4586 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4906 22764
rect 4586 21196 4906 22708
rect 4586 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4906 21196
rect 4586 19628 4906 21140
rect 4586 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4906 19628
rect 4586 18060 4906 19572
rect 4586 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4906 18060
rect 4586 16492 4906 18004
rect 4586 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4906 16492
rect 4586 14924 4906 16436
rect 4586 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4906 14924
rect 4586 13356 4906 14868
rect 4586 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4906 13356
rect 4586 11788 4906 13300
rect 4586 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4906 11788
rect 4586 10220 4906 11732
rect 4586 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4906 10220
rect 4586 8652 4906 10164
rect 4586 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4906 8652
rect 4586 7084 4906 8596
rect 4586 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4906 7084
rect 4586 5516 4906 7028
rect 4586 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4906 5516
rect 4586 3948 4906 5460
rect 4586 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4906 3948
rect 4586 3076 4906 3892
rect 7988 26684 8308 26716
rect 7988 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8308 26684
rect 7988 25116 8308 26628
rect 7988 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8308 25116
rect 7988 23548 8308 25060
rect 7988 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8308 23548
rect 7988 21980 8308 23492
rect 7988 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8308 21980
rect 7988 20412 8308 21924
rect 7988 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8308 20412
rect 7988 18844 8308 20356
rect 7988 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8308 18844
rect 7988 17276 8308 18788
rect 7988 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8308 17276
rect 7988 15708 8308 17220
rect 7988 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8308 15708
rect 7988 14140 8308 15652
rect 7988 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8308 14140
rect 7988 12572 8308 14084
rect 7988 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8308 12572
rect 7988 11004 8308 12516
rect 7988 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8308 11004
rect 7988 9436 8308 10948
rect 7988 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8308 9436
rect 7988 7868 8308 9380
rect 7988 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8308 7868
rect 7988 6300 8308 7812
rect 7988 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8308 6300
rect 7988 4732 8308 6244
rect 7988 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8308 4732
rect 7988 3164 8308 4676
rect 7988 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8308 3164
rect 7988 3076 8308 3108
rect 11390 25900 11710 26716
rect 11390 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11710 25900
rect 11390 24332 11710 25844
rect 11390 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11710 24332
rect 11390 22764 11710 24276
rect 11390 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11710 22764
rect 11390 21196 11710 22708
rect 11390 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11710 21196
rect 11390 19628 11710 21140
rect 11390 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11710 19628
rect 11390 18060 11710 19572
rect 11390 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11710 18060
rect 11390 16492 11710 18004
rect 11390 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11710 16492
rect 11390 14924 11710 16436
rect 11390 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11710 14924
rect 11390 13356 11710 14868
rect 11390 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11710 13356
rect 11390 11788 11710 13300
rect 11390 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11710 11788
rect 11390 10220 11710 11732
rect 11390 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11710 10220
rect 11390 8652 11710 10164
rect 11390 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11710 8652
rect 11390 7084 11710 8596
rect 11390 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11710 7084
rect 11390 5516 11710 7028
rect 11390 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11710 5516
rect 11390 3948 11710 5460
rect 11390 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11710 3948
rect 11390 3076 11710 3892
rect 14792 26684 15112 26716
rect 14792 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15112 26684
rect 14792 25116 15112 26628
rect 14792 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15112 25116
rect 14792 23548 15112 25060
rect 14792 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15112 23548
rect 14792 21980 15112 23492
rect 14792 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15112 21980
rect 14792 20412 15112 21924
rect 14792 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15112 20412
rect 14792 18844 15112 20356
rect 14792 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15112 18844
rect 14792 17276 15112 18788
rect 14792 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15112 17276
rect 14792 15708 15112 17220
rect 14792 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15112 15708
rect 14792 14140 15112 15652
rect 14792 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15112 14140
rect 14792 12572 15112 14084
rect 14792 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15112 12572
rect 14792 11004 15112 12516
rect 14792 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15112 11004
rect 14792 9436 15112 10948
rect 14792 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15112 9436
rect 14792 7868 15112 9380
rect 14792 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15112 7868
rect 14792 6300 15112 7812
rect 14792 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15112 6300
rect 14792 4732 15112 6244
rect 14792 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15112 4732
rect 14792 3164 15112 4676
rect 14792 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15112 3164
rect 14792 3076 15112 3108
rect 18194 25900 18514 26716
rect 18194 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18514 25900
rect 18194 24332 18514 25844
rect 18194 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18514 24332
rect 18194 22764 18514 24276
rect 18194 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18514 22764
rect 18194 21196 18514 22708
rect 18194 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18514 21196
rect 18194 19628 18514 21140
rect 18194 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18514 19628
rect 18194 18060 18514 19572
rect 18194 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18514 18060
rect 18194 16492 18514 18004
rect 18194 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18514 16492
rect 18194 14924 18514 16436
rect 18194 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18514 14924
rect 18194 13356 18514 14868
rect 18194 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18514 13356
rect 18194 11788 18514 13300
rect 18194 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18514 11788
rect 18194 10220 18514 11732
rect 18194 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18514 10220
rect 18194 8652 18514 10164
rect 18194 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18514 8652
rect 18194 7084 18514 8596
rect 18194 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18514 7084
rect 18194 5516 18514 7028
rect 18194 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18514 5516
rect 18194 3948 18514 5460
rect 18194 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18514 3948
rect 18194 3076 18514 3892
rect 21596 26684 21916 26716
rect 21596 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21916 26684
rect 21596 25116 21916 26628
rect 24998 25900 25318 26716
rect 24998 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25318 25900
rect 21596 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21916 25116
rect 21596 23548 21916 25060
rect 21596 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21916 23548
rect 21596 21980 21916 23492
rect 24220 25284 24276 25294
rect 24220 23268 24276 25228
rect 24220 23202 24276 23212
rect 24998 24332 25318 25844
rect 24998 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25318 24332
rect 21596 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21916 21980
rect 21596 20412 21916 21924
rect 21596 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21916 20412
rect 21596 18844 21916 20356
rect 21596 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21916 18844
rect 21596 17276 21916 18788
rect 21596 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21916 17276
rect 21596 15708 21916 17220
rect 21596 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21916 15708
rect 21596 14140 21916 15652
rect 21596 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21916 14140
rect 21596 12572 21916 14084
rect 21596 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21916 12572
rect 21596 11004 21916 12516
rect 21596 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21916 11004
rect 21596 9436 21916 10948
rect 21596 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21916 9436
rect 21596 7868 21916 9380
rect 21596 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21916 7868
rect 21596 6300 21916 7812
rect 21596 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21916 6300
rect 21596 4732 21916 6244
rect 21596 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21916 4732
rect 21596 3164 21916 4676
rect 21596 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21916 3164
rect 21596 3076 21916 3108
rect 24998 22764 25318 24276
rect 24998 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25318 22764
rect 24998 21196 25318 22708
rect 24998 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25318 21196
rect 24998 19628 25318 21140
rect 24998 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25318 19628
rect 24998 18060 25318 19572
rect 24998 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25318 18060
rect 24998 16492 25318 18004
rect 24998 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25318 16492
rect 24998 14924 25318 16436
rect 24998 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25318 14924
rect 24998 13356 25318 14868
rect 24998 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25318 13356
rect 24998 11788 25318 13300
rect 24998 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25318 11788
rect 24998 10220 25318 11732
rect 24998 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25318 10220
rect 24998 8652 25318 10164
rect 24998 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25318 8652
rect 24998 7084 25318 8596
rect 24998 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25318 7084
rect 24998 5516 25318 7028
rect 24998 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25318 5516
rect 24998 3948 25318 5460
rect 24998 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25318 3948
rect 24998 3076 25318 3892
rect 28400 26684 28720 26716
rect 28400 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28720 26684
rect 28400 25116 28720 26628
rect 28400 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28720 25116
rect 28400 23548 28720 25060
rect 28400 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28720 23548
rect 28400 21980 28720 23492
rect 28400 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28720 21980
rect 28400 20412 28720 21924
rect 28400 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28720 20412
rect 28400 18844 28720 20356
rect 28400 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28720 18844
rect 28400 17276 28720 18788
rect 28400 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28720 17276
rect 28400 15708 28720 17220
rect 28400 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28720 15708
rect 28400 14140 28720 15652
rect 28400 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28720 14140
rect 28400 12572 28720 14084
rect 28400 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28720 12572
rect 28400 11004 28720 12516
rect 28400 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28720 11004
rect 28400 9436 28720 10948
rect 28400 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28720 9436
rect 28400 7868 28720 9380
rect 28400 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28720 7868
rect 28400 6300 28720 7812
rect 28400 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28720 6300
rect 28400 4732 28720 6244
rect 28400 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28720 4732
rect 28400 3164 28720 4676
rect 28400 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28720 3164
rect 28400 3076 28720 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _047_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _048_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13664 0 -1 10976
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _049_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _050_
timestamp 1698431365
transform -1 0 8848 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _051_
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _052_
timestamp 1698431365
transform -1 0 6384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _053_
timestamp 1698431365
transform -1 0 5264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _054_
timestamp 1698431365
transform 1 0 3136 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _055_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _056_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _057_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _058_
timestamp 1698431365
transform -1 0 4704 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _059_
timestamp 1698431365
transform -1 0 15568 0 -1 14112
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _060_
timestamp 1698431365
transform -1 0 14224 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _061_
timestamp 1698431365
transform -1 0 11984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _062_
timestamp 1698431365
transform 1 0 15680 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _063_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _064_
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _065_
timestamp 1698431365
transform 1 0 9520 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _066_
timestamp 1698431365
transform -1 0 10304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _067_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _068_
timestamp 1698431365
transform -1 0 16128 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _069_
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _070_
timestamp 1698431365
transform 1 0 14336 0 1 10976
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _071_
timestamp 1698431365
transform -1 0 26880 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _072_
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _073_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _074_
timestamp 1698431365
transform -1 0 22064 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _075_
timestamp 1698431365
transform -1 0 27440 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _076_
timestamp 1698431365
transform -1 0 26544 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _077_
timestamp 1698431365
transform -1 0 24752 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _078_
timestamp 1698431365
transform -1 0 22848 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _079_
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _080_
timestamp 1698431365
transform -1 0 20832 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _081_
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _082_
timestamp 1698431365
transform -1 0 23520 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _083_
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _084_
timestamp 1698431365
transform -1 0 27664 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _085_
timestamp 1698431365
transform 1 0 20048 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _086_
timestamp 1698431365
transform -1 0 24080 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _087_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _088_
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _089_
timestamp 1698431365
transform 1 0 21280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _090_
timestamp 1698431365
transform 1 0 18592 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _091_
timestamp 1698431365
transform -1 0 18816 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16016 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _093_
timestamp 1698431365
transform -1 0 14336 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _095_
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _096_
timestamp 1698431365
transform 1 0 4032 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _097_
timestamp 1698431365
transform 1 0 2688 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _098_
timestamp 1698431365
transform -1 0 5376 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _099_
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _100_
timestamp 1698431365
transform 1 0 3360 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _101_
timestamp 1698431365
transform -1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _102_
timestamp 1698431365
transform -1 0 5824 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _103_
timestamp 1698431365
transform -1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _104_
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _105_
timestamp 1698431365
transform -1 0 12880 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _106_
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _107_
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _108_
timestamp 1698431365
transform 1 0 9296 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _109_
timestamp 1698431365
transform 1 0 7504 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _110_
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _111_
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _112_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _113_
timestamp 1698431365
transform -1 0 15792 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _114_
timestamp 1698431365
transform -1 0 27104 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _115_
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _116_
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _117_
timestamp 1698431365
transform 1 0 17360 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _118_
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _119_
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _120_
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _121_
timestamp 1698431365
transform 1 0 19824 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _122_
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _123_
timestamp 1698431365
transform 1 0 16128 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _124_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _125_
timestamp 1698431365
transform 1 0 22624 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _126_
timestamp 1698431365
transform 1 0 21280 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _127_
timestamp 1698431365
transform 1 0 19376 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _128_
timestamp 1698431365
transform -1 0 23520 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _129_
timestamp 1698431365
transform -1 0 27328 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _130_
timestamp 1698431365
transform 1 0 22400 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _131_
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _132_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _133_
timestamp 1698431365
transform 1 0 14672 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _134_
timestamp 1698431365
transform 1 0 12208 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _135_
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _144_
timestamp 1698431365
transform 1 0 21280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _145_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1698431365
transform -1 0 10864 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _147_
timestamp 1698431365
transform 1 0 11088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _148_
timestamp 1698431365
transform 1 0 24416 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1698431365
transform 1 0 21952 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _150_
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1698431365
transform 1 0 9744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _152_
timestamp 1698431365
transform 1 0 25760 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _153_
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_
timestamp 1698431365
transform 1 0 11760 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _156_
timestamp 1698431365
transform 1 0 25424 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _157_
timestamp 1698431365
transform -1 0 11424 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _159_
timestamp 1698431365
transform 1 0 23744 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _160_
timestamp 1698431365
transform 1 0 21728 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _161_
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _162_
timestamp 1698431365
transform 1 0 14336 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _163_
timestamp 1698431365
transform -1 0 12208 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _164_
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _165_
timestamp 1698431365
transform -1 0 4032 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _166_
timestamp 1698431365
transform 1 0 25088 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _167_
timestamp 1698431365
transform 1 0 14784 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _168_
timestamp 1698431365
transform -1 0 9520 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _169_
timestamp 1698431365
transform 1 0 10864 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _170_
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _171_
timestamp 1698431365
transform 1 0 26096 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _172_
timestamp 1698431365
transform -1 0 11088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_
timestamp 1698431365
transform 1 0 16352 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _174_
timestamp 1698431365
transform 1 0 25760 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _175_
timestamp 1698431365
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _176_
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _177_
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _178_
timestamp 1698431365
transform 1 0 12432 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1698431365
transform 1 0 15456 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _180_
timestamp 1698431365
transform 1 0 10080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1698431365
transform -1 0 10080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__049__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I
timestamp 1698431365
transform 1 0 8960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1698431365
transform 1 0 6608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1698431365
transform -1 0 5936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1698431365
transform 1 0 2912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1698431365
transform 1 0 6608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1698431365
transform -1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1698431365
transform -1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1698431365
transform -1 0 21616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__I
timestamp 1698431365
transform 1 0 25424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I
timestamp 1698431365
transform 1 0 23072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__CLK
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__CLK
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__CLK
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__CLK
timestamp 1698431365
transform -1 0 24080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__CLK
timestamp 1698431365
transform 1 0 21840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__CLK
timestamp 1698431365
transform -1 0 26096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__CLK
timestamp 1698431365
transform -1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__CLK
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__CLK
timestamp 1698431365
transform 1 0 21952 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__CLK
timestamp 1698431365
transform 1 0 28112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__CLK
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__CLK
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__CLK
timestamp 1698431365
transform 1 0 28112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__CLK
timestamp 1698431365
transform 1 0 23296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__CLK
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__CLK
timestamp 1698431365
transform 1 0 18480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform 1 0 15232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 11312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 8848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 3360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 15568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 23744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 7504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 6160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 14896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 17920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 20832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 14224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 26320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 19600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 27664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 11760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 4704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 24640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 18368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 22848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 4256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__84 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__85
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__86
timestamp 1698431365
transform -1 0 26432 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__87
timestamp 1698431365
transform 1 0 26320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__88
timestamp 1698431365
transform -1 0 2688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__89
timestamp 1698431365
transform -1 0 20384 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cbx_1__0__90
timestamp 1698431365
transform -1 0 2016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_44 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_54 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_118
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_132
timestamp 1698431365
transform 1 0 16128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_148
timestamp 1698431365
transform 1 0 17920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_154
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_166
timestamp 1698431365
transform 1 0 19936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_200
timestamp 1698431365
transform 1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_220
timestamp 1698431365
transform 1 0 25984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_234
timestamp 1698431365
transform 1 0 27552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_34 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_50
timestamp 1698431365
transform 1 0 6944 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_62
timestamp 1698431365
transform 1 0 8288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_85
timestamp 1698431365
transform 1 0 10864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_91
timestamp 1698431365
transform 1 0 11536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_105
timestamp 1698431365
transform 1 0 13104 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_119
timestamp 1698431365
transform 1 0 14672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_129
timestamp 1698431365
transform 1 0 15792 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_137
timestamp 1698431365
transform 1 0 16688 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_160
timestamp 1698431365
transform 1 0 19264 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_164
timestamp 1698431365
transform 1 0 19712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_222
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_239
timestamp 1698431365
transform 1 0 28112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_69
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_73
timestamp 1698431365
transform 1 0 9520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_113
timestamp 1698431365
transform 1 0 14000 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_122
timestamp 1698431365
transform 1 0 15008 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_138
timestamp 1698431365
transform 1 0 16800 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_148
timestamp 1698431365
transform 1 0 17920 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_237
timestamp 1698431365
transform 1 0 27888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_158
timestamp 1698431365
transform 1 0 19040 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_175
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_183
timestamp 1698431365
transform 1 0 21840 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_200
timestamp 1698431365
transform 1 0 23744 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_237
timestamp 1698431365
transform 1 0 27888 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_6
timestamp 1698431365
transform 1 0 2016 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_22
timestamp 1698431365
transform 1 0 3808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_30
timestamp 1698431365
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_132
timestamp 1698431365
transform 1 0 16128 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_140
timestamp 1698431365
transform 1 0 17024 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_157
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_173
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_224
timestamp 1698431365
transform 1 0 26432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_237
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_38
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_116
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_152
timestamp 1698431365
transform 1 0 18368 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_155
timestamp 1698431365
transform 1 0 18704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_159
timestamp 1698431365
transform 1 0 19152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_194
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_198
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_237
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_18
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_63
timestamp 1698431365
transform 1 0 8400 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_95
timestamp 1698431365
transform 1 0 11984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_115
timestamp 1698431365
transform 1 0 14224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_153
timestamp 1698431365
transform 1 0 18480 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_162
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_170
timestamp 1698431365
transform 1 0 20384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_186
timestamp 1698431365
transform 1 0 22176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_10
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_46
timestamp 1698431365
transform 1 0 6496 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_62
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_88
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_96
timestamp 1698431365
transform 1 0 12096 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_216
timestamp 1698431365
transform 1 0 25536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_237
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_49
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_66
timestamp 1698431365
transform 1 0 8736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_70
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_78
timestamp 1698431365
transform 1 0 10080 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_148
timestamp 1698431365
transform 1 0 17920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_156
timestamp 1698431365
transform 1 0 18816 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_212
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_216
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_220
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_6
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_110
timestamp 1698431365
transform 1 0 13664 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_118
timestamp 1698431365
transform 1 0 14560 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_135
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_156
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_160
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_203
timestamp 1698431365
transform 1 0 24080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_237
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_51
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_89
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_109
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_154
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_162
timestamp 1698431365
transform 1 0 19488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_166
timestamp 1698431365
transform 1 0 19936 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_235
timestamp 1698431365
transform 1 0 27664 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_126
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_134
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_198
timestamp 1698431365
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_237
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_43
timestamp 1698431365
transform 1 0 6160 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_60
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_68
timestamp 1698431365
transform 1 0 8960 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_103
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_167
timestamp 1698431365
transform 1 0 20048 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_239
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_44
timestamp 1698431365
transform 1 0 6272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_61
timestamp 1698431365
transform 1 0 8176 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_74
timestamp 1698431365
transform 1 0 9632 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_83
timestamp 1698431365
transform 1 0 10640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_87
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_127
timestamp 1698431365
transform 1 0 15568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_135
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_167
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_175
timestamp 1698431365
transform 1 0 20944 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_214
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_217
timestamp 1698431365
transform 1 0 25648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_237
timestamp 1698431365
transform 1 0 27888 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_132
timestamp 1698431365
transform 1 0 16128 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_164
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_52
timestamp 1698431365
transform 1 0 7168 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_60
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_162
timestamp 1698431365
transform 1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_164
timestamp 1698431365
transform 1 0 19712 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_237
timestamp 1698431365
transform 1 0 27888 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_65
timestamp 1698431365
transform 1 0 8624 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_73
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_90
timestamp 1698431365
transform 1 0 11424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_98
timestamp 1698431365
transform 1 0 12320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_155
timestamp 1698431365
transform 1 0 18704 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_235
timestamp 1698431365
transform 1 0 27664 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_239
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_182
timestamp 1698431365
transform 1 0 21728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_186
timestamp 1698431365
transform 1 0 22176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_190
timestamp 1698431365
transform 1 0 22624 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_224
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_49
timestamp 1698431365
transform 1 0 6832 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_121
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_192
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_234
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_81
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_89
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_240
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_149
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_157
timestamp 1698431365
transform 1 0 18928 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_228
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_126
timestamp 1698431365
transform 1 0 15456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_177
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_181
timestamp 1698431365
transform 1 0 21616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_185
timestamp 1698431365
transform 1 0 22064 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_224
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_131
timestamp 1698431365
transform 1 0 16016 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_148
timestamp 1698431365
transform 1 0 17920 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_164
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_203
timestamp 1698431365
transform 1 0 24080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_221
timestamp 1698431365
transform 1 0 26096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_108
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_126
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_134
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_209
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_213
timestamp 1698431365
transform 1 0 25200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_90
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_122
timestamp 1698431365
transform 1 0 15008 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_166
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_176
timestamp 1698431365
transform 1 0 21056 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_200
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_224
timestamp 1698431365
transform 1 0 26432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_237
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_97
timestamp 1698431365
transform 1 0 12208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_117
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_119
timestamp 1698431365
transform 1 0 14672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_132
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_140
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_156
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_160
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_162
timestamp 1698431365
transform 1 0 19488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_191
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_197
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_224
timestamp 1698431365
transform 1 0 26432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_226
timestamp 1698431365
transform 1 0 26656 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_237
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_24
timestamp 1698431365
transform 1 0 4032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_40
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_43
timestamp 1698431365
transform 1 0 6160 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_51
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_55
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_63
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_83
timestamp 1698431365
transform 1 0 10640 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_99
timestamp 1698431365
transform 1 0 12432 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_107
timestamp 1698431365
transform 1 0 13328 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_111
timestamp 1698431365
transform 1 0 13776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_121
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698431365
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_16
timestamp 1698431365
transform 1 0 3136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_117
timestamp 1698431365
transform 1 0 14448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_127
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_135
timestamp 1698431365
transform 1 0 16464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_145
timestamp 1698431365
transform 1 0 17584 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_149
timestamp 1698431365
transform 1 0 18032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_183
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_223
timestamp 1698431365
transform 1 0 26320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_237
timestamp 1698431365
transform 1 0 27888 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_6
timestamp 1698431365
transform 1 0 2016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_21
timestamp 1698431365
transform 1 0 3696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_51
timestamp 1698431365
transform 1 0 7056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_53
timestamp 1698431365
transform 1 0 7280 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_70
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_108
timestamp 1698431365
transform 1 0 13440 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_119
timestamp 1698431365
transform 1 0 14672 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_123
timestamp 1698431365
transform 1 0 15120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_135
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_148
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_162
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_182
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_200
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_240
timestamp 1698431365
transform 1 0 28224 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20720 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 16464 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 27888 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 20832 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 20048 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 17920 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 20944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 15456 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform 1 0 18256 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 11424 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 26096 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform 1 0 6272 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 27888 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 27888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 23968 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 28336 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform 1 0 6384 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 27888 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 8624 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 23744 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform -1 0 27888 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 13216 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform -1 0 16128 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 8400 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 16128 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 28112 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 9296 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 5264 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform 1 0 26096 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 18928 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 24528 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 11424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 28336 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 25200 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 8848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 3472 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 16240 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 22848 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 24528 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 7504 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 14896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 18592 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 27664 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 14896 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 17584 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 15792 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 26992 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 10864 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 20496 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 23296 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 28336 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 3808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 17920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 22624 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 19264 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform -1 0 28336 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform -1 0 28336 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 4144 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input42 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform -1 0 10752 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform 1 0 20608 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform 1 0 23296 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output49
timestamp 1698431365
transform 1 0 25200 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output50
timestamp 1698431365
transform 1 0 11984 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output51 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698431365
transform 1 0 15008 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform 1 0 22624 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform 1 0 18816 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output55
timestamp 1698431365
transform 1 0 26768 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output56
timestamp 1698431365
transform 1 0 26432 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output57
timestamp 1698431365
transform 1 0 26768 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform -1 0 11536 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output60
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output62
timestamp 1698431365
transform 1 0 13552 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output63
timestamp 1698431365
transform 1 0 9520 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output64
timestamp 1698431365
transform 1 0 11536 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform -1 0 26768 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform 1 0 22176 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output68
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output69
timestamp 1698431365
transform -1 0 8960 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output70
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output71
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output72
timestamp 1698431365
transform -1 0 3136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output73
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output74
timestamp 1698431365
transform -1 0 7056 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output75
timestamp 1698431365
transform -1 0 3696 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output76
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output77
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output78
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output79
timestamp 1698431365
transform 1 0 26768 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output80
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output81
timestamp 1698431365
transform 1 0 13552 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output82
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output83
timestamp 1698431365
transform 1 0 18368 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_30 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 28560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_31
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_32
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_33
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_34
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_35
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_36
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_37
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_38
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_39
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_40
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_41
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 28560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_42
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_43
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_44
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_45
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_46
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_47
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_48
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_49
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_50
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 28560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 28560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_61
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_62
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_63
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_64
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_65
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_66
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_67
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_68
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_69
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_70
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_71
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_72
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_73
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_74
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_75
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_76
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_77
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_78
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_81
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_86
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_87
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_88
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_89
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_90
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_91
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_92
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_93
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_94
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_95
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_96
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_97
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_98
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_99
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_100
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_101
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_102
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_103
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_104
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_105
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_106
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_107
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_108
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_109
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_110
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_111
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_112
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_113
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_114
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_115
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_116
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_117
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_118
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_119
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_120
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_121
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_122
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_123
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_124
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_125
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_126
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_127
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_128
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_129
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_130
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_131
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_132
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_133
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_134
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_135
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_136
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_137
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_138
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_139
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_140
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_141
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_142
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_143
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_144
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_145
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_146
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_147
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_148
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_149
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_150
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_151
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_152
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_153
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_154
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_155
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_156
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_157
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 310 870
<< labels >>
flabel metal3 s 29200 1344 30000 1456 0 FreeSans 448 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
port 0 nsew signal tristate
flabel metal2 s 24864 29200 24976 30000 0 FreeSans 448 90 0 0 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
port 1 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
port 2 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
port 3 nsew signal tristate
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 29200 8736 30000 8848 0 FreeSans 448 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 1344 29200 1456 30000 0 FreeSans 448 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 29200 20832 30000 20944 0 FreeSans 448 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal2 s 24192 29200 24304 30000 0 FreeSans 448 90 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 8736 29200 8848 30000 0 FreeSans 448 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 3360 29200 3472 30000 0 FreeSans 448 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal2 s 15456 29200 15568 30000 0 FreeSans 448 90 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 29200 29568 30000 29680 0 FreeSans 448 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 23520 29200 23632 30000 0 FreeSans 448 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 7392 29200 7504 30000 0 FreeSans 448 90 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal2 s 6048 29200 6160 30000 0 FreeSans 448 90 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal2 s 4704 29200 4816 30000 0 FreeSans 448 90 0 0 chanx_left_in[2]
port 18 nsew signal input
flabel metal2 s 14784 29200 14896 30000 0 FreeSans 448 90 0 0 chanx_left_in[3]
port 19 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chanx_left_in[4]
port 20 nsew signal input
flabel metal3 s 29200 21504 30000 21616 0 FreeSans 448 0 0 0 chanx_left_in[5]
port 21 nsew signal input
flabel metal3 s 29200 2016 30000 2128 0 FreeSans 448 0 0 0 chanx_left_in[6]
port 22 nsew signal input
flabel metal2 s 14112 29200 14224 30000 0 FreeSans 448 90 0 0 chanx_left_in[7]
port 23 nsew signal input
flabel metal3 s 29200 28224 30000 28336 0 FreeSans 448 0 0 0 chanx_left_in[8]
port 24 nsew signal input
flabel metal2 s 16800 29200 16912 30000 0 FreeSans 448 90 0 0 chanx_left_in[9]
port 25 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chanx_left_out[0]
port 26 nsew signal tristate
flabel metal3 s 29200 22176 30000 22288 0 FreeSans 448 0 0 0 chanx_left_out[10]
port 27 nsew signal tristate
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chanx_left_out[11]
port 28 nsew signal tristate
flabel metal2 s 20160 29200 20272 30000 0 FreeSans 448 90 0 0 chanx_left_out[12]
port 29 nsew signal tristate
flabel metal3 s 29200 6048 30000 6160 0 FreeSans 448 0 0 0 chanx_left_out[13]
port 30 nsew signal tristate
flabel metal3 s 29200 26880 30000 26992 0 FreeSans 448 0 0 0 chanx_left_out[14]
port 31 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 chanx_left_out[15]
port 32 nsew signal tristate
flabel metal2 s 10752 29200 10864 30000 0 FreeSans 448 90 0 0 chanx_left_out[16]
port 33 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 chanx_left_out[17]
port 34 nsew signal tristate
flabel metal3 s 29200 5376 30000 5488 0 FreeSans 448 0 0 0 chanx_left_out[18]
port 35 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chanx_left_out[19]
port 36 nsew signal tristate
flabel metal3 s 29200 8064 30000 8176 0 FreeSans 448 0 0 0 chanx_left_out[1]
port 37 nsew signal tristate
flabel metal3 s 29200 7392 30000 7504 0 FreeSans 448 0 0 0 chanx_left_out[2]
port 38 nsew signal tristate
flabel metal3 s 29200 24192 30000 24304 0 FreeSans 448 0 0 0 chanx_left_out[3]
port 39 nsew signal tristate
flabel metal2 s 22176 29200 22288 30000 0 FreeSans 448 90 0 0 chanx_left_out[4]
port 40 nsew signal tristate
flabel metal2 s 10080 29200 10192 30000 0 FreeSans 448 90 0 0 chanx_left_out[5]
port 41 nsew signal tristate
flabel metal3 s 29200 20160 30000 20272 0 FreeSans 448 0 0 0 chanx_left_out[6]
port 42 nsew signal tristate
flabel metal3 s 29200 28896 30000 29008 0 FreeSans 448 0 0 0 chanx_left_out[7]
port 43 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chanx_left_out[8]
port 44 nsew signal tristate
flabel metal2 s 9408 29200 9520 30000 0 FreeSans 448 90 0 0 chanx_left_out[9]
port 45 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chanx_right_in[0]
port 46 nsew signal input
flabel metal3 s 29200 22848 30000 22960 0 FreeSans 448 0 0 0 chanx_right_in[10]
port 47 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chanx_right_in[11]
port 48 nsew signal input
flabel metal2 s 19488 29200 19600 30000 0 FreeSans 448 90 0 0 chanx_right_in[12]
port 49 nsew signal input
flabel metal3 s 29200 4704 30000 4816 0 FreeSans 448 0 0 0 chanx_right_in[13]
port 50 nsew signal input
flabel metal3 s 29200 19488 30000 19600 0 FreeSans 448 0 0 0 chanx_right_in[14]
port 51 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chanx_right_in[15]
port 52 nsew signal input
flabel metal2 s 4032 29200 4144 30000 0 FreeSans 448 90 0 0 chanx_right_in[16]
port 53 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chanx_right_in[17]
port 54 nsew signal input
flabel metal3 s 29200 4032 30000 4144 0 FreeSans 448 0 0 0 chanx_right_in[18]
port 55 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chanx_right_in[19]
port 56 nsew signal input
flabel metal3 s 29200 3360 30000 3472 0 FreeSans 448 0 0 0 chanx_right_in[1]
port 57 nsew signal input
flabel metal3 s 29200 2688 30000 2800 0 FreeSans 448 0 0 0 chanx_right_in[2]
port 58 nsew signal input
flabel metal3 s 29200 23520 30000 23632 0 FreeSans 448 0 0 0 chanx_right_in[3]
port 59 nsew signal input
flabel metal2 s 20832 29200 20944 30000 0 FreeSans 448 90 0 0 chanx_right_in[4]
port 60 nsew signal input
flabel metal2 s 6720 29200 6832 30000 0 FreeSans 448 90 0 0 chanx_right_in[5]
port 61 nsew signal input
flabel metal3 s 29200 18816 30000 18928 0 FreeSans 448 0 0 0 chanx_right_in[6]
port 62 nsew signal input
flabel metal3 s 29200 18144 30000 18256 0 FreeSans 448 0 0 0 chanx_right_in[7]
port 63 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chanx_right_in[8]
port 64 nsew signal input
flabel metal2 s 2688 29200 2800 30000 0 FreeSans 448 90 0 0 chanx_right_in[9]
port 65 nsew signal input
flabel metal2 s 11424 29200 11536 30000 0 FreeSans 448 90 0 0 chanx_right_out[0]
port 66 nsew signal tristate
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chanx_right_out[10]
port 67 nsew signal tristate
flabel metal3 s 29200 26208 30000 26320 0 FreeSans 448 0 0 0 chanx_right_out[11]
port 68 nsew signal tristate
flabel metal2 s 21504 29200 21616 30000 0 FreeSans 448 90 0 0 chanx_right_out[12]
port 69 nsew signal tristate
flabel metal2 s 12096 29200 12208 30000 0 FreeSans 448 90 0 0 chanx_right_out[13]
port 70 nsew signal tristate
flabel metal2 s 8064 29200 8176 30000 0 FreeSans 448 90 0 0 chanx_right_out[14]
port 71 nsew signal tristate
flabel metal2 s 18144 29200 18256 30000 0 FreeSans 448 90 0 0 chanx_right_out[15]
port 72 nsew signal tristate
flabel metal3 s 29200 24864 30000 24976 0 FreeSans 448 0 0 0 chanx_right_out[16]
port 73 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 chanx_right_out[17]
port 74 nsew signal tristate
flabel metal2 s 22848 29200 22960 30000 0 FreeSans 448 90 0 0 chanx_right_out[18]
port 75 nsew signal tristate
flabel metal2 s 5376 29200 5488 30000 0 FreeSans 448 90 0 0 chanx_right_out[19]
port 76 nsew signal tristate
flabel metal2 s 2016 29200 2128 30000 0 FreeSans 448 90 0 0 chanx_right_out[1]
port 77 nsew signal tristate
flabel metal2 s 12768 29200 12880 30000 0 FreeSans 448 90 0 0 chanx_right_out[2]
port 78 nsew signal tristate
flabel metal2 s 16128 29200 16240 30000 0 FreeSans 448 90 0 0 chanx_right_out[3]
port 79 nsew signal tristate
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chanx_right_out[4]
port 80 nsew signal tristate
flabel metal3 s 29200 27552 30000 27664 0 FreeSans 448 0 0 0 chanx_right_out[5]
port 81 nsew signal tristate
flabel metal3 s 29200 6720 30000 6832 0 FreeSans 448 0 0 0 chanx_right_out[6]
port 82 nsew signal tristate
flabel metal2 s 13440 29200 13552 30000 0 FreeSans 448 90 0 0 chanx_right_out[7]
port 83 nsew signal tristate
flabel metal3 s 29200 25536 30000 25648 0 FreeSans 448 0 0 0 chanx_right_out[8]
port 84 nsew signal tristate
flabel metal2 s 17472 29200 17584 30000 0 FreeSans 448 90 0 0 chanx_right_out[9]
port 85 nsew signal tristate
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 pReset
port 86 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 prog_clk
port 87 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 88 nsew signal tristate
flabel metal2 s 18816 29200 18928 30000 0 FreeSans 448 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 89 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 90 nsew signal tristate
flabel metal4 s 4586 3076 4906 26716 0 FreeSans 1280 90 0 0 vdd
port 91 nsew power bidirectional
flabel metal4 s 11390 3076 11710 26716 0 FreeSans 1280 90 0 0 vdd
port 91 nsew power bidirectional
flabel metal4 s 18194 3076 18514 26716 0 FreeSans 1280 90 0 0 vdd
port 91 nsew power bidirectional
flabel metal4 s 24998 3076 25318 26716 0 FreeSans 1280 90 0 0 vdd
port 91 nsew power bidirectional
flabel metal4 s 7988 3076 8308 26716 0 FreeSans 1280 90 0 0 vss
port 92 nsew ground bidirectional
flabel metal4 s 14792 3076 15112 26716 0 FreeSans 1280 90 0 0 vss
port 92 nsew ground bidirectional
flabel metal4 s 21596 3076 21916 26716 0 FreeSans 1280 90 0 0 vss
port 92 nsew ground bidirectional
flabel metal4 s 28400 3076 28720 26716 0 FreeSans 1280 90 0 0 vss
port 92 nsew ground bidirectional
rlabel metal1 14952 25872 14952 25872 0 vdd
rlabel via1 15032 26656 15032 26656 0 vss
rlabel metal2 10472 12376 10472 12376 0 _000_
rlabel metal3 7168 10808 7168 10808 0 _001_
rlabel metal2 7000 10976 7000 10976 0 _002_
rlabel metal2 5656 9408 5656 9408 0 _003_
rlabel metal2 2408 11312 2408 11312 0 _004_
rlabel metal2 4760 7728 4760 7728 0 _005_
rlabel metal2 6328 16464 6328 16464 0 _006_
rlabel metal2 2296 15904 2296 15904 0 _007_
rlabel metal2 2632 14560 2632 14560 0 _008_
rlabel metal3 4928 16632 4928 16632 0 _009_
rlabel metal2 12488 13720 12488 13720 0 _010_
rlabel metal2 11256 14280 11256 14280 0 _011_
rlabel metal2 16408 19432 16408 19432 0 _012_
rlabel metal2 14056 19768 14056 19768 0 _013_
rlabel metal2 12040 18424 12040 18424 0 _014_
rlabel metal2 10472 17864 10472 17864 0 _015_
rlabel metal2 8568 19208 8568 19208 0 _016_
rlabel metal2 8344 16520 8344 16520 0 _017_
rlabel metal2 15848 18200 15848 18200 0 _018_
rlabel metal2 12824 16464 12824 16464 0 _019_
rlabel metal2 23912 18200 23912 18200 0 _020_
rlabel metal2 24696 18816 24696 18816 0 _021_
rlabel metal2 23240 19208 23240 19208 0 _022_
rlabel metal2 20552 20188 20552 20188 0 _023_
rlabel metal2 24248 14112 24248 14112 0 _024_
rlabel metal2 25928 13720 25928 13720 0 _025_
rlabel metal2 24808 14728 24808 14728 0 _026_
rlabel metal2 22792 16464 22792 16464 0 _027_
rlabel metal2 20832 14728 20832 14728 0 _028_
rlabel metal3 19712 17416 19712 17416 0 _029_
rlabel metal2 22792 8792 22792 8792 0 _030_
rlabel metal2 25816 7224 25816 7224 0 _031_
rlabel metal2 24472 10360 24472 10360 0 _032_
rlabel metal2 22344 10976 22344 10976 0 _033_
rlabel metal2 23800 11144 23800 11144 0 _034_
rlabel metal2 24192 9352 24192 9352 0 _035_
rlabel metal2 25368 5152 25368 5152 0 _036_
rlabel metal2 22232 7840 22232 7840 0 _037_
rlabel metal2 19320 8736 19320 8736 0 _038_
rlabel metal2 17976 8008 17976 8008 0 _039_
rlabel metal2 15848 9240 15848 9240 0 _040_
rlabel metal2 13720 9464 13720 9464 0 _041_
rlabel metal2 16184 8848 16184 8848 0 _042_
rlabel metal2 2072 14392 2072 14392 0 _043_
rlabel metal2 15736 18816 15736 18816 0 _044_
rlabel metal3 27664 14504 27664 14504 0 _045_
rlabel metal2 21448 8176 21448 8176 0 _046_
rlabel metal3 1302 10808 1302 10808 0 ccff_head
rlabel metal3 28490 8792 28490 8792 0 ccff_tail
rlabel metal2 1848 25984 1848 25984 0 chanx_left_in[0]
rlabel metal2 10808 1246 10808 1246 0 chanx_left_in[10]
rlabel metal2 28168 21224 28168 21224 0 chanx_left_in[11]
rlabel metal2 24192 26488 24192 26488 0 chanx_left_in[12]
rlabel metal2 9016 25536 9016 25536 0 chanx_left_in[13]
rlabel metal2 3304 25200 3304 25200 0 chanx_left_in[14]
rlabel metal2 15512 27874 15512 27874 0 chanx_left_in[15]
rlabel metal2 23128 24920 23128 24920 0 chanx_left_in[16]
rlabel metal2 1736 23688 1736 23688 0 chanx_left_in[17]
rlabel metal2 23632 25480 23632 25480 0 chanx_left_in[18]
rlabel metal2 7448 28070 7448 28070 0 chanx_left_in[19]
rlabel metal2 6104 28070 6104 28070 0 chanx_left_in[1]
rlabel metal2 4760 26208 4760 26208 0 chanx_left_in[2]
rlabel metal2 14840 28070 14840 28070 0 chanx_left_in[3]
rlabel metal2 18312 4200 18312 4200 0 chanx_left_in[4]
rlabel metal3 28378 21560 28378 21560 0 chanx_left_in[5]
rlabel metal2 20216 3192 20216 3192 0 chanx_left_in[6]
rlabel metal2 14392 27048 14392 27048 0 chanx_left_in[7]
rlabel metal2 25480 25480 25480 25480 0 chanx_left_in[8]
rlabel metal2 16856 27426 16856 27426 0 chanx_left_in[9]
rlabel metal2 16184 2198 16184 2198 0 chanx_left_out[0]
rlabel metal3 28658 22232 28658 22232 0 chanx_left_out[10]
rlabel metal2 9800 2464 9800 2464 0 chanx_left_out[11]
rlabel metal2 21224 26488 21224 26488 0 chanx_left_out[12]
rlabel metal2 24248 5320 24248 5320 0 chanx_left_out[13]
rlabel metal2 25928 26264 25928 26264 0 chanx_left_out[14]
rlabel metal2 12824 2478 12824 2478 0 chanx_left_out[15]
rlabel metal2 10808 28070 10808 28070 0 chanx_left_out[16]
rlabel metal2 15512 2198 15512 2198 0 chanx_left_out[17]
rlabel metal2 23240 4424 23240 4424 0 chanx_left_out[18]
rlabel metal2 18872 854 18872 854 0 chanx_left_out[19]
rlabel metal2 27776 5320 27776 5320 0 chanx_left_out[1]
rlabel metal2 27384 5600 27384 5600 0 chanx_left_out[2]
rlabel metal2 28056 24416 28056 24416 0 chanx_left_out[3]
rlabel metal2 22904 26208 22904 26208 0 chanx_left_out[4]
rlabel metal2 10360 27272 10360 27272 0 chanx_left_out[5]
rlabel metal2 28056 20440 28056 20440 0 chanx_left_out[6]
rlabel metal2 27776 24136 27776 24136 0 chanx_left_out[7]
rlabel metal2 13496 854 13496 854 0 chanx_left_out[8]
rlabel metal3 9968 24920 9968 24920 0 chanx_left_out[9]
rlabel metal2 14840 910 14840 910 0 chanx_right_in[0]
rlabel metal2 26824 22288 26824 22288 0 chanx_right_in[10]
rlabel metal2 10136 854 10136 854 0 chanx_right_in[11]
rlabel metal2 20216 25536 20216 25536 0 chanx_right_in[12]
rlabel metal3 26824 4536 26824 4536 0 chanx_right_in[13]
rlabel metal2 28168 19768 28168 19768 0 chanx_right_in[14]
rlabel metal2 11816 3864 11816 3864 0 chanx_right_in[15]
rlabel metal2 4088 26096 4088 26096 0 chanx_right_in[16]
rlabel metal2 16856 2478 16856 2478 0 chanx_right_in[17]
rlabel metal2 24696 3864 24696 3864 0 chanx_right_in[18]
rlabel metal2 18424 3360 18424 3360 0 chanx_right_in[19]
rlabel metal3 26698 3416 26698 3416 0 chanx_right_in[1]
rlabel metal2 20888 3136 20888 3136 0 chanx_right_in[2]
rlabel metal2 24696 24248 24696 24248 0 chanx_right_in[3]
rlabel metal2 20888 27426 20888 27426 0 chanx_right_in[4]
rlabel metal2 6776 28070 6776 28070 0 chanx_right_in[5]
rlabel metal2 28168 19040 28168 19040 0 chanx_right_in[6]
rlabel metal2 27720 18256 27720 18256 0 chanx_right_in[7]
rlabel metal2 12152 1246 12152 1246 0 chanx_right_in[8]
rlabel metal2 2744 27202 2744 27202 0 chanx_right_in[9]
rlabel metal2 12152 25816 12152 25816 0 chanx_right_out[0]
rlabel metal2 7952 3304 7952 3304 0 chanx_right_out[10]
rlabel metal2 26152 25424 26152 25424 0 chanx_right_out[11]
rlabel metal2 22792 26488 22792 26488 0 chanx_right_out[12]
rlabel metal2 12152 28070 12152 28070 0 chanx_right_out[13]
rlabel metal2 8008 27720 8008 27720 0 chanx_right_out[14]
rlabel metal2 18872 26096 18872 26096 0 chanx_right_out[15]
rlabel metal2 27720 25088 27720 25088 0 chanx_right_out[16]
rlabel metal3 1470 24920 1470 24920 0 chanx_right_out[17]
rlabel metal2 25032 26488 25032 26488 0 chanx_right_out[18]
rlabel metal2 5656 26152 5656 26152 0 chanx_right_out[19]
rlabel metal2 2632 26600 2632 26600 0 chanx_right_out[1]
rlabel metal2 13944 25648 13944 25648 0 chanx_right_out[2]
rlabel metal2 17416 26320 17416 26320 0 chanx_right_out[3]
rlabel metal2 14280 3304 14280 3304 0 chanx_right_out[4]
rlabel metal2 27496 25312 27496 25312 0 chanx_right_out[5]
rlabel metal2 25704 5152 25704 5152 0 chanx_right_out[6]
rlabel metal2 14168 26488 14168 26488 0 chanx_right_out[7]
rlabel metal2 27720 25872 27720 25872 0 chanx_right_out[8]
rlabel metal2 18984 26488 18984 26488 0 chanx_right_out[9]
rlabel metal2 22008 13720 22008 13720 0 clknet_0_prog_clk
rlabel metal2 2072 7336 2072 7336 0 clknet_2_0__leaf_prog_clk
rlabel metal3 4368 16856 4368 16856 0 clknet_2_1__leaf_prog_clk
rlabel metal2 22680 5880 22680 5880 0 clknet_2_2__leaf_prog_clk
rlabel metal2 27720 13664 27720 13664 0 clknet_2_3__leaf_prog_clk
rlabel metal2 5544 8008 5544 8008 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal3 2184 11256 2184 11256 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal3 7112 8120 7112 8120 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal2 7560 10024 7560 10024 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal2 5544 12376 5544 12376 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal2 15848 10920 15848 10920 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal3 8064 13160 8064 13160 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel metal3 14280 14392 14280 14392 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal3 4312 14392 4312 14392 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel metal2 2408 12824 2408 12824 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal2 2744 16296 2744 16296 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal2 7112 15736 7112 15736 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal2 9072 17080 9072 17080 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal3 10024 15960 10024 15960 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal2 11256 18200 11256 18200 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal2 13048 20552 13048 20552 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal3 16352 20664 16352 20664 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal3 19096 19096 19096 19096 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal3 22344 19992 22344 19992 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal2 25480 20412 25480 20412 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal2 25928 18760 25928 18760 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal3 23688 16968 23688 16968 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal2 12040 15736 12040 15736 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 16968 18480 16968 18480 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal2 19880 16688 19880 16688 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal2 27272 16240 27272 16240 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal2 27272 14448 27272 14448 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal2 25592 15176 25592 15176 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal3 27048 12264 27048 12264 0 mem_top_ipin_1.DFFR_4_.Q
rlabel metal2 26376 11592 26376 11592 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal3 25424 9128 25424 9128 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal2 19768 13104 19768 13104 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal3 25200 10696 25200 10696 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal3 26096 7560 26096 7560 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal3 26936 4424 26936 4424 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal2 21112 7840 21112 7840 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal2 14280 6888 14280 6888 0 mem_top_ipin_3.DFFR_0_.Q
rlabel metal2 20440 9352 20440 9352 0 mem_top_ipin_3.DFFR_1_.Q
rlabel metal2 20328 6328 20328 6328 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal3 22064 7224 22064 7224 0 mem_top_ipin_3.DFFR_3_.Q
rlabel metal2 27272 6384 27272 6384 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal2 2408 7924 2408 7924 0 net1
rlabel metal2 3752 24248 3752 24248 0 net10
rlabel metal3 18760 8344 18760 8344 0 net100
rlabel metal2 12376 20720 12376 20720 0 net101
rlabel metal2 19880 12096 19880 12096 0 net102
rlabel metal2 8232 17528 8232 17528 0 net103
rlabel metal3 23688 20888 23688 20888 0 net104
rlabel metal2 7896 12208 7896 12208 0 net105
rlabel metal2 22568 14056 22568 14056 0 net106
rlabel metal2 22008 10136 22008 10136 0 net107
rlabel metal2 20776 19152 20776 19152 0 net108
rlabel metal2 18648 16520 18648 16520 0 net109
rlabel metal2 20552 24584 20552 24584 0 net11
rlabel metal3 26768 17640 26768 17640 0 net110
rlabel metal2 23688 13832 23688 13832 0 net111
rlabel metal2 8008 13776 8008 13776 0 net112
rlabel metal2 23128 5432 23128 5432 0 net113
rlabel metal2 6104 16520 6104 16520 0 net114
rlabel metal2 19992 6608 19992 6608 0 net115
rlabel metal3 23408 15288 23408 15288 0 net116
rlabel metal2 10024 18760 10024 18760 0 net117
rlabel metal2 12936 8456 12936 8456 0 net118
rlabel metal2 4872 10584 4872 10584 0 net119
rlabel metal2 11928 24640 11928 24640 0 net12
rlabel metal2 8456 11032 8456 11032 0 net120
rlabel metal2 3976 15736 3976 15736 0 net121
rlabel metal2 8680 14560 8680 14560 0 net122
rlabel metal3 25312 8792 25312 8792 0 net123
rlabel metal2 6104 18872 6104 18872 0 net124
rlabel metal2 23352 6776 23352 6776 0 net125
rlabel metal2 3472 9016 3472 9016 0 net126
rlabel metal2 3920 9912 3920 9912 0 net127
rlabel metal3 27104 9912 27104 9912 0 net128
rlabel metal2 11256 7112 11256 7112 0 net129
rlabel metal2 9800 24304 9800 24304 0 net13
rlabel metal2 22904 12040 22904 12040 0 net130
rlabel metal2 22904 16128 22904 16128 0 net131
rlabel metal3 7616 23240 7616 23240 0 net14
rlabel metal2 15624 24584 15624 24584 0 net15
rlabel metal2 18088 4816 18088 4816 0 net16
rlabel metal3 25816 21672 25816 21672 0 net17
rlabel metal2 20608 4424 20608 4424 0 net18
rlabel metal2 13832 24360 13832 24360 0 net19
rlabel metal2 2072 24472 2072 24472 0 net2
rlabel metal2 25928 24360 25928 24360 0 net20
rlabel metal2 16520 24584 16520 24584 0 net21
rlabel metal2 15288 4760 15288 4760 0 net22
rlabel metal2 26488 22120 26488 22120 0 net23
rlabel metal2 10360 4592 10360 4592 0 net24
rlabel metal2 19880 24584 19880 24584 0 net25
rlabel metal2 22232 4256 22232 4256 0 net26
rlabel metal3 26208 20104 26208 20104 0 net27
rlabel metal3 11368 3304 11368 3304 0 net28
rlabel metal2 10696 25032 10696 25032 0 net29
rlabel metal2 10920 4200 10920 4200 0 net3
rlabel metal2 13496 4704 13496 4704 0 net30
rlabel metal2 22120 3640 22120 3640 0 net31
rlabel metal2 18592 4536 18592 4536 0 net32
rlabel metal2 21784 3584 21784 3584 0 net33
rlabel metal2 21168 3416 21168 3416 0 net34
rlabel metal2 24080 23912 24080 23912 0 net35
rlabel metal2 21448 24584 21448 24584 0 net36
rlabel metal2 10976 23128 10976 23128 0 net37
rlabel metal3 26656 21224 26656 21224 0 net38
rlabel metal2 25536 21672 25536 21672 0 net39
rlabel metal3 27048 21784 27048 21784 0 net4
rlabel metal2 12320 3416 12320 3416 0 net40
rlabel metal2 8456 24584 8456 24584 0 net41
rlabel metal2 9968 4424 9968 4424 0 net42
rlabel metal2 26152 5880 26152 5880 0 net43
rlabel metal2 14728 4200 14728 4200 0 net44
rlabel metal2 26264 23016 26264 23016 0 net45
rlabel metal2 10472 4200 10472 4200 0 net46
rlabel metal2 20468 26264 20468 26264 0 net47
rlabel metal3 22960 4424 22960 4424 0 net48
rlabel metal2 24920 24136 24920 24136 0 net49
rlabel metal2 20664 23184 20664 23184 0 net5
rlabel metal2 11592 4704 11592 4704 0 net50
rlabel metal2 10360 25032 10360 25032 0 net51
rlabel metal2 15176 4200 15176 4200 0 net52
rlabel metal2 22904 3808 22904 3808 0 net53
rlabel metal2 18984 4200 18984 4200 0 net54
rlabel metal2 26936 5544 26936 5544 0 net55
rlabel metal2 26600 4088 26600 4088 0 net56
rlabel metal2 24248 23968 24248 23968 0 net57
rlabel metal2 21672 24360 21672 24360 0 net58
rlabel metal2 10920 23912 10920 23912 0 net59
rlabel metal2 11032 24472 11032 24472 0 net6
rlabel metal2 25928 21448 25928 21448 0 net60
rlabel metal2 25648 23352 25648 23352 0 net61
rlabel metal2 12264 4704 12264 4704 0 net62
rlabel metal2 8680 24304 8680 24304 0 net63
rlabel metal2 10024 24640 10024 24640 0 net64
rlabel metal2 8624 3528 8624 3528 0 net65
rlabel metal2 26600 23464 26600 23464 0 net66
rlabel metal2 20888 24024 20888 24024 0 net67
rlabel metal2 11312 23800 11312 23800 0 net68
rlabel metal2 9016 23632 9016 23632 0 net69
rlabel metal2 9240 24808 9240 24808 0 net7
rlabel metal2 15288 24528 15288 24528 0 net70
rlabel metal2 25592 24528 25592 24528 0 net71
rlabel metal2 3528 25088 3528 25088 0 net72
rlabel metal2 20776 24584 20776 24584 0 net73
rlabel metal3 9296 23800 9296 23800 0 net74
rlabel metal2 9576 24808 9576 24808 0 net75
rlabel metal2 10584 23408 10584 23408 0 net76
rlabel metal2 15960 24808 15960 24808 0 net77
rlabel metal2 13608 4200 13608 4200 0 net78
rlabel metal3 25816 23240 25816 23240 0 net79
rlabel metal2 15176 25200 15176 25200 0 net8
rlabel metal2 25032 3640 25032 3640 0 net80
rlabel metal2 13552 23800 13552 23800 0 net81
rlabel metal2 26264 25032 26264 25032 0 net82
rlabel metal2 16856 24584 16856 24584 0 net83
rlabel metal2 7448 2030 7448 2030 0 net84
rlabel metal2 6776 2030 6776 2030 0 net85
rlabel metal3 25536 26488 25536 26488 0 net86
rlabel metal2 26656 4872 26656 4872 0 net87
rlabel metal3 1582 24248 1582 24248 0 net88
rlabel metal2 20104 26656 20104 26656 0 net89
rlabel metal3 24304 23912 24304 23912 0 net9
rlabel metal3 1246 6104 1246 6104 0 net90
rlabel metal3 17248 8904 17248 8904 0 net91
rlabel metal2 12264 11704 12264 11704 0 net92
rlabel metal3 24136 13720 24136 13720 0 net93
rlabel metal2 18088 19656 18088 19656 0 net94
rlabel metal2 16856 17920 16856 17920 0 net95
rlabel metal2 4536 16856 4536 16856 0 net96
rlabel metal2 4088 14168 4088 14168 0 net97
rlabel metal2 13944 17864 13944 17864 0 net98
rlabel metal2 16296 20552 16296 20552 0 net99
rlabel metal2 9464 854 9464 854 0 pReset
rlabel metal2 15288 12656 15288 12656 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
