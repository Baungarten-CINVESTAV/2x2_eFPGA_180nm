* NGSPICE file created from sb_2__1_.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

.subckt sb_2__1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18]
+ chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[10]
+ chany_bottom_out[11] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[9] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
+ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ pReset prog_clk top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ vdd vss chany_bottom_out[8]
+ chanx_left_out[8] chany_bottom_out[12] chany_bottom_out[16] chanx_left_out[9] chany_top_out[0]
+ chanx_left_out[10] chany_top_out[4] chanx_left_out[11] chany_top_out[8] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chany_top_out[16] chanx_left_out[15] chany_bottom_out[0]
+ chany_bottom_out[4] chanx_left_out[7]
XFILLER_0_17_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_294_ net109 _050_ clknet_3_3__leaf_prog_clk mem_bottom_track_17.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_346_ net191 _102_ clknet_3_5__leaf_prog_clk mem_left_track_15.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_11_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_277_ net118 _033_ clknet_3_4__leaf_prog_clk mem_top_track_24.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input36_I pReset vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_200_ _110_ _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_131_ _111_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xsb_2__1__82 chanx_left_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__93 chanx_left_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_329_ net138 _085_ clknet_3_7__leaf_prog_clk mem_left_track_7.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_10_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold63 mem_top_track_24.DFFR_4_.Q net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold52 mem_top_track_24.DFFR_1_.Q net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold74 mem_bottom_track_1.DFFR_1_.Q net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold30 mem_left_track_5.DFFR_1_.Q net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold41 mem_left_track_7.DFFR_1_.Q net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold96 mem_bottom_track_1.DFFR_6_.Q net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__167__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold85 mem_left_track_3.DFFR_3_.Q net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__247__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput64 net64 chany_top_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput53 net53 chany_bottom_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput42 net42 chany_bottom_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_3_7__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_293_ net119 _049_ clknet_3_2__leaf_prog_clk mem_bottom_track_17.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_23_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_276_ net145 _032_ clknet_3_4__leaf_prog_clk mem_top_track_24.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_345_ net101 _101_ clknet_3_5__leaf_prog_clk mem_left_track_13.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_11_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input29_I chany_top_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_4_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_130_ _111_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xsb_2__1__94 chanx_left_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_259_ net200 _015_ clknet_3_2__leaf_prog_clk mem_bottom_track_1.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ net146 _084_ clknet_3_7__leaf_prog_clk mem_left_track_7.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xsb_2__1__83 chanx_left_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__72 chany_top_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_10_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold75 mem_top_track_24.DFFR_2_.Q net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold20 mem_top_track_8.DFFR_1_.Q net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 mem_top_track_0.DFFR_5_.Q net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold64 mem_top_track_16.DFFR_0_.D net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 mem_left_track_21.DFFR_1_.Q net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 mem_left_track_1.DFFR_5_.Q net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold97 mem_bottom_track_33.DFFR_0_.Q net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold31 mem_bottom_track_17.DFFR_5_.Q net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_7_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input11_I chany_bottom_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput65 net65 chany_top_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput54 net54 chany_bottom_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput43 net43 chany_bottom_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_33_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__178__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I chany_bottom_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_292_ net199 _048_ clknet_3_2__leaf_prog_clk mem_bottom_track_17.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_23_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_413_ net2 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_344_ net186 _100_ clknet_3_5__leaf_prog_clk mem_left_track_13.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_275_ net149 _031_ clknet_3_4__leaf_prog_clk mem_top_track_24.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_20_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsb_2__1__95 chanx_left_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_9_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_2__1__84 chanx_left_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__73 chany_top_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_258_ net104 _014_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_189_ _110_ _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_327_ net163 _083_ clknet_3_7__leaf_prog_clk mem_left_track_7.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__270__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold76 mem_top_track_8.DFFR_0_.Q net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold32 mem_left_track_15.DFFR_1_.Q net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold21 mem_top_track_16.DFFR_5_.Q net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold54 mem_left_track_1.DFFR_0_.Q net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold43 mem_bottom_track_17.DFFR_0_.D net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold98 mem_bottom_track_17.DFFR_3_.Q net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 mem_bottom_track_33.DFFR_4_.Q net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 mem_bottom_track_25.DFFR_4_.Q net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 mem_left_track_7.DFFR_4_.Q net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_8_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput55 net55 chany_bottom_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput66 net66 chany_top_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput44 net44 chany_bottom_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_291_ net195 _047_ clknet_3_2__leaf_prog_clk mem_bottom_track_17.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_31_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__189__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_412_ net10 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_274_ net172 _030_ clknet_3_4__leaf_prog_clk mem_top_track_24.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_343_ net126 _099_ clknet_3_7__leaf_prog_clk mem_left_track_27.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_326_ net162 _082_ clknet_3_7__leaf_prog_clk mem_left_track_7.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_257_ net171 _013_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_188_ _116_ _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xsb_2__1__74 chany_top_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__96 chanx_left_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__85 chanx_left_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_0_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input34_I chany_top_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_309_ net158 _065_ clknet_3_3__leaf_prog_clk mem_left_track_1.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold22 mem_bottom_track_17.DFFR_1_.Q net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold11 mem_left_track_5.DFFR_5_.Q net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 mem_top_track_16.DFFR_0_.Q net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold44 mem_top_track_8.DFFR_2_.Q net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 mem_top_track_32.DFFR_3_.Q net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 mem_left_track_3.DFFR_0_.Q net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold99 mem_left_track_3.DFFR_4_.Q net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 mem_left_track_5.DFFR_3_.Q net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 mem_left_track_7.DFFR_3_.Q net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_38_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput56 net56 chany_bottom_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput45 net45 chany_bottom_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_9_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput67 net67 chany_top_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__260__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_290_ net169 _046_ clknet_3_2__leaf_prog_clk mem_bottom_track_17.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_8_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_342_ net99 _098_ clknet_3_5__leaf_prog_clk mem_left_track_27.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_411_ net11 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_273_ net134 _029_ clknet_3_1__leaf_prog_clk mem_top_track_24.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_325_ net106 _081_ clknet_3_7__leaf_prog_clk mem_left_track_5.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xsb_2__1__75 chany_top_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__97 chanx_left_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_256_ net121 _012_ clknet_3_1__leaf_prog_clk mem_bottom_track_1.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_187_ _116_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xsb_2__1__86 chanx_left_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input27_I chany_top_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_239_ _121_ _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_308_ net120 _064_ clknet_3_6__leaf_prog_clk mem_left_track_1.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_30_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold45 mem_bottom_track_1.DFFR_7_.Q net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold23 mem_left_track_1.DFFR_4_.Q net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold56 mem_left_track_1.DFFR_2_.Q net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold12 mem_bottom_track_17.DFFR_0_.Q net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 mem_bottom_track_25.DFFR_1_.Q net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold89 mem_left_track_13.DFFR_0_.Q net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold67 mem_top_track_16.DFFR_4_.Q net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold78 mem_bottom_track_9.DFFR_4_.Q net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_38_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput46 net46 chany_bottom_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput57 net57 chany_top_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput68 net68 chany_top_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input1_I ccff_head vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__250__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_410_ net12 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_272_ net160 _028_ clknet_3_1__leaf_prog_clk mem_top_track_24.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_341_ net136 _097_ clknet_3_5__leaf_prog_clk mem_left_track_25.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_42_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__273__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xsb_2__1__87 chanx_left_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__76 chany_top_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_255_ net102 _011_ clknet_3_3__leaf_prog_clk mem_bottom_track_1.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_324_ net155 _080_ clknet_3_7__leaf_prog_clk mem_left_track_5.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_24_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_186_ _116_ _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_0_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_238_ _121_ _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_24_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_169_ _115_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_307_ net143 _063_ clknet_3_3__leaf_prog_clk mem_bottom_track_33.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold35 mem_top_track_16.DFFR_1_.Q net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 mem_left_track_17.DFFR_0_.Q net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold57 mem_top_track_0.DFFR_3_.Q net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold24 mem_bottom_track_1.DFFR_2_.Q net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 mem_left_track_5.DFFR_2_.Q net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 mem_bottom_track_25.DFFR_5_.Q net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold13 mem_bottom_track_25.DFFR_3_.Q net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput47 net47 chany_bottom_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput58 net58 chany_top_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput69 net69 chany_top_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_271_ net161 _027_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_340_ net190 _096_ clknet_3_5__leaf_prog_clk mem_left_track_25.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__200__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_2__1__88 chanx_left_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__77 chany_bottom_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_254_ net113 _010_ clknet_3_1__leaf_prog_clk mem_bottom_track_1.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_323_ net127 _079_ clknet_3_6__leaf_prog_clk mem_left_track_5.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_185_ _116_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_306_ net194 _062_ clknet_3_3__leaf_prog_clk mem_bottom_track_33.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_12_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_237_ _121_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__263__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_168_ _115_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input32_I chany_top_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold36 mem_top_track_8.DFFR_4_.Q net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 mem_top_track_0.DFFR_7_.Q net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 mem_left_track_19.DFFR_0_.Q net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold14 mem_bottom_track_9.DFFR_1_.Q net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold47 mem_left_track_3.DFFR_2_.Q net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold58 mem_left_track_5.DFFR_0_.Q net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__286__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput48 net48 chany_bottom_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput59 net59 chany_top_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput37 net37 ccff_tail vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_4_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold100 mem_left_track_7.DFFR_5_.Q net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_5_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_270_ net185 _026_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_42_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_399_ net9 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_322_ net165 _078_ clknet_3_6__leaf_prog_clk mem_left_track_5.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xsb_2__1__78 chany_bottom_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__89 chanx_left_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_10_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_253_ net202 _009_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_6_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_184_ _116_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_15_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__211__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_305_ net180 _061_ clknet_3_3__leaf_prog_clk mem_bottom_track_33.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_236_ _121_ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_167_ _110_ _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_24_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold37 mem_top_track_24.DFFR_3_.Q net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold59 mem_bottom_track_9.DFFR_2_.Q net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 mem_top_track_24.DFFR_0_.Q net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold26 mem_top_track_32.DFFR_2_.Q net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold15 mem_left_track_11.DFFR_0_.Q net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input25_I chany_top_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_219_ _119_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput49 net49 chany_bottom_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput38 net38 chanx_left_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__253__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold101 mem_left_track_27.DFFR_1_.Q net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_5_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_398_ net17 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_252_ net193 _008_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_7_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_321_ net130 _077_ clknet_3_6__leaf_prog_clk mem_left_track_5.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xsb_2__1__79 chany_bottom_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_10_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_183_ _116_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_235_ _121_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_304_ net115 _060_ clknet_3_6__leaf_prog_clk mem_bottom_track_33.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_166_ _114_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_11_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold38 mem_top_track_0.DFFR_6_.Q net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold16 mem_bottom_track_1.DFFR_4_.Q net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__222__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold27 mem_bottom_track_33.DFFR_3_.Q net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input18_I chany_top_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold49 mem_left_track_7.DFFR_2_.Q net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_3_1__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_149_ _113_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_218_ _119_ _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput39 net39 chanx_left_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_17_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold102 mem_bottom_track_17.DFFR_2_.Q net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_5_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_397_ net28 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__266__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_18_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__289__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_251_ net1 _007_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_182_ _116_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_320_ net178 _076_ clknet_3_6__leaf_prog_clk mem_left_track_5.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_234_ _121_ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_165_ _114_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_303_ net124 _059_ clknet_3_2__leaf_prog_clk mem_bottom_track_33.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold17 mem_top_track_16.DFFR_2_.Q net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold39 mem_left_track_23.DFFR_1_.Q net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 mem_bottom_track_9.DFFR_3_.Q net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_148_ _113_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_217_ _119_ _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input30_I chany_top_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold103 mem_bottom_track_1.DFFR_0_.D net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_396_ net29 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_250_ net203 _006_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_181_ _116_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__256__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_302_ net107 _058_ clknet_3_3__leaf_prog_clk mem_bottom_track_33.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_233_ net36 _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_164_ _114_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold29 mem_left_track_25.DFFR_1_.Q net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold18 mem_bottom_track_33.DFFR_2_.Q net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_147_ _113_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_216_ _119_ _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input23_I chany_top_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold104 mem_top_track_0.DFFR_2_.Q net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_13_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_395_ net30 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_180_ _116_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_232_ _120_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_301_ net128 _057_ clknet_3_2__leaf_prog_clk mem_bottom_track_25.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_163_ _114_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold19 mem_top_track_24.DFFR_5_.Q net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_215_ _119_ _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_146_ _113_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__246__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I chany_bottom_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__269__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I chany_bottom_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_129_ _111_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_17_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold105 mem_bottom_track_1.DFFR_5_.Q net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_394_ net31 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_162_ _114_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_231_ _120_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_300_ net137 _056_ clknet_3_2__leaf_prog_clk mem_bottom_track_25.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 ccff_head net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_0_prog_clk prog_clk clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_145_ _110_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_214_ _119_ _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_128_ _111_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold106 mem_top_track_0.DFFR_0_.Q net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_393_ net32 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_161_ _114_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_230_ _120_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput2 chany_bottom_in[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_144_ _112_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_213_ _119_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_28_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_127_ _111_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_25_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input21_I chany_top_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold107 mem_left_track_19.DFFR_1_.Q net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_6__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_392_ net34 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__249__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_160_ _114_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_17_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_289_ net142 _045_ clknet_3_0__leaf_prog_clk mem_bottom_track_9.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 chany_bottom_in[10] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_40_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_212_ _119_ _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_143_ _112_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_126_ _111_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_16_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input14_I chany_bottom_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold108 mem_left_track_17.DFFR_1_.Q net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__282__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I chany_bottom_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_391_ net35 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_288_ net177 _044_ clknet_3_2__leaf_prog_clk mem_bottom_track_9.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 chany_bottom_in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_142_ _112_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_211_ _110_ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_409_ net13 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_125_ _111_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_39_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold109 mem_top_track_0.DFFR_1_.Q net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_8_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_390_ net18 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__272__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_287_ net111 _043_ clknet_3_0__leaf_prog_clk mem_bottom_track_9.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput5 chany_bottom_in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_141_ _112_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_210_ _118_ _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_408_ net14 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_339_ net150 _095_ clknet_3_5__leaf_prog_clk mem_left_track_23.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_36_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_124_ _111_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_0_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput30 chany_top_in[4] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_17_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_286_ net156 _042_ clknet_3_0__leaf_prog_clk mem_bottom_track_9.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput6 chany_bottom_in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__262__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_140_ _112_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_407_ net15 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_338_ net187 _094_ clknet_3_5__leaf_prog_clk mem_left_track_23.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_269_ net132 _025_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_123_ _110_ _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_33_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 chany_top_in[5] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 chany_top_in[12] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_3__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input12_I chany_bottom_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input4_I chany_bottom_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_285_ net125 _041_ clknet_3_2__leaf_prog_clk mem_bottom_track_9.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_1_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 chany_bottom_in[16] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_406_ net16 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_337_ net204 _093_ clknet_3_4__leaf_prog_clk mem_left_track_21.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_268_ net114 _024_ clknet_3_4__leaf_prog_clk mem_top_track_16.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_199_ _117_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_122_ net36 _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__252__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput32 chany_top_in[6] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 chany_top_in[13] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput10 chany_bottom_in[1] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_353_ net198 _109_ clknet_3_5__leaf_prog_clk mem_left_track_29.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_284_ net175 _040_ clknet_3_2__leaf_prog_clk mem_bottom_track_17.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput8 chany_bottom_in[17] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_405_ net3 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_267_ net100 _023_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_336_ net98 _092_ clknet_3_5__leaf_prog_clk mem_left_track_21.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_198_ _117_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_6_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input35_I chany_top_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 chany_top_in[7] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 chany_top_in[14] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_319_ net139 _075_ clknet_3_6__leaf_prog_clk mem_left_track_3.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput11 chany_bottom_in[2] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_7_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__265__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_352_ net170 _108_ clknet_3_5__leaf_prog_clk net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_283_ net116 _039_ clknet_3_4__leaf_prog_clk mem_top_track_32.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput9 chany_bottom_in[18] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_404_ net4 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_266_ net164 _022_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_197_ _117_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_335_ net167 _091_ clknet_3_7__leaf_prog_clk mem_left_track_11.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_22_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input28_I chany_top_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_249_ net206 _005_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput23 chany_top_in[15] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 chany_bottom_in[4] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_318_ net174 _074_ clknet_3_6__leaf_prog_clk mem_left_track_3.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput34 chany_top_in[8] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_7_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold1 mem_left_track_21.DFFR_0_.Q net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input10_I chany_bottom_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I chany_bottom_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_351_ net205 _107_ clknet_3_5__leaf_prog_clk mem_left_track_19.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_282_ net103 _038_ clknet_3_1__leaf_prog_clk mem_top_track_32.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_1_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_403_ net5 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_334_ net112 _090_ clknet_3_4__leaf_prog_clk mem_left_track_11.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_265_ net122 _021_ clknet_3_1__leaf_prog_clk mem_top_track_8.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_196_ _117_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_22_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 chany_bottom_in[5] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_317_ net188 _073_ clknet_3_6__leaf_prog_clk mem_left_track_3.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput24 chany_top_in[16] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_248_ net201 _004_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput35 chany_top_in[9] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_179_ _116_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_24_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold2 mem_left_track_27.DFFR_0_.Q net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_32_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_350_ net166 _106_ clknet_3_5__leaf_prog_clk mem_left_track_19.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_281_ net105 _037_ clknet_3_3__leaf_prog_clk mem_top_track_32.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_402_ net6 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_264_ net173 _020_ clknet_3_1__leaf_prog_clk mem_top_track_8.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_333_ net197 _089_ clknet_3_7__leaf_prog_clk mem_left_track_9.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_195_ _117_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_19_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__245__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput14 chany_bottom_in[6] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_247_ net154 _003_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput36 pReset net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_316_ net144 _072_ clknet_3_6__leaf_prog_clk mem_left_track_3.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput25 chany_top_in[17] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_178_ _110_ _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input33_I chany_top_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold3 mem_top_track_16.DFFR_3_.Q net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_280_ net123 _036_ clknet_3_4__leaf_prog_clk mem_top_track_32.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_401_ net7 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_263_ net117 _019_ clknet_3_0__leaf_prog_clk mem_top_track_8.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_332_ net157 _088_ clknet_3_7__leaf_prog_clk mem_left_track_11.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_36_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_194_ _117_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_19_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput26 chany_top_in[18] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput15 chany_bottom_in[8] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_246_ net168 _002_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_315_ net182 _071_ clknet_3_6__leaf_prog_clk mem_left_track_3.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_177_ _115_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_15_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input26_I chany_top_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_229_ _120_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk clknet_3_7__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_4_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold4 mem_left_track_11.DFFR_1_.Q net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__258__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_prog_clk_I prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ net8 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_331_ net108 _087_ clknet_3_7__leaf_prog_clk mem_left_track_7.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_262_ net141 _018_ clknet_3_0__leaf_prog_clk mem_top_track_8.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_193_ _117_ _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_42_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_314_ net196 _070_ clknet_3_6__leaf_prog_clk mem_left_track_3.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput27 chany_top_in[19] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput16 chany_bottom_in[9] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_245_ net183 _001_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_6_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk clknet_3_6__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_176_ _115_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input19_I chany_top_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_159_ _114_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_228_ _120_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 mem_bottom_track_1.DFFR_3_.Q net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__248__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_330_ net179 _086_ clknet_3_7__leaf_prog_clk mem_left_track_7.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_261_ net147 _017_ clknet_3_0__leaf_prog_clk mem_top_track_8.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk clknet_3_5__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_192_ _117_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_42_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_1_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_244_ net135 _000_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_7_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_313_ net192 _069_ clknet_3_3__leaf_prog_clk mem_left_track_1.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput28 chany_top_in[1] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput17 chany_top_in[0] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_175_ _115_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_38_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_227_ _120_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_158_ _114_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input31_I chany_top_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold6 mem_top_track_32.DFFR_0_.Q net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_32_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk clknet_3_4__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_260_ net133 _016_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_0_.D vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_191_ _117_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_389_ net20 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_243_ _121_ _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_312_ net151 _068_ clknet_3_3__leaf_prog_clk mem_left_track_1.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput18 chany_top_in[10] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 chany_top_in[2] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_174_ _115_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_226_ _120_ _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_157_ _114_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input24_I chany_top_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold7 mem_bottom_track_1.DFFR_0_.Q net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ _118_ _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_40_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk clknet_3_3__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__271__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_3_5__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_190_ _117_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_388_ net21 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_242_ _121_ _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_311_ net181 _067_ clknet_3_3__leaf_prog_clk mem_left_track_1.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_173_ _115_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput19 chany_top_in[11] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_225_ _120_ _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_156_ _110_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk clknet_3_2__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_35_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input17_I chany_top_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold8 mem_top_track_32.DFFR_1_.Q net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_139_ _112_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_208_ _118_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input9_I chany_bottom_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__261__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_387_ net22 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_310_ net153 _066_ clknet_3_3__leaf_prog_clk mem_left_track_1.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_241_ _121_ _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_172_ _115_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_24_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk clknet_3_1__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_224_ _120_ _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_12_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_155_ _113_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_35_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold9 mem_left_track_3.DFFR_5_.Q net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_40_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_207_ _118_ _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_40_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_138_ _112_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_28_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_8_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_34_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ net24 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk clknet_3_0__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_240_ _121_ _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_17_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_171_ _115_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_24_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_223_ _120_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_37_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_154_ _113_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_20_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_137_ _112_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_206_ _118_ _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_31_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input22_I chany_top_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold90 mem_left_track_23.DFFR_0_.Q net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ net25 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_170_ _115_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_9_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_299_ net131 _055_ clknet_3_2__leaf_prog_clk mem_bottom_track_25.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_153_ _113_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_222_ _110_ _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_136_ _112_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_205_ _118_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_29_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_2__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input15_I chany_bottom_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__264__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input7_I chany_bottom_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__287__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold80 mem_bottom_track_9.DFFR_0_.Q net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold91 mem_left_track_3.DFFR_1_.Q net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_384_ net26 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 chany_top_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__123__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_298_ net189 _054_ clknet_3_2__leaf_prog_clk mem_bottom_track_25.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_1_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_152_ _113_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_20_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_221_ _119_ _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_204_ _118_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_25_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_135_ _112_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold70 mem_left_track_11.DFFR_0_.D net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold81 mem_left_track_5.DFFR_4_.Q net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold92 mem_bottom_track_25.DFFR_2_.Q net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__254__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_383_ net27 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput60 net60 chany_top_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput71 net71 chany_top_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_9_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_297_ net110 _053_ clknet_3_3__leaf_prog_clk mem_bottom_track_25.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_220_ _119_ _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_151_ _113_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__134__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_349_ net129 _105_ clknet_3_5__leaf_prog_clk mem_left_track_17.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_203_ _118_ _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_134_ _110_ _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_2__1__90 chanx_left_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_28_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I chany_top_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold71 mem_top_track_0.DFFR_4_.Q net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold93 mem_left_track_25.DFFR_0_.Q net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold60 mem_left_track_9.DFFR_0_.Q net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold82 mem_left_track_7.DFFR_0_.Q net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_42_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_382_ net23 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput61 net61 chany_top_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput50 net50 chany_bottom_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_296_ net184 _052_ clknet_3_3__leaf_prog_clk mem_bottom_track_25.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__244__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_150_ _113_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__267__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_0_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_348_ net176 _104_ clknet_3_5__leaf_prog_clk mem_left_track_17.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_279_ net152 _035_ clknet_3_4__leaf_prog_clk mem_top_track_32.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_133_ _111_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__145__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_202_ _118_ _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_2__1__80 chany_bottom_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_2__1__91 chanx_left_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_10_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I chany_bottom_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold94 mem_left_track_15.DFFR_0_.Q net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold50 mem_top_track_8.DFFR_3_.Q net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold61 mem_left_track_1.DFFR_3_.Q net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold72 mem_bottom_track_17.DFFR_4_.Q net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold83 mem_bottom_track_33.DFFR_1_.Q net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I chany_bottom_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_381_ net19 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput62 net62 chany_top_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput40 net40 chanx_left_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput51 net51 chany_bottom_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_2_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_295_ net140 _051_ clknet_3_2__leaf_prog_clk mem_bottom_track_17.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_347_ net148 _103_ clknet_3_5__leaf_prog_clk mem_left_track_15.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_278_ net159 _034_ clknet_3_4__leaf_prog_clk mem_bottom_track_1.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_34_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_132_ _111_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_201_ _118_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xsb_2__1__92 chanx_left_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_2__1__81 chany_bottom_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__257__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__156__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold40 mem_bottom_track_25.DFFR_0_.Q net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold51 mem_left_track_13.DFFR_1_.Q net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold73 mem_left_track_29.DFFR_0_.Q net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 mem_top_track_32.DFFR_4_.Q net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold84 mem_left_track_1.DFFR_1_.Q net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold95 mem_bottom_track_33.DFFR_5_.Q net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_380_ net33 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput52 net52 chany_bottom_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput41 net41 chanx_left_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput63 net63 chany_top_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_5_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

