magic
tech gf180mcuD
magscale 1 10
timestamp 1702149425
<< metal1 >>
rect 32274 45166 32286 45218
rect 32338 45215 32350 45218
rect 33394 45215 33406 45218
rect 32338 45169 33406 45215
rect 32338 45166 32350 45169
rect 33394 45166 33406 45169
rect 33458 45166 33470 45218
rect 14130 44830 14142 44882
rect 14194 44879 14206 44882
rect 14914 44879 14926 44882
rect 14194 44833 14926 44879
rect 14194 44830 14206 44833
rect 14914 44830 14926 44833
rect 14978 44830 14990 44882
rect 16818 44830 16830 44882
rect 16882 44879 16894 44882
rect 17490 44879 17502 44882
rect 16882 44833 17502 44879
rect 16882 44830 16894 44833
rect 17490 44830 17502 44833
rect 17554 44830 17566 44882
rect 20178 44830 20190 44882
rect 20242 44879 20254 44882
rect 20962 44879 20974 44882
rect 20242 44833 20974 44879
rect 20242 44830 20254 44833
rect 20962 44830 20974 44833
rect 21026 44830 21038 44882
rect 26898 44830 26910 44882
rect 26962 44879 26974 44882
rect 27570 44879 27582 44882
rect 26962 44833 27582 44879
rect 26962 44830 26974 44833
rect 27570 44830 27582 44833
rect 27634 44830 27646 44882
rect 28914 44830 28926 44882
rect 28978 44879 28990 44882
rect 30034 44879 30046 44882
rect 28978 44833 30046 44879
rect 28978 44830 28990 44833
rect 30034 44830 30046 44833
rect 30098 44830 30110 44882
rect 36978 44830 36990 44882
rect 37042 44879 37054 44882
rect 38098 44879 38110 44882
rect 37042 44833 38110 44879
rect 37042 44830 37054 44833
rect 38098 44830 38110 44833
rect 38162 44830 38174 44882
rect 40338 44830 40350 44882
rect 40402 44879 40414 44882
rect 41906 44879 41918 44882
rect 40402 44833 41918 44879
rect 40402 44830 40414 44833
rect 41906 44830 41918 44833
rect 41970 44830 41982 44882
rect 1344 44714 46592 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 46592 44714
rect 1344 44628 46592 44662
rect 17502 44546 17554 44558
rect 17502 44482 17554 44494
rect 25566 44546 25618 44558
rect 25566 44482 25618 44494
rect 7422 44434 7474 44446
rect 13470 44434 13522 44446
rect 25342 44434 25394 44446
rect 33406 44434 33458 44446
rect 9762 44382 9774 44434
rect 9826 44382 9838 44434
rect 14914 44382 14926 44434
rect 14978 44382 14990 44434
rect 19506 44382 19518 44434
rect 19570 44382 19582 44434
rect 20962 44382 20974 44434
rect 21026 44382 21038 44434
rect 23426 44382 23438 44434
rect 23490 44382 23502 44434
rect 28802 44382 28814 44434
rect 28866 44382 28878 44434
rect 30370 44382 30382 44434
rect 30434 44382 30446 44434
rect 32610 44382 32622 44434
rect 32674 44382 32686 44434
rect 7422 44370 7474 44382
rect 13470 44370 13522 44382
rect 25342 44370 25394 44382
rect 33406 44370 33458 44382
rect 36766 44434 36818 44446
rect 37090 44382 37102 44434
rect 37154 44382 37166 44434
rect 40338 44382 40350 44434
rect 40402 44382 40414 44434
rect 41906 44382 41918 44434
rect 41970 44382 41982 44434
rect 44034 44382 44046 44434
rect 44098 44382 44110 44434
rect 36766 44370 36818 44382
rect 13694 44322 13746 44334
rect 34526 44322 34578 44334
rect 38110 44322 38162 44334
rect 7858 44270 7870 44322
rect 7922 44270 7934 44322
rect 20178 44270 20190 44322
rect 20242 44270 20254 44322
rect 21970 44270 21982 44322
rect 22034 44270 22046 44322
rect 23874 44270 23886 44322
rect 23938 44270 23950 44322
rect 26226 44270 26238 44322
rect 26290 44270 26302 44322
rect 26898 44270 26910 44322
rect 26962 44270 26974 44322
rect 27570 44270 27582 44322
rect 27634 44270 27646 44322
rect 33954 44270 33966 44322
rect 34018 44270 34030 44322
rect 37650 44270 37662 44322
rect 37714 44270 37726 44322
rect 13694 44258 13746 44270
rect 34526 44258 34578 44270
rect 38110 44258 38162 44270
rect 38782 44322 38834 44334
rect 43698 44270 43710 44322
rect 43762 44270 43774 44322
rect 38782 44258 38834 44270
rect 15934 44210 15986 44222
rect 15934 44146 15986 44158
rect 35982 44210 36034 44222
rect 35982 44146 36034 44158
rect 46174 44210 46226 44222
rect 46174 44146 46226 44158
rect 7646 44098 7698 44110
rect 7646 44034 7698 44046
rect 9326 44098 9378 44110
rect 9326 44034 9378 44046
rect 14030 44098 14082 44110
rect 14030 44034 14082 44046
rect 14366 44098 14418 44110
rect 14366 44034 14418 44046
rect 18286 44098 18338 44110
rect 18286 44034 18338 44046
rect 26686 44098 26738 44110
rect 26686 44034 26738 44046
rect 27358 44098 27410 44110
rect 27358 44034 27410 44046
rect 28366 44098 28418 44110
rect 28366 44034 28418 44046
rect 29934 44098 29986 44110
rect 29934 44034 29986 44046
rect 32174 44098 32226 44110
rect 32174 44034 32226 44046
rect 33742 44098 33794 44110
rect 33742 44034 33794 44046
rect 34862 44098 34914 44110
rect 34862 44034 34914 44046
rect 38446 44098 38498 44110
rect 38446 44034 38498 44046
rect 39118 44098 39170 44110
rect 39118 44034 39170 44046
rect 39790 44098 39842 44110
rect 39790 44034 39842 44046
rect 41358 44098 41410 44110
rect 41358 44034 41410 44046
rect 45614 44098 45666 44110
rect 45614 44034 45666 44046
rect 45838 44098 45890 44110
rect 45838 44034 45890 44046
rect 1344 43930 46592 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 46592 43930
rect 1344 43844 46592 43878
rect 17726 43762 17778 43774
rect 17726 43698 17778 43710
rect 27694 43762 27746 43774
rect 27694 43698 27746 43710
rect 30046 43762 30098 43774
rect 30046 43698 30098 43710
rect 34302 43762 34354 43774
rect 34302 43698 34354 43710
rect 37886 43762 37938 43774
rect 37886 43698 37938 43710
rect 18734 43650 18786 43662
rect 18734 43586 18786 43598
rect 19070 43650 19122 43662
rect 19070 43586 19122 43598
rect 20414 43650 20466 43662
rect 20414 43586 20466 43598
rect 21086 43650 21138 43662
rect 21086 43586 21138 43598
rect 21422 43650 21474 43662
rect 21422 43586 21474 43598
rect 21758 43650 21810 43662
rect 21758 43586 21810 43598
rect 23998 43650 24050 43662
rect 23998 43586 24050 43598
rect 25230 43650 25282 43662
rect 25230 43586 25282 43598
rect 25566 43650 25618 43662
rect 25566 43586 25618 43598
rect 30494 43650 30546 43662
rect 30494 43586 30546 43598
rect 31614 43650 31666 43662
rect 31614 43586 31666 43598
rect 31838 43650 31890 43662
rect 31838 43586 31890 43598
rect 34974 43650 35026 43662
rect 34974 43586 35026 43598
rect 35198 43650 35250 43662
rect 35198 43586 35250 43598
rect 35534 43650 35586 43662
rect 35534 43586 35586 43598
rect 38334 43650 38386 43662
rect 38334 43586 38386 43598
rect 39678 43650 39730 43662
rect 39678 43586 39730 43598
rect 39902 43650 39954 43662
rect 39902 43586 39954 43598
rect 40238 43650 40290 43662
rect 40238 43586 40290 43598
rect 42590 43650 42642 43662
rect 42590 43586 42642 43598
rect 42814 43650 42866 43662
rect 42814 43586 42866 43598
rect 18398 43538 18450 43550
rect 19854 43538 19906 43550
rect 19282 43486 19294 43538
rect 19346 43486 19358 43538
rect 18398 43474 18450 43486
rect 19854 43474 19906 43486
rect 20862 43538 20914 43550
rect 20862 43474 20914 43486
rect 22094 43538 22146 43550
rect 22094 43474 22146 43486
rect 22430 43538 22482 43550
rect 22430 43474 22482 43486
rect 23774 43538 23826 43550
rect 23774 43474 23826 43486
rect 24334 43538 24386 43550
rect 24334 43474 24386 43486
rect 26462 43538 26514 43550
rect 26462 43474 26514 43486
rect 28478 43538 28530 43550
rect 28478 43474 28530 43486
rect 29822 43538 29874 43550
rect 41246 43538 41298 43550
rect 30706 43486 30718 43538
rect 30770 43486 30782 43538
rect 32050 43486 32062 43538
rect 32114 43486 32126 43538
rect 38994 43486 39006 43538
rect 39058 43486 39070 43538
rect 43026 43486 43038 43538
rect 43090 43486 43102 43538
rect 45042 43486 45054 43538
rect 45106 43486 45118 43538
rect 29822 43474 29874 43486
rect 41246 43474 41298 43486
rect 22866 43374 22878 43426
rect 22930 43374 22942 43426
rect 26898 43374 26910 43426
rect 26962 43374 26974 43426
rect 28914 43374 28926 43426
rect 28978 43374 28990 43426
rect 41682 43374 41694 43426
rect 41746 43374 41758 43426
rect 46050 43374 46062 43426
rect 46114 43374 46126 43426
rect 1344 43146 46592 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 46592 43146
rect 1344 43060 46592 43094
rect 45726 42978 45778 42990
rect 45726 42914 45778 42926
rect 18174 42866 18226 42878
rect 18174 42802 18226 42814
rect 25006 42866 25058 42878
rect 25006 42802 25058 42814
rect 25566 42754 25618 42766
rect 7522 42702 7534 42754
rect 7586 42702 7598 42754
rect 13906 42702 13918 42754
rect 13970 42702 13982 42754
rect 19058 42702 19070 42754
rect 19122 42702 19134 42754
rect 20626 42702 20638 42754
rect 20690 42702 20702 42754
rect 21634 42702 21646 42754
rect 21698 42702 21710 42754
rect 22418 42702 22430 42754
rect 22482 42702 22494 42754
rect 23314 42702 23326 42754
rect 23378 42702 23390 42754
rect 25566 42690 25618 42702
rect 26574 42754 26626 42766
rect 26574 42690 26626 42702
rect 38222 42754 38274 42766
rect 40238 42754 40290 42766
rect 38994 42702 39006 42754
rect 39058 42702 39070 42754
rect 39666 42702 39678 42754
rect 39730 42702 39742 42754
rect 44034 42702 44046 42754
rect 44098 42702 44110 42754
rect 38222 42690 38274 42702
rect 40238 42690 40290 42702
rect 7758 42642 7810 42654
rect 7758 42578 7810 42590
rect 14142 42642 14194 42654
rect 14142 42578 14194 42590
rect 18846 42642 18898 42654
rect 18846 42578 18898 42590
rect 20414 42642 20466 42654
rect 20414 42578 20466 42590
rect 22206 42642 22258 42654
rect 22206 42578 22258 42590
rect 23550 42642 23602 42654
rect 23550 42578 23602 42590
rect 25902 42642 25954 42654
rect 25902 42578 25954 42590
rect 26238 42642 26290 42654
rect 26238 42578 26290 42590
rect 38558 42642 38610 42654
rect 38558 42578 38610 42590
rect 39230 42642 39282 42654
rect 39230 42578 39282 42590
rect 39902 42642 39954 42654
rect 39902 42578 39954 42590
rect 40574 42642 40626 42654
rect 40574 42578 40626 42590
rect 1710 42530 1762 42542
rect 1710 42466 1762 42478
rect 21870 42530 21922 42542
rect 21870 42466 21922 42478
rect 44270 42530 44322 42542
rect 44270 42466 44322 42478
rect 44942 42530 44994 42542
rect 44942 42466 44994 42478
rect 1344 42362 46592 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 46592 42362
rect 1344 42276 46592 42310
rect 27134 42194 27186 42206
rect 27134 42130 27186 42142
rect 27806 42194 27858 42206
rect 27806 42130 27858 42142
rect 28142 42194 28194 42206
rect 28142 42130 28194 42142
rect 30494 42194 30546 42206
rect 30494 42130 30546 42142
rect 37438 42194 37490 42206
rect 37438 42130 37490 42142
rect 38782 42194 38834 42206
rect 38782 42130 38834 42142
rect 28478 42082 28530 42094
rect 28478 42018 28530 42030
rect 38446 42082 38498 42094
rect 44146 42030 44158 42082
rect 44210 42030 44222 42082
rect 38446 42018 38498 42030
rect 37102 41970 37154 41982
rect 26898 41918 26910 41970
rect 26962 41918 26974 41970
rect 27570 41918 27582 41970
rect 27634 41918 27646 41970
rect 30258 41918 30270 41970
rect 30322 41918 30334 41970
rect 37102 41906 37154 41918
rect 46286 41858 46338 41870
rect 44930 41806 44942 41858
rect 44994 41806 45006 41858
rect 46286 41794 46338 41806
rect 1344 41578 46592 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 46592 41578
rect 1344 41492 46592 41526
rect 44830 41074 44882 41086
rect 44830 41010 44882 41022
rect 45166 41074 45218 41086
rect 45166 41010 45218 41022
rect 45838 41074 45890 41086
rect 45838 41010 45890 41022
rect 46174 41074 46226 41086
rect 46174 41010 46226 41022
rect 1344 40794 46592 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 46592 40794
rect 1344 40708 46592 40742
rect 46062 40626 46114 40638
rect 46062 40562 46114 40574
rect 45378 40462 45390 40514
rect 45442 40462 45454 40514
rect 44146 40238 44158 40290
rect 44210 40238 44222 40290
rect 1344 40010 46592 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 46592 40010
rect 1344 39924 46592 39958
rect 43026 39678 43038 39730
rect 43090 39678 43102 39730
rect 46174 39506 46226 39518
rect 42242 39454 42254 39506
rect 42306 39454 42318 39506
rect 46174 39442 46226 39454
rect 1344 39226 46592 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 46592 39226
rect 1344 39140 46592 39174
rect 43250 38894 43262 38946
rect 43314 38894 43326 38946
rect 45714 38894 45726 38946
rect 45778 38894 45790 38946
rect 41906 38670 41918 38722
rect 41970 38670 41982 38722
rect 44706 38670 44718 38722
rect 44770 38670 44782 38722
rect 1344 38442 46592 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 46592 38442
rect 1344 38356 46592 38390
rect 17826 38110 17838 38162
rect 17890 38110 17902 38162
rect 41346 38110 41358 38162
rect 41410 38110 41422 38162
rect 18834 37886 18846 37938
rect 18898 37886 18910 37938
rect 42354 37886 42366 37938
rect 42418 37886 42430 37938
rect 1344 37658 46592 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 46592 37658
rect 1344 37572 46592 37606
rect 13794 37326 13806 37378
rect 13858 37326 13870 37378
rect 17490 37326 17502 37378
rect 17554 37326 17566 37378
rect 38098 37326 38110 37378
rect 38162 37326 38174 37378
rect 43810 37326 43822 37378
rect 43874 37326 43886 37378
rect 15138 37102 15150 37154
rect 15202 37102 15214 37154
rect 18610 37102 18622 37154
rect 18674 37102 18686 37154
rect 39218 37102 39230 37154
rect 39282 37102 39294 37154
rect 42466 37102 42478 37154
rect 42530 37102 42542 37154
rect 1344 36874 46592 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 46592 36874
rect 1344 36788 46592 36822
rect 14802 36542 14814 36594
rect 14866 36542 14878 36594
rect 18722 36542 18734 36594
rect 18786 36542 18798 36594
rect 22418 36542 22430 36594
rect 22482 36542 22494 36594
rect 38546 36542 38558 36594
rect 38610 36542 38622 36594
rect 40898 36542 40910 36594
rect 40962 36542 40974 36594
rect 15810 36318 15822 36370
rect 15874 36318 15886 36370
rect 19730 36318 19742 36370
rect 19794 36318 19806 36370
rect 23538 36318 23550 36370
rect 23602 36318 23614 36370
rect 37426 36318 37438 36370
rect 37490 36318 37502 36370
rect 41906 36318 41918 36370
rect 41970 36318 41982 36370
rect 1344 36090 46592 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 46592 36090
rect 1344 36004 46592 36038
rect 42466 35870 42478 35922
rect 42530 35870 42542 35922
rect 6178 35758 6190 35810
rect 6242 35758 6254 35810
rect 16034 35758 16046 35810
rect 16098 35758 16110 35810
rect 19506 35758 19518 35810
rect 19570 35758 19582 35810
rect 22642 35758 22654 35810
rect 22706 35758 22718 35810
rect 39890 35758 39902 35810
rect 39954 35758 39966 35810
rect 41694 35698 41746 35710
rect 44930 35646 44942 35698
rect 44994 35646 45006 35698
rect 45378 35646 45390 35698
rect 45442 35646 45454 35698
rect 41694 35634 41746 35646
rect 16830 35586 16882 35598
rect 5170 35534 5182 35586
rect 5234 35534 5246 35586
rect 14690 35534 14702 35586
rect 14754 35534 14766 35586
rect 16482 35534 16494 35586
rect 16546 35534 16558 35586
rect 20626 35534 20638 35586
rect 20690 35534 20702 35586
rect 23650 35534 23662 35586
rect 23714 35534 23726 35586
rect 38882 35534 38894 35586
rect 38946 35534 38958 35586
rect 16830 35522 16882 35534
rect 41806 35474 41858 35486
rect 41806 35410 41858 35422
rect 1344 35306 46592 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 46592 35306
rect 1344 35220 46592 35254
rect 8642 34974 8654 35026
rect 8706 34974 8718 35026
rect 11442 34974 11454 35026
rect 11506 34974 11518 35026
rect 14690 34974 14702 35026
rect 14754 34974 14766 35026
rect 17602 34974 17614 35026
rect 17666 34974 17678 35026
rect 22306 34974 22318 35026
rect 22370 34974 22382 35026
rect 25106 34974 25118 35026
rect 25170 34974 25182 35026
rect 32610 34974 32622 35026
rect 32674 34974 32686 35026
rect 38098 34974 38110 35026
rect 38162 34974 38174 35026
rect 40786 34974 40798 35026
rect 40850 34974 40862 35026
rect 7298 34750 7310 34802
rect 7362 34750 7374 34802
rect 12674 34750 12686 34802
rect 12738 34750 12750 34802
rect 15922 34750 15934 34802
rect 15986 34750 15998 34802
rect 18498 34750 18510 34802
rect 18562 34750 18574 34802
rect 23538 34750 23550 34802
rect 23602 34750 23614 34802
rect 26114 34750 26126 34802
rect 26178 34750 26190 34802
rect 31490 34750 31502 34802
rect 31554 34750 31566 34802
rect 38994 34750 39006 34802
rect 39058 34750 39070 34802
rect 42130 34750 42142 34802
rect 42194 34750 42206 34802
rect 16606 34690 16658 34702
rect 16606 34626 16658 34638
rect 1344 34522 46592 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 46592 34522
rect 1344 34436 46592 34470
rect 1710 34354 1762 34366
rect 45502 34354 45554 34366
rect 2258 34302 2270 34354
rect 2322 34302 2334 34354
rect 44930 34302 44942 34354
rect 44994 34302 45006 34354
rect 1710 34290 1762 34302
rect 45502 34290 45554 34302
rect 8530 34190 8542 34242
rect 8594 34190 8606 34242
rect 13570 34190 13582 34242
rect 13634 34190 13646 34242
rect 15698 34190 15710 34242
rect 15762 34190 15774 34242
rect 19730 34190 19742 34242
rect 19794 34190 19806 34242
rect 21522 34190 21534 34242
rect 21586 34190 21598 34242
rect 27234 34190 27246 34242
rect 27298 34190 27310 34242
rect 30258 34190 30270 34242
rect 30322 34190 30334 34242
rect 33394 34190 33406 34242
rect 33458 34190 33470 34242
rect 37314 34190 37326 34242
rect 37378 34190 37390 34242
rect 5406 34130 5458 34142
rect 4834 34078 4846 34130
rect 4898 34078 4910 34130
rect 5406 34066 5458 34078
rect 41806 34130 41858 34142
rect 42354 34078 42366 34130
rect 42418 34078 42430 34130
rect 41806 34066 41858 34078
rect 5854 34018 5906 34030
rect 11342 34018 11394 34030
rect 7522 33966 7534 34018
rect 7586 33966 7598 34018
rect 5854 33954 5906 33966
rect 11342 33954 11394 33966
rect 12350 34018 12402 34030
rect 17502 34018 17554 34030
rect 12562 33966 12574 34018
rect 12626 33966 12638 34018
rect 14354 33966 14366 34018
rect 14418 33966 14430 34018
rect 12350 33954 12402 33966
rect 17502 33954 17554 33966
rect 17950 34018 18002 34030
rect 30830 34018 30882 34030
rect 40350 34018 40402 34030
rect 18386 33966 18398 34018
rect 18450 33966 18462 34018
rect 22642 33966 22654 34018
rect 22706 33966 22718 34018
rect 26226 33966 26238 34018
rect 26290 33966 26302 34018
rect 29026 33966 29038 34018
rect 29090 33966 29102 34018
rect 31042 33966 31054 34018
rect 31106 33966 31118 34018
rect 34514 33966 34526 34018
rect 34578 33966 34590 34018
rect 38658 33966 38670 34018
rect 38722 33966 38734 34018
rect 17950 33954 18002 33966
rect 30830 33954 30882 33966
rect 40350 33954 40402 33966
rect 41246 34018 41298 34030
rect 41246 33954 41298 33966
rect 41234 33854 41246 33906
rect 41298 33903 41310 33906
rect 41682 33903 41694 33906
rect 41298 33857 41694 33903
rect 41298 33854 41310 33857
rect 41682 33854 41694 33857
rect 41746 33854 41758 33906
rect 1344 33738 46592 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 46592 33738
rect 1344 33652 46592 33686
rect 17054 33570 17106 33582
rect 12338 33518 12350 33570
rect 12402 33567 12414 33570
rect 12898 33567 12910 33570
rect 12402 33521 12910 33567
rect 12402 33518 12414 33521
rect 12898 33518 12910 33521
rect 12962 33518 12974 33570
rect 17054 33506 17106 33518
rect 44382 33570 44434 33582
rect 44382 33506 44434 33518
rect 3602 33406 3614 33458
rect 3666 33406 3678 33458
rect 8866 33406 8878 33458
rect 8930 33406 8942 33458
rect 11890 33406 11902 33458
rect 11954 33406 11966 33458
rect 19506 33406 19518 33458
rect 19570 33406 19582 33458
rect 24658 33406 24670 33458
rect 24722 33406 24734 33458
rect 30146 33406 30158 33458
rect 30210 33406 30222 33458
rect 33170 33406 33182 33458
rect 33234 33406 33246 33458
rect 37986 33406 37998 33458
rect 38050 33406 38062 33458
rect 13358 33346 13410 33358
rect 40686 33346 40738 33358
rect 14018 33294 14030 33346
rect 14082 33294 14094 33346
rect 41346 33294 41358 33346
rect 41410 33294 41422 33346
rect 13358 33282 13410 33294
rect 40686 33282 40738 33294
rect 17726 33234 17778 33246
rect 21646 33234 21698 33246
rect 23326 33234 23378 33246
rect 28254 33234 28306 33246
rect 4946 33182 4958 33234
rect 5010 33182 5022 33234
rect 9650 33182 9662 33234
rect 9714 33182 9726 33234
rect 10882 33182 10894 33234
rect 10946 33182 10958 33234
rect 17378 33182 17390 33234
rect 17442 33182 17454 33234
rect 18386 33182 18398 33234
rect 18450 33182 18462 33234
rect 22978 33182 22990 33234
rect 23042 33182 23054 33234
rect 25666 33182 25678 33234
rect 25730 33182 25742 33234
rect 31154 33182 31166 33234
rect 31218 33182 31230 33234
rect 34066 33182 34078 33234
rect 34130 33182 34142 33234
rect 38994 33182 39006 33234
rect 39058 33182 39070 33234
rect 17726 33170 17778 33182
rect 21646 33170 21698 33182
rect 23326 33170 23378 33182
rect 28254 33170 28306 33182
rect 6190 33122 6242 33134
rect 6190 33058 6242 33070
rect 12350 33122 12402 33134
rect 12350 33058 12402 33070
rect 12910 33122 12962 33134
rect 21534 33122 21586 33134
rect 16482 33070 16494 33122
rect 16546 33070 16558 33122
rect 12910 33058 12962 33070
rect 21534 33058 21586 33070
rect 28366 33122 28418 33134
rect 28366 33058 28418 33070
rect 40014 33122 40066 33134
rect 40014 33058 40066 33070
rect 40462 33122 40514 33134
rect 43586 33070 43598 33122
rect 43650 33070 43662 33122
rect 40462 33058 40514 33070
rect 1344 32954 46592 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 46592 32954
rect 1344 32868 46592 32902
rect 6078 32786 6130 32798
rect 5506 32734 5518 32786
rect 5570 32734 5582 32786
rect 6078 32722 6130 32734
rect 13246 32786 13298 32798
rect 13246 32722 13298 32734
rect 17502 32786 17554 32798
rect 24334 32786 24386 32798
rect 30270 32786 30322 32798
rect 45166 32786 45218 32798
rect 23762 32734 23774 32786
rect 23826 32734 23838 32786
rect 29698 32734 29710 32786
rect 29762 32734 29774 32786
rect 44482 32734 44494 32786
rect 44546 32734 44558 32786
rect 17502 32722 17554 32734
rect 24334 32722 24386 32734
rect 30270 32722 30322 32734
rect 45166 32722 45218 32734
rect 9438 32674 9490 32686
rect 6962 32622 6974 32674
rect 7026 32622 7038 32674
rect 9438 32610 9490 32622
rect 10222 32674 10274 32686
rect 10222 32610 10274 32622
rect 14030 32674 14082 32686
rect 18162 32622 18174 32674
rect 18226 32622 18238 32674
rect 30482 32622 30494 32674
rect 30546 32622 30558 32674
rect 33842 32622 33854 32674
rect 33906 32622 33918 32674
rect 38770 32622 38782 32674
rect 38834 32622 38846 32674
rect 14030 32610 14082 32622
rect 2382 32562 2434 32574
rect 13134 32562 13186 32574
rect 16942 32562 16994 32574
rect 2930 32510 2942 32562
rect 2994 32510 3006 32562
rect 12450 32510 12462 32562
rect 12514 32510 12526 32562
rect 16370 32510 16382 32562
rect 16434 32510 16446 32562
rect 2382 32498 2434 32510
rect 13134 32498 13186 32510
rect 16942 32498 16994 32510
rect 20638 32562 20690 32574
rect 26574 32562 26626 32574
rect 31838 32562 31890 32574
rect 41022 32562 41074 32574
rect 21298 32510 21310 32562
rect 21362 32510 21374 32562
rect 27234 32510 27246 32562
rect 27298 32510 27310 32562
rect 30706 32510 30718 32562
rect 30770 32510 30782 32562
rect 31378 32510 31390 32562
rect 31442 32510 31454 32562
rect 33282 32510 33294 32562
rect 33346 32510 33358 32562
rect 20638 32498 20690 32510
rect 26574 32498 26626 32510
rect 31838 32498 31890 32510
rect 41022 32498 41074 32510
rect 41694 32562 41746 32574
rect 42018 32510 42030 32562
rect 42082 32510 42094 32562
rect 41694 32498 41746 32510
rect 8990 32450 9042 32462
rect 39678 32450 39730 32462
rect 7970 32398 7982 32450
rect 8034 32398 8046 32450
rect 19170 32398 19182 32450
rect 19234 32398 19246 32450
rect 31154 32398 31166 32450
rect 31218 32398 31230 32450
rect 32162 32398 32174 32450
rect 32226 32398 32238 32450
rect 33058 32398 33070 32450
rect 33122 32398 33134 32450
rect 35186 32398 35198 32450
rect 35250 32398 35262 32450
rect 37650 32398 37662 32450
rect 37714 32398 37726 32450
rect 8990 32386 9042 32398
rect 39678 32386 39730 32398
rect 40014 32450 40066 32462
rect 40226 32398 40238 32450
rect 40290 32398 40302 32450
rect 40014 32386 40066 32398
rect 1344 32170 46592 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 46592 32170
rect 1344 32084 46592 32118
rect 17054 32002 17106 32014
rect 17054 31938 17106 31950
rect 5518 31890 5570 31902
rect 3490 31838 3502 31890
rect 3554 31838 3566 31890
rect 5518 31826 5570 31838
rect 13022 31890 13074 31902
rect 13022 31826 13074 31838
rect 20862 31890 20914 31902
rect 20862 31826 20914 31838
rect 21198 31890 21250 31902
rect 21198 31826 21250 31838
rect 28702 31890 28754 31902
rect 28702 31826 28754 31838
rect 29038 31890 29090 31902
rect 35758 31890 35810 31902
rect 33954 31838 33966 31890
rect 34018 31838 34030 31890
rect 29038 31826 29090 31838
rect 35758 31826 35810 31838
rect 42590 31890 42642 31902
rect 42590 31826 42642 31838
rect 9214 31778 9266 31790
rect 8642 31726 8654 31778
rect 8706 31726 8718 31778
rect 9214 31714 9266 31726
rect 9550 31778 9602 31790
rect 13358 31778 13410 31790
rect 17166 31778 17218 31790
rect 25230 31778 25282 31790
rect 32510 31778 32562 31790
rect 9986 31726 9998 31778
rect 10050 31726 10062 31778
rect 13906 31726 13918 31778
rect 13970 31726 13982 31778
rect 17826 31726 17838 31778
rect 17890 31726 17902 31778
rect 24210 31726 24222 31778
rect 24274 31726 24286 31778
rect 24770 31726 24782 31778
rect 24834 31726 24846 31778
rect 25666 31726 25678 31778
rect 25730 31726 25742 31778
rect 32050 31726 32062 31778
rect 32114 31726 32126 31778
rect 9550 31714 9602 31726
rect 13358 31714 13410 31726
rect 17166 31714 17218 31726
rect 25230 31714 25282 31726
rect 32510 31714 32562 31726
rect 39118 31778 39170 31790
rect 39442 31726 39454 31778
rect 39506 31726 39518 31778
rect 43026 31726 43038 31778
rect 43090 31726 43102 31778
rect 39118 31714 39170 31726
rect 21982 31666 22034 31678
rect 2370 31614 2382 31666
rect 2434 31614 2446 31666
rect 21982 31602 22034 31614
rect 29822 31666 29874 31678
rect 43710 31666 43762 31678
rect 34962 31614 34974 31666
rect 35026 31614 35038 31666
rect 42802 31614 42814 31666
rect 42866 31614 42878 31666
rect 29822 31602 29874 31614
rect 43710 31602 43762 31614
rect 35870 31554 35922 31566
rect 6066 31502 6078 31554
rect 6130 31502 6142 31554
rect 12338 31502 12350 31554
rect 12402 31502 12414 31554
rect 16482 31502 16494 31554
rect 16546 31502 16558 31554
rect 20290 31502 20302 31554
rect 20354 31502 20366 31554
rect 28130 31502 28142 31554
rect 28194 31502 28206 31554
rect 35870 31490 35922 31502
rect 37102 31554 37154 31566
rect 37102 31490 37154 31502
rect 38782 31554 38834 31566
rect 43822 31554 43874 31566
rect 42018 31502 42030 31554
rect 42082 31502 42094 31554
rect 38782 31490 38834 31502
rect 43822 31490 43874 31502
rect 44942 31554 44994 31566
rect 44942 31490 44994 31502
rect 1344 31386 46592 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 46592 31386
rect 1344 31300 46592 31334
rect 5742 31218 5794 31230
rect 5742 31154 5794 31166
rect 15710 31218 15762 31230
rect 15710 31154 15762 31166
rect 17278 31218 17330 31230
rect 24782 31218 24834 31230
rect 30046 31218 30098 31230
rect 36654 31218 36706 31230
rect 44606 31218 44658 31230
rect 18050 31166 18062 31218
rect 18114 31166 18126 31218
rect 24210 31166 24222 31218
rect 24274 31166 24286 31218
rect 28914 31166 28926 31218
rect 28978 31166 28990 31218
rect 35858 31166 35870 31218
rect 35922 31166 35934 31218
rect 43810 31166 43822 31218
rect 43874 31166 43886 31218
rect 17278 31154 17330 31166
rect 24782 31154 24834 31166
rect 30046 31154 30098 31166
rect 36654 31154 36706 31166
rect 44606 31154 44658 31166
rect 4958 31106 5010 31118
rect 14926 31106 14978 31118
rect 29710 31106 29762 31118
rect 39678 31106 39730 31118
rect 8530 31054 8542 31106
rect 8594 31054 8606 31106
rect 10770 31054 10782 31106
rect 10834 31054 10846 31106
rect 25218 31054 25230 31106
rect 25282 31054 25294 31106
rect 31938 31054 31950 31106
rect 32002 31054 32014 31106
rect 38882 31054 38894 31106
rect 38946 31054 38958 31106
rect 4958 31042 5010 31054
rect 14926 31042 14978 31054
rect 29710 31042 29762 31054
rect 39678 31042 39730 31054
rect 2270 30994 2322 31006
rect 6078 30994 6130 31006
rect 2706 30942 2718 30994
rect 2770 30942 2782 30994
rect 2270 30930 2322 30942
rect 6078 30930 6130 30942
rect 9998 30994 10050 31006
rect 20750 30994 20802 31006
rect 10994 30942 11006 30994
rect 11058 30942 11070 30994
rect 12114 30942 12126 30994
rect 12178 30942 12190 30994
rect 12562 30942 12574 30994
rect 12626 30942 12638 30994
rect 20290 30942 20302 30994
rect 20354 30942 20366 30994
rect 9998 30930 10050 30942
rect 20750 30930 20802 30942
rect 21086 30994 21138 31006
rect 26014 30994 26066 31006
rect 41134 30994 41186 31006
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 26674 30942 26686 30994
rect 26738 30942 26750 30994
rect 33058 30942 33070 30994
rect 33122 30942 33134 30994
rect 33618 30942 33630 30994
rect 33682 30942 33694 30994
rect 41570 30942 41582 30994
rect 41634 30942 41646 30994
rect 45042 30942 45054 30994
rect 45106 30942 45118 30994
rect 21086 30930 21138 30942
rect 26014 30930 26066 30942
rect 41134 30930 41186 30942
rect 7198 30882 7250 30894
rect 10446 30882 10498 30894
rect 7522 30830 7534 30882
rect 7586 30830 7598 30882
rect 7198 30818 7250 30830
rect 10446 30818 10498 30830
rect 11454 30882 11506 30894
rect 16158 30882 16210 30894
rect 16830 30882 16882 30894
rect 11666 30830 11678 30882
rect 11730 30830 11742 30882
rect 16482 30830 16494 30882
rect 16546 30830 16558 30882
rect 11454 30818 11506 30830
rect 16158 30818 16210 30830
rect 16830 30818 16882 30830
rect 25566 30882 25618 30894
rect 36990 30882 37042 30894
rect 30930 30830 30942 30882
rect 30994 30830 31006 30882
rect 25566 30818 25618 30830
rect 36990 30818 37042 30830
rect 37438 30882 37490 30894
rect 45614 30882 45666 30894
rect 37874 30830 37886 30882
rect 37938 30830 37950 30882
rect 39890 30830 39902 30882
rect 39954 30830 39966 30882
rect 44818 30830 44830 30882
rect 44882 30830 44894 30882
rect 37438 30818 37490 30830
rect 45614 30818 45666 30830
rect 1344 30602 46592 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 46592 30602
rect 1344 30516 46592 30550
rect 4050 30270 4062 30322
rect 4114 30270 4126 30322
rect 14914 30270 14926 30322
rect 14978 30270 14990 30322
rect 26898 30270 26910 30322
rect 26962 30270 26974 30322
rect 42130 30270 42142 30322
rect 42194 30270 42206 30322
rect 45714 30270 45726 30322
rect 45778 30270 45790 30322
rect 9214 30210 9266 30222
rect 5618 30158 5630 30210
rect 5682 30158 5694 30210
rect 6066 30158 6078 30210
rect 6130 30158 6142 30210
rect 9214 30146 9266 30158
rect 9550 30210 9602 30222
rect 13022 30210 13074 30222
rect 15598 30210 15650 30222
rect 19070 30210 19122 30222
rect 25678 30210 25730 30222
rect 9874 30158 9886 30210
rect 9938 30158 9950 30210
rect 13682 30158 13694 30210
rect 13746 30158 13758 30210
rect 14242 30158 14254 30210
rect 14306 30158 14318 30210
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 20402 30158 20414 30210
rect 20466 30158 20478 30210
rect 21522 30158 21534 30210
rect 21586 30158 21598 30210
rect 25106 30158 25118 30210
rect 25170 30158 25182 30210
rect 9550 30146 9602 30158
rect 13022 30146 13074 30158
rect 15598 30146 15650 30158
rect 19070 30146 19122 30158
rect 25678 30146 25730 30158
rect 29262 30210 29314 30222
rect 32734 30210 32786 30222
rect 29698 30158 29710 30210
rect 29762 30158 29774 30210
rect 29262 30146 29314 30158
rect 32734 30146 32786 30158
rect 32846 30210 32898 30222
rect 36542 30210 36594 30222
rect 40910 30210 40962 30222
rect 35970 30158 35982 30210
rect 36034 30158 36046 30210
rect 37314 30158 37326 30210
rect 37378 30158 37390 30210
rect 37762 30158 37774 30210
rect 37826 30158 37838 30210
rect 32846 30146 32898 30158
rect 36542 30146 36594 30158
rect 40910 30146 40962 30158
rect 41694 30210 41746 30222
rect 41694 30146 41746 30158
rect 44270 30210 44322 30222
rect 45042 30158 45054 30210
rect 45106 30158 45118 30210
rect 44270 30146 44322 30158
rect 1934 30098 1986 30110
rect 14590 30098 14642 30110
rect 3042 30046 3054 30098
rect 3106 30046 3118 30098
rect 13458 30046 13470 30098
rect 13522 30046 13534 30098
rect 1934 30034 1986 30046
rect 14590 30034 14642 30046
rect 15262 30098 15314 30110
rect 15262 30034 15314 30046
rect 16382 30098 16434 30110
rect 16382 30034 16434 30046
rect 20750 30098 20802 30110
rect 45502 30098 45554 30110
rect 21746 30046 21758 30098
rect 21810 30046 21822 30098
rect 27906 30046 27918 30098
rect 27970 30046 27982 30098
rect 43138 30046 43150 30098
rect 43202 30046 43214 30098
rect 43922 30046 43934 30098
rect 43986 30046 43998 30098
rect 44818 30046 44830 30098
rect 44882 30046 44894 30098
rect 20750 30034 20802 30046
rect 45502 30034 45554 30046
rect 2046 29986 2098 29998
rect 21982 29986 22034 29998
rect 41246 29986 41298 29998
rect 8642 29934 8654 29986
rect 8706 29934 8718 29986
rect 12450 29934 12462 29986
rect 12514 29934 12526 29986
rect 22754 29934 22766 29986
rect 22818 29934 22830 29986
rect 32162 29934 32174 29986
rect 32226 29934 32238 29986
rect 33506 29934 33518 29986
rect 33570 29934 33582 29986
rect 40226 29934 40238 29986
rect 40290 29934 40302 29986
rect 2046 29922 2098 29934
rect 21982 29922 22034 29934
rect 41246 29922 41298 29934
rect 1344 29818 46592 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 46592 29818
rect 1344 29732 46592 29766
rect 8206 29650 8258 29662
rect 7522 29598 7534 29650
rect 7586 29598 7598 29650
rect 8206 29586 8258 29598
rect 8654 29650 8706 29662
rect 13134 29650 13186 29662
rect 16942 29650 16994 29662
rect 12338 29598 12350 29650
rect 12402 29598 12414 29650
rect 16370 29598 16382 29650
rect 16434 29598 16446 29650
rect 8654 29586 8706 29598
rect 13134 29586 13186 29598
rect 16942 29586 16994 29598
rect 21982 29650 22034 29662
rect 21982 29586 22034 29598
rect 26014 29650 26066 29662
rect 31502 29650 31554 29662
rect 30930 29598 30942 29650
rect 30994 29598 31006 29650
rect 26014 29586 26066 29598
rect 31502 29586 31554 29598
rect 38782 29650 38834 29662
rect 38782 29586 38834 29598
rect 40798 29650 40850 29662
rect 44942 29650 44994 29662
rect 41570 29598 41582 29650
rect 41634 29598 41646 29650
rect 40798 29586 40850 29598
rect 44942 29586 44994 29598
rect 21198 29538 21250 29550
rect 27582 29538 27634 29550
rect 2258 29486 2270 29538
rect 2322 29486 2334 29538
rect 17378 29486 17390 29538
rect 17442 29486 17454 29538
rect 22642 29486 22654 29538
rect 22706 29486 22718 29538
rect 25218 29486 25230 29538
rect 25282 29486 25294 29538
rect 21198 29474 21250 29486
rect 27582 29474 27634 29486
rect 32062 29538 32114 29550
rect 32062 29474 32114 29486
rect 33182 29538 33234 29550
rect 37998 29538 38050 29550
rect 33506 29486 33518 29538
rect 33570 29486 33582 29538
rect 45826 29486 45838 29538
rect 45890 29486 45902 29538
rect 33182 29474 33234 29486
rect 37998 29474 38050 29486
rect 4734 29426 4786 29438
rect 9662 29426 9714 29438
rect 25902 29426 25954 29438
rect 35310 29426 35362 29438
rect 5058 29374 5070 29426
rect 5122 29374 5134 29426
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 13346 29374 13358 29426
rect 13410 29374 13422 29426
rect 13906 29374 13918 29426
rect 13970 29374 13982 29426
rect 17602 29374 17614 29426
rect 17666 29374 17678 29426
rect 18386 29374 18398 29426
rect 18450 29374 18462 29426
rect 18834 29374 18846 29426
rect 18898 29374 18910 29426
rect 25442 29374 25454 29426
rect 25506 29374 25518 29426
rect 27906 29374 27918 29426
rect 27970 29374 27982 29426
rect 28466 29374 28478 29426
rect 28530 29374 28542 29426
rect 35746 29374 35758 29426
rect 35810 29374 35822 29426
rect 39106 29374 39118 29426
rect 39170 29374 39182 29426
rect 43810 29374 43822 29426
rect 43874 29374 43886 29426
rect 44370 29374 44382 29426
rect 44434 29374 44446 29426
rect 4734 29362 4786 29374
rect 9662 29362 9714 29374
rect 25902 29362 25954 29374
rect 35310 29362 35362 29374
rect 8766 29314 8818 29326
rect 27022 29314 27074 29326
rect 40014 29314 40066 29326
rect 3266 29262 3278 29314
rect 3330 29262 3342 29314
rect 23650 29262 23662 29314
rect 23714 29262 23726 29314
rect 27346 29262 27358 29314
rect 27410 29262 27422 29314
rect 31714 29262 31726 29314
rect 31778 29262 31790 29314
rect 8766 29250 8818 29262
rect 27022 29250 27074 29262
rect 40014 29250 40066 29262
rect 45054 29314 45106 29326
rect 45054 29250 45106 29262
rect 45502 29314 45554 29326
rect 45502 29250 45554 29262
rect 1344 29034 46592 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 46592 29034
rect 1344 28948 46592 28982
rect 11790 28866 11842 28878
rect 11790 28802 11842 28814
rect 18846 28866 18898 28878
rect 18846 28802 18898 28814
rect 29038 28866 29090 28878
rect 29038 28802 29090 28814
rect 36542 28866 36594 28878
rect 36542 28802 36594 28814
rect 40574 28866 40626 28878
rect 44930 28814 44942 28866
rect 44994 28863 45006 28866
rect 45378 28863 45390 28866
rect 44994 28817 45390 28863
rect 44994 28814 45006 28817
rect 45378 28814 45390 28817
rect 45442 28814 45454 28866
rect 40574 28802 40626 28814
rect 1934 28754 1986 28766
rect 14030 28754 14082 28766
rect 2146 28702 2158 28754
rect 2210 28702 2222 28754
rect 4050 28702 4062 28754
rect 4114 28702 4126 28754
rect 5618 28702 5630 28754
rect 5682 28702 5694 28754
rect 7522 28702 7534 28754
rect 7586 28702 7598 28754
rect 1934 28690 1986 28702
rect 14030 28690 14082 28702
rect 14478 28754 14530 28766
rect 44942 28754 44994 28766
rect 19058 28702 19070 28754
rect 19122 28702 19134 28754
rect 21634 28702 21646 28754
rect 21698 28702 21710 28754
rect 24210 28702 24222 28754
rect 24274 28702 24286 28754
rect 28130 28702 28142 28754
rect 28194 28702 28206 28754
rect 14478 28690 14530 28702
rect 44942 28690 44994 28702
rect 45390 28754 45442 28766
rect 45390 28690 45442 28702
rect 6638 28642 6690 28654
rect 8318 28642 8370 28654
rect 12910 28642 12962 28654
rect 6290 28590 6302 28642
rect 6354 28590 6366 28642
rect 7410 28590 7422 28642
rect 7474 28590 7486 28642
rect 8754 28590 8766 28642
rect 8818 28590 8830 28642
rect 12002 28590 12014 28642
rect 12066 28590 12078 28642
rect 12226 28590 12238 28642
rect 12290 28590 12302 28642
rect 6638 28578 6690 28590
rect 8318 28578 8370 28590
rect 12910 28578 12962 28590
rect 13582 28642 13634 28654
rect 13582 28578 13634 28590
rect 14926 28642 14978 28654
rect 14926 28578 14978 28590
rect 15150 28642 15202 28654
rect 20750 28642 20802 28654
rect 25006 28642 25058 28654
rect 32510 28642 32562 28654
rect 15810 28590 15822 28642
rect 15874 28590 15886 28642
rect 19282 28590 19294 28642
rect 19346 28590 19358 28642
rect 23762 28590 23774 28642
rect 23826 28590 23838 28642
rect 24434 28590 24446 28642
rect 24498 28590 24510 28642
rect 26562 28590 26574 28642
rect 26626 28590 26638 28642
rect 32162 28590 32174 28642
rect 32226 28590 32238 28642
rect 15150 28578 15202 28590
rect 20750 28578 20802 28590
rect 25006 28578 25058 28590
rect 32510 28578 32562 28590
rect 32846 28642 32898 28654
rect 33394 28590 33406 28642
rect 33458 28590 33470 28642
rect 36978 28590 36990 28642
rect 37042 28590 37054 28642
rect 37538 28590 37550 28642
rect 37602 28590 37614 28642
rect 40786 28590 40798 28642
rect 40850 28590 40862 28642
rect 41346 28590 41358 28642
rect 41410 28590 41422 28642
rect 32846 28578 32898 28590
rect 5966 28530 6018 28542
rect 3042 28478 3054 28530
rect 3106 28478 3118 28530
rect 5966 28466 6018 28478
rect 29822 28530 29874 28542
rect 29822 28466 29874 28478
rect 44382 28418 44434 28430
rect 11218 28366 11230 28418
rect 11282 28366 11294 28418
rect 18050 28366 18062 28418
rect 18114 28366 18126 28418
rect 35970 28366 35982 28418
rect 36034 28366 36046 28418
rect 39890 28366 39902 28418
rect 39954 28366 39966 28418
rect 43586 28366 43598 28418
rect 43650 28366 43662 28418
rect 44382 28354 44434 28366
rect 1344 28250 46592 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 46592 28250
rect 1344 28164 46592 28198
rect 3502 28082 3554 28094
rect 8318 28082 8370 28094
rect 16942 28082 16994 28094
rect 4274 28030 4286 28082
rect 4338 28030 4350 28082
rect 16370 28030 16382 28082
rect 16434 28030 16446 28082
rect 3502 28018 3554 28030
rect 8318 28018 8370 28030
rect 16942 28018 16994 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 20750 28082 20802 28094
rect 30606 28082 30658 28094
rect 21522 28030 21534 28082
rect 21586 28030 21598 28082
rect 29810 28030 29822 28082
rect 29874 28030 29886 28082
rect 20750 28018 20802 28030
rect 30606 28018 30658 28030
rect 31502 28082 31554 28094
rect 31502 28018 31554 28030
rect 37326 28082 37378 28094
rect 44594 28030 44606 28082
rect 44658 28030 44670 28082
rect 37326 28018 37378 28030
rect 3278 27970 3330 27982
rect 3278 27906 3330 27918
rect 36542 27970 36594 27982
rect 41246 27970 41298 27982
rect 40898 27918 40910 27970
rect 40962 27918 40974 27970
rect 45826 27918 45838 27970
rect 45890 27918 45902 27970
rect 36542 27906 36594 27918
rect 41246 27906 41298 27918
rect 7198 27858 7250 27870
rect 24446 27858 24498 27870
rect 27134 27858 27186 27870
rect 33854 27858 33906 27870
rect 41470 27858 41522 27870
rect 6514 27806 6526 27858
rect 6578 27806 6590 27858
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 13346 27806 13358 27858
rect 13410 27806 13422 27858
rect 13906 27806 13918 27858
rect 13970 27806 13982 27858
rect 18274 27806 18286 27858
rect 18338 27806 18350 27858
rect 23874 27806 23886 27858
rect 23938 27806 23950 27858
rect 25442 27806 25454 27858
rect 25506 27806 25518 27858
rect 27458 27806 27470 27858
rect 27522 27806 27534 27858
rect 31826 27806 31838 27858
rect 31890 27806 31902 27858
rect 34290 27806 34302 27858
rect 34354 27806 34366 27858
rect 37538 27806 37550 27858
rect 37602 27806 37614 27858
rect 42130 27806 42142 27858
rect 42194 27806 42206 27858
rect 46050 27806 46062 27858
rect 46114 27806 46126 27858
rect 7198 27794 7250 27806
rect 24446 27794 24498 27806
rect 27134 27794 27186 27806
rect 33854 27794 33906 27806
rect 41470 27794 41522 27806
rect 9886 27746 9938 27758
rect 45614 27746 45666 27758
rect 2930 27694 2942 27746
rect 2994 27694 3006 27746
rect 11778 27694 11790 27746
rect 11842 27694 11854 27746
rect 19058 27694 19070 27746
rect 19122 27694 19134 27746
rect 25218 27694 25230 27746
rect 25282 27694 25294 27746
rect 38658 27694 38670 27746
rect 38722 27694 38734 27746
rect 9886 27682 9938 27694
rect 45614 27682 45666 27694
rect 45166 27634 45218 27646
rect 45166 27570 45218 27582
rect 1344 27466 46592 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 46592 27466
rect 1344 27380 46592 27414
rect 16270 27298 16322 27310
rect 16270 27234 16322 27246
rect 24894 27298 24946 27310
rect 24894 27234 24946 27246
rect 25006 27298 25058 27310
rect 25006 27234 25058 27246
rect 40574 27298 40626 27310
rect 40574 27234 40626 27246
rect 44382 27298 44434 27310
rect 44382 27234 44434 27246
rect 5966 27186 6018 27198
rect 4050 27134 4062 27186
rect 4114 27134 4126 27186
rect 5618 27134 5630 27186
rect 5682 27134 5694 27186
rect 5966 27122 6018 27134
rect 12126 27186 12178 27198
rect 20526 27186 20578 27198
rect 46174 27186 46226 27198
rect 14914 27134 14926 27186
rect 14978 27134 14990 27186
rect 20290 27134 20302 27186
rect 20354 27134 20366 27186
rect 34514 27134 34526 27186
rect 34578 27134 34590 27186
rect 12126 27122 12178 27134
rect 20526 27122 20578 27134
rect 46174 27122 46226 27134
rect 7982 27074 8034 27086
rect 19742 27074 19794 27086
rect 6962 27022 6974 27074
rect 7026 27022 7038 27074
rect 8530 27022 8542 27074
rect 8594 27022 8606 27074
rect 13458 27022 13470 27074
rect 13522 27022 13534 27074
rect 19394 27022 19406 27074
rect 19458 27022 19470 27074
rect 7982 27010 8034 27022
rect 19742 27010 19794 27022
rect 21198 27074 21250 27086
rect 28702 27074 28754 27086
rect 40686 27074 40738 27086
rect 44942 27074 44994 27086
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 28130 27022 28142 27074
rect 28194 27022 28206 27074
rect 30146 27022 30158 27074
rect 30210 27022 30222 27074
rect 31826 27022 31838 27074
rect 31890 27022 31902 27074
rect 36978 27022 36990 27074
rect 37042 27022 37054 27074
rect 37426 27022 37438 27074
rect 37490 27022 37502 27074
rect 41346 27022 41358 27074
rect 41410 27022 41422 27074
rect 21198 27010 21250 27022
rect 28702 27010 28754 27022
rect 40686 27010 40738 27022
rect 44942 27010 44994 27022
rect 6414 26962 6466 26974
rect 11678 26962 11730 26974
rect 12910 26962 12962 26974
rect 3042 26910 3054 26962
rect 3106 26910 3118 26962
rect 6738 26910 6750 26962
rect 6802 26910 6814 26962
rect 12562 26910 12574 26962
rect 12626 26910 12638 26962
rect 6414 26898 6466 26910
rect 11678 26898 11730 26910
rect 12910 26898 12962 26910
rect 24110 26962 24162 26974
rect 36430 26962 36482 26974
rect 35522 26910 35534 26962
rect 35586 26910 35598 26962
rect 24110 26898 24162 26910
rect 36430 26898 36482 26910
rect 39790 26962 39842 26974
rect 39790 26898 39842 26910
rect 45726 26962 45778 26974
rect 45726 26898 45778 26910
rect 11106 26798 11118 26850
rect 11170 26798 11182 26850
rect 17042 26798 17054 26850
rect 17106 26798 17118 26850
rect 25778 26798 25790 26850
rect 25842 26798 25854 26850
rect 43810 26798 43822 26850
rect 43874 26798 43886 26850
rect 1344 26682 46592 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 46592 26682
rect 1344 26596 46592 26630
rect 1598 26514 1650 26526
rect 9102 26514 9154 26526
rect 2370 26462 2382 26514
rect 2434 26462 2446 26514
rect 8530 26462 8542 26514
rect 8594 26462 8606 26514
rect 1598 26450 1650 26462
rect 9102 26450 9154 26462
rect 9662 26514 9714 26526
rect 17502 26514 17554 26526
rect 14914 26462 14926 26514
rect 14978 26462 14990 26514
rect 9662 26450 9714 26462
rect 17502 26450 17554 26462
rect 18062 26514 18114 26526
rect 23214 26514 23266 26526
rect 32958 26514 33010 26526
rect 22418 26462 22430 26514
rect 22482 26462 22494 26514
rect 28242 26462 28254 26514
rect 28306 26462 28318 26514
rect 18062 26450 18114 26462
rect 23214 26450 23266 26462
rect 32958 26450 33010 26462
rect 36766 26514 36818 26526
rect 43810 26462 43822 26514
rect 43874 26462 43886 26514
rect 36766 26450 36818 26462
rect 33742 26402 33794 26414
rect 11218 26350 11230 26402
rect 11282 26350 11294 26402
rect 16482 26350 16494 26402
rect 16546 26350 16558 26402
rect 18834 26350 18846 26402
rect 18898 26350 18910 26402
rect 33742 26338 33794 26350
rect 37550 26402 37602 26414
rect 45378 26350 45390 26402
rect 45442 26350 45454 26402
rect 37550 26338 37602 26350
rect 5630 26290 5682 26302
rect 11790 26290 11842 26302
rect 25118 26290 25170 26302
rect 36654 26290 36706 26302
rect 40462 26290 40514 26302
rect 4722 26238 4734 26290
rect 4786 26238 4798 26290
rect 5170 26238 5182 26290
rect 5234 26238 5246 26290
rect 6066 26238 6078 26290
rect 6130 26238 6142 26290
rect 12338 26238 12350 26290
rect 12402 26238 12414 26290
rect 19058 26238 19070 26290
rect 19122 26238 19134 26290
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 23874 26238 23886 26290
rect 23938 26238 23950 26290
rect 25666 26238 25678 26290
rect 25730 26238 25742 26290
rect 29026 26238 29038 26290
rect 29090 26238 29102 26290
rect 36082 26238 36094 26290
rect 36146 26238 36158 26290
rect 39890 26238 39902 26290
rect 39954 26238 39966 26290
rect 5630 26226 5682 26238
rect 11790 26226 11842 26238
rect 25118 26226 25170 26238
rect 36654 26226 36706 26238
rect 40462 26226 40514 26238
rect 41022 26290 41074 26302
rect 46174 26290 46226 26302
rect 41458 26238 41470 26290
rect 41522 26238 41534 26290
rect 41022 26226 41074 26238
rect 46174 26226 46226 26238
rect 9550 26178 9602 26190
rect 9550 26114 9602 26126
rect 11566 26178 11618 26190
rect 11566 26114 11618 26126
rect 15822 26178 15874 26190
rect 16830 26178 16882 26190
rect 16034 26126 16046 26178
rect 16098 26126 16110 26178
rect 15822 26114 15874 26126
rect 16830 26114 16882 26126
rect 17950 26178 18002 26190
rect 45054 26178 45106 26190
rect 23986 26126 23998 26178
rect 24050 26126 24062 26178
rect 31378 26126 31390 26178
rect 31442 26126 31454 26178
rect 44706 26126 44718 26178
rect 44770 26126 44782 26178
rect 17950 26114 18002 26126
rect 45054 26114 45106 26126
rect 45726 26178 45778 26190
rect 45726 26114 45778 26126
rect 15486 26066 15538 26078
rect 15486 26002 15538 26014
rect 28814 26066 28866 26078
rect 28814 26002 28866 26014
rect 44494 26066 44546 26078
rect 44494 26002 44546 26014
rect 1344 25898 46592 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 46592 25898
rect 1344 25812 46592 25846
rect 13022 25730 13074 25742
rect 13022 25666 13074 25678
rect 35310 25730 35362 25742
rect 35310 25666 35362 25678
rect 45502 25618 45554 25630
rect 4050 25566 4062 25618
rect 4114 25566 4126 25618
rect 6962 25566 6974 25618
rect 7026 25566 7038 25618
rect 16370 25566 16382 25618
rect 16434 25566 16446 25618
rect 18946 25566 18958 25618
rect 19010 25566 19022 25618
rect 23090 25566 23102 25618
rect 23154 25566 23166 25618
rect 28242 25566 28254 25618
rect 28306 25566 28318 25618
rect 37986 25566 37998 25618
rect 38050 25566 38062 25618
rect 43810 25566 43822 25618
rect 43874 25566 43886 25618
rect 44818 25566 44830 25618
rect 44882 25566 44894 25618
rect 45502 25554 45554 25566
rect 9550 25506 9602 25518
rect 24558 25506 24610 25518
rect 31614 25506 31666 25518
rect 8530 25454 8542 25506
rect 8594 25454 8606 25506
rect 9874 25454 9886 25506
rect 9938 25454 9950 25506
rect 13682 25454 13694 25506
rect 13746 25454 13758 25506
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 20290 25454 20302 25506
rect 20354 25454 20366 25506
rect 24994 25454 25006 25506
rect 25058 25454 25070 25506
rect 31042 25454 31054 25506
rect 31106 25454 31118 25506
rect 32274 25454 32286 25506
rect 32338 25454 32350 25506
rect 37762 25454 37774 25506
rect 37826 25454 37838 25506
rect 38434 25454 38446 25506
rect 38498 25454 38510 25506
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 43138 25454 43150 25506
rect 43202 25454 43214 25506
rect 9550 25442 9602 25454
rect 24558 25442 24610 25454
rect 31614 25442 31666 25454
rect 28590 25394 28642 25406
rect 35870 25394 35922 25406
rect 3042 25342 3054 25394
rect 3106 25342 3118 25394
rect 13458 25342 13470 25394
rect 13522 25342 13534 25394
rect 14130 25342 14142 25394
rect 14194 25342 14206 25394
rect 15362 25342 15374 25394
rect 15426 25342 15438 25394
rect 22082 25342 22094 25394
rect 22146 25342 22158 25394
rect 29586 25342 29598 25394
rect 29650 25342 29662 25394
rect 30370 25342 30382 25394
rect 30434 25342 30446 25394
rect 30818 25342 30830 25394
rect 30882 25342 30894 25394
rect 28590 25330 28642 25342
rect 35870 25330 35922 25342
rect 37326 25394 37378 25406
rect 37326 25330 37378 25342
rect 42254 25394 42306 25406
rect 43598 25394 43650 25406
rect 42914 25342 42926 25394
rect 42978 25342 42990 25394
rect 42254 25330 42306 25342
rect 43598 25330 43650 25342
rect 45166 25394 45218 25406
rect 45166 25330 45218 25342
rect 8990 25282 9042 25294
rect 20750 25282 20802 25294
rect 28030 25282 28082 25294
rect 35758 25282 35810 25294
rect 12450 25230 12462 25282
rect 12514 25230 12526 25282
rect 27234 25230 27246 25282
rect 27298 25230 27310 25282
rect 34738 25230 34750 25282
rect 34802 25230 34814 25282
rect 8990 25218 9042 25230
rect 20750 25218 20802 25230
rect 28030 25218 28082 25230
rect 35758 25218 35810 25230
rect 37214 25282 37266 25294
rect 42030 25282 42082 25294
rect 41458 25230 41470 25282
rect 41522 25230 41534 25282
rect 37214 25218 37266 25230
rect 42030 25218 42082 25230
rect 42366 25282 42418 25294
rect 42366 25218 42418 25230
rect 45614 25282 45666 25294
rect 45614 25218 45666 25230
rect 1344 25114 46592 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 46592 25114
rect 1344 25028 46592 25062
rect 3950 24946 4002 24958
rect 20974 24946 21026 24958
rect 24782 24946 24834 24958
rect 4722 24894 4734 24946
rect 4786 24894 4798 24946
rect 12562 24894 12574 24946
rect 12626 24894 12638 24946
rect 16146 24894 16158 24946
rect 16210 24894 16222 24946
rect 20402 24894 20414 24946
rect 20466 24894 20478 24946
rect 23986 24894 23998 24946
rect 24050 24894 24062 24946
rect 3950 24882 4002 24894
rect 20974 24882 21026 24894
rect 24782 24882 24834 24894
rect 29374 24946 29426 24958
rect 45054 24946 45106 24958
rect 35970 24894 35982 24946
rect 36034 24894 36046 24946
rect 44482 24894 44494 24946
rect 44546 24894 44558 24946
rect 29374 24882 29426 24894
rect 45054 24882 45106 24894
rect 2046 24834 2098 24846
rect 2046 24770 2098 24782
rect 28590 24834 28642 24846
rect 28590 24770 28642 24782
rect 41022 24834 41074 24846
rect 41022 24770 41074 24782
rect 45502 24834 45554 24846
rect 45502 24770 45554 24782
rect 7646 24722 7698 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 3490 24670 3502 24722
rect 3554 24670 3566 24722
rect 6962 24670 6974 24722
rect 7026 24670 7038 24722
rect 7646 24658 7698 24670
rect 9662 24722 9714 24734
rect 13246 24722 13298 24734
rect 17502 24722 17554 24734
rect 25678 24722 25730 24734
rect 32958 24722 33010 24734
rect 41358 24722 41410 24734
rect 10098 24670 10110 24722
rect 10162 24670 10174 24722
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 21186 24670 21198 24722
rect 21250 24670 21262 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 26338 24670 26350 24722
rect 26402 24670 26414 24722
rect 32162 24670 32174 24722
rect 32226 24670 32238 24722
rect 33618 24670 33630 24722
rect 33682 24670 33694 24722
rect 39442 24670 39454 24722
rect 39506 24670 39518 24722
rect 42018 24670 42030 24722
rect 42082 24670 42094 24722
rect 9662 24658 9714 24670
rect 13246 24658 13298 24670
rect 17502 24658 17554 24670
rect 25678 24658 25730 24670
rect 32958 24658 33010 24670
rect 41358 24658 41410 24670
rect 2494 24610 2546 24622
rect 37102 24610 37154 24622
rect 3602 24558 3614 24610
rect 3666 24558 3678 24610
rect 31042 24558 31054 24610
rect 31106 24558 31118 24610
rect 38546 24558 38558 24610
rect 38610 24558 38622 24610
rect 45714 24558 45726 24610
rect 45778 24558 45790 24610
rect 2494 24546 2546 24558
rect 37102 24546 37154 24558
rect 13134 24498 13186 24510
rect 13134 24434 13186 24446
rect 16942 24498 16994 24510
rect 16942 24434 16994 24446
rect 36654 24498 36706 24510
rect 36654 24434 36706 24446
rect 1344 24330 46592 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 46592 24330
rect 1344 24244 46592 24278
rect 8430 24050 8482 24062
rect 22206 24050 22258 24062
rect 36206 24050 36258 24062
rect 4050 23998 4062 24050
rect 4114 23998 4126 24050
rect 7858 23998 7870 24050
rect 7922 23998 7934 24050
rect 14914 23998 14926 24050
rect 14978 23998 14990 24050
rect 20402 23998 20414 24050
rect 20466 23998 20478 24050
rect 30146 23998 30158 24050
rect 30210 23998 30222 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 8430 23986 8482 23998
rect 22206 23986 22258 23998
rect 36206 23986 36258 23998
rect 36990 24050 37042 24062
rect 36990 23986 37042 23998
rect 42478 24050 42530 24062
rect 42802 23998 42814 24050
rect 42866 23998 42878 24050
rect 42478 23986 42530 23998
rect 9326 23938 9378 23950
rect 19966 23938 20018 23950
rect 29262 23938 29314 23950
rect 37886 23938 37938 23950
rect 41582 23938 41634 23950
rect 2034 23886 2046 23938
rect 2098 23886 2110 23938
rect 9650 23886 9662 23938
rect 9714 23886 9726 23938
rect 19282 23886 19294 23938
rect 19346 23886 19358 23938
rect 23314 23886 23326 23938
rect 23378 23886 23390 23938
rect 35410 23886 35422 23938
rect 35474 23886 35486 23938
rect 38546 23886 38558 23938
rect 38610 23886 38622 23938
rect 45042 23886 45054 23938
rect 45106 23886 45118 23938
rect 9326 23874 9378 23886
rect 19966 23874 20018 23886
rect 29262 23874 29314 23886
rect 37886 23874 37938 23886
rect 41582 23874 41634 23886
rect 5966 23826 6018 23838
rect 20750 23826 20802 23838
rect 21646 23826 21698 23838
rect 2258 23774 2270 23826
rect 2322 23774 2334 23826
rect 3042 23774 3054 23826
rect 3106 23774 3118 23826
rect 5618 23774 5630 23826
rect 5682 23774 5694 23826
rect 6626 23774 6638 23826
rect 6690 23774 6702 23826
rect 14018 23774 14030 23826
rect 14082 23774 14094 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 5966 23762 6018 23774
rect 20750 23762 20802 23774
rect 21646 23762 21698 23774
rect 22430 23826 22482 23838
rect 26786 23774 26798 23826
rect 26850 23774 26862 23826
rect 31154 23774 31166 23826
rect 31218 23774 31230 23826
rect 33954 23774 33966 23826
rect 34018 23774 34030 23826
rect 43810 23774 43822 23826
rect 43874 23774 43886 23826
rect 44818 23774 44830 23826
rect 44882 23774 44894 23826
rect 22430 23762 22482 23774
rect 8878 23714 8930 23726
rect 12798 23714 12850 23726
rect 12226 23662 12238 23714
rect 12290 23662 12302 23714
rect 8878 23650 8930 23662
rect 12798 23650 12850 23662
rect 16270 23714 16322 23726
rect 22542 23714 22594 23726
rect 17042 23662 17054 23714
rect 17106 23662 17118 23714
rect 16270 23650 16322 23662
rect 22542 23650 22594 23662
rect 37102 23714 37154 23726
rect 45614 23714 45666 23726
rect 40786 23662 40798 23714
rect 40850 23662 40862 23714
rect 37102 23650 37154 23662
rect 45614 23650 45666 23662
rect 46062 23714 46114 23726
rect 46062 23650 46114 23662
rect 1344 23546 46592 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 46592 23546
rect 1344 23460 46592 23494
rect 17502 23378 17554 23390
rect 23326 23378 23378 23390
rect 5506 23326 5518 23378
rect 5570 23326 5582 23378
rect 22530 23326 22542 23378
rect 22594 23326 22606 23378
rect 17502 23314 17554 23326
rect 23326 23314 23378 23326
rect 24334 23378 24386 23390
rect 24334 23314 24386 23326
rect 26574 23378 26626 23390
rect 30606 23378 30658 23390
rect 46062 23378 46114 23390
rect 30034 23326 30046 23378
rect 30098 23326 30110 23378
rect 37090 23326 37102 23378
rect 37154 23326 37166 23378
rect 45154 23326 45166 23378
rect 45218 23326 45230 23378
rect 26574 23314 26626 23326
rect 30606 23314 30658 23326
rect 46062 23314 46114 23326
rect 13918 23266 13970 23278
rect 13918 23202 13970 23214
rect 19406 23266 19458 23278
rect 19406 23202 19458 23214
rect 23886 23266 23938 23278
rect 23886 23202 23938 23214
rect 26014 23266 26066 23278
rect 32050 23214 32062 23266
rect 32114 23214 32126 23266
rect 33058 23214 33070 23266
rect 33122 23214 33134 23266
rect 38098 23214 38110 23266
rect 38162 23214 38174 23266
rect 39666 23214 39678 23266
rect 39730 23214 39742 23266
rect 40898 23214 40910 23266
rect 40962 23214 40974 23266
rect 26014 23202 26066 23214
rect 2606 23154 2658 23166
rect 16830 23154 16882 23166
rect 2034 23102 2046 23154
rect 2098 23102 2110 23154
rect 2930 23102 2942 23154
rect 2994 23102 3006 23154
rect 8866 23102 8878 23154
rect 8930 23102 8942 23154
rect 12562 23102 12574 23154
rect 12626 23102 12638 23154
rect 16146 23102 16158 23154
rect 16210 23102 16222 23154
rect 2606 23090 2658 23102
rect 16830 23090 16882 23102
rect 19630 23154 19682 23166
rect 26686 23154 26738 23166
rect 20178 23102 20190 23154
rect 20242 23102 20254 23154
rect 19630 23090 19682 23102
rect 26686 23090 26738 23102
rect 26910 23154 26962 23166
rect 34414 23154 34466 23166
rect 40014 23154 40066 23166
rect 42030 23154 42082 23166
rect 27570 23102 27582 23154
rect 27634 23102 27646 23154
rect 33282 23102 33294 23154
rect 33346 23102 33358 23154
rect 34850 23102 34862 23154
rect 34914 23102 34926 23154
rect 41122 23102 41134 23154
rect 41186 23102 41198 23154
rect 42578 23102 42590 23154
rect 42642 23102 42654 23154
rect 26910 23090 26962 23102
rect 34414 23090 34466 23102
rect 40014 23090 40066 23102
rect 42030 23090 42082 23102
rect 6526 23042 6578 23054
rect 1922 22990 1934 23042
rect 1986 22990 1998 23042
rect 6526 22978 6578 22990
rect 9662 23042 9714 23054
rect 9662 22978 9714 22990
rect 10222 23042 10274 23054
rect 10222 22978 10274 22990
rect 17390 23042 17442 23054
rect 17390 22978 17442 22990
rect 18174 23042 18226 23054
rect 31054 23042 31106 23054
rect 19058 22990 19070 23042
rect 19122 22990 19134 23042
rect 23538 22990 23550 23042
rect 23602 22990 23614 23042
rect 25778 22990 25790 23042
rect 25842 22990 25854 23042
rect 18174 22978 18226 22990
rect 31054 22978 31106 22990
rect 39118 23042 39170 23054
rect 39118 22978 39170 22990
rect 6078 22930 6130 22942
rect 6078 22866 6130 22878
rect 13134 22930 13186 22942
rect 13134 22866 13186 22878
rect 37886 22930 37938 22942
rect 37886 22866 37938 22878
rect 45726 22930 45778 22942
rect 45726 22866 45778 22878
rect 1344 22762 46592 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 46592 22762
rect 1344 22676 46592 22710
rect 16718 22482 16770 22494
rect 2146 22430 2158 22482
rect 2210 22430 2222 22482
rect 4050 22430 4062 22482
rect 4114 22430 4126 22482
rect 16718 22418 16770 22430
rect 40574 22482 40626 22494
rect 40574 22418 40626 22430
rect 5518 22370 5570 22382
rect 9550 22370 9602 22382
rect 17166 22370 17218 22382
rect 21422 22370 21474 22382
rect 25006 22370 25058 22382
rect 32734 22370 32786 22382
rect 2034 22318 2046 22370
rect 2098 22318 2110 22370
rect 6066 22318 6078 22370
rect 6130 22318 6142 22370
rect 9874 22318 9886 22370
rect 9938 22318 9950 22370
rect 13794 22318 13806 22370
rect 13858 22318 13870 22370
rect 17826 22318 17838 22370
rect 17890 22318 17902 22370
rect 21858 22318 21870 22370
rect 21922 22318 21934 22370
rect 25666 22318 25678 22370
rect 25730 22318 25742 22370
rect 32162 22318 32174 22370
rect 32226 22318 32238 22370
rect 5518 22306 5570 22318
rect 9550 22306 9602 22318
rect 17166 22306 17218 22318
rect 21422 22306 21474 22318
rect 25006 22306 25058 22318
rect 32734 22306 32786 22318
rect 33070 22370 33122 22382
rect 37102 22370 37154 22382
rect 33506 22318 33518 22370
rect 33570 22318 33582 22370
rect 37538 22318 37550 22370
rect 37602 22318 37614 22370
rect 40786 22318 40798 22370
rect 40850 22318 40862 22370
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 45042 22318 45054 22370
rect 45106 22318 45118 22370
rect 33070 22306 33122 22318
rect 37102 22306 37154 22318
rect 13022 22258 13074 22270
rect 3042 22206 3054 22258
rect 3106 22206 3118 22258
rect 16370 22206 16382 22258
rect 16434 22206 16446 22258
rect 13022 22194 13074 22206
rect 9214 22146 9266 22158
rect 14478 22146 14530 22158
rect 20862 22146 20914 22158
rect 24894 22146 24946 22158
rect 28702 22146 28754 22158
rect 8418 22094 8430 22146
rect 8482 22094 8494 22146
rect 12226 22094 12238 22146
rect 12290 22094 12302 22146
rect 20290 22094 20302 22146
rect 20354 22094 20366 22146
rect 24322 22094 24334 22146
rect 24386 22094 24398 22146
rect 28018 22094 28030 22146
rect 28082 22094 28094 22146
rect 9214 22082 9266 22094
rect 14478 22082 14530 22094
rect 20862 22082 20914 22094
rect 24894 22082 24946 22094
rect 28702 22082 28754 22094
rect 29038 22146 29090 22158
rect 36542 22146 36594 22158
rect 44382 22146 44434 22158
rect 46286 22146 46338 22158
rect 29810 22094 29822 22146
rect 29874 22094 29886 22146
rect 35746 22094 35758 22146
rect 35810 22094 35822 22146
rect 39890 22094 39902 22146
rect 39954 22094 39966 22146
rect 43810 22094 43822 22146
rect 43874 22094 43886 22146
rect 44818 22094 44830 22146
rect 44882 22094 44894 22146
rect 29038 22082 29090 22094
rect 36542 22082 36594 22094
rect 44382 22082 44434 22094
rect 46286 22082 46338 22094
rect 1344 21978 46592 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 46592 21978
rect 1344 21892 46592 21926
rect 2482 21758 2494 21810
rect 2546 21758 2558 21810
rect 15026 21758 15038 21810
rect 15090 21758 15102 21810
rect 21186 21758 21198 21810
rect 21250 21758 21262 21810
rect 28466 21758 28478 21810
rect 28530 21758 28542 21810
rect 39890 21758 39902 21810
rect 39954 21758 39966 21810
rect 11230 21698 11282 21710
rect 6066 21646 6078 21698
rect 6130 21646 6142 21698
rect 11230 21634 11282 21646
rect 11566 21698 11618 21710
rect 16718 21698 16770 21710
rect 32510 21698 32562 21710
rect 11890 21646 11902 21698
rect 11954 21646 11966 21698
rect 16370 21646 16382 21698
rect 16434 21646 16446 21698
rect 24322 21646 24334 21698
rect 24386 21646 24398 21698
rect 32162 21646 32174 21698
rect 32226 21646 32238 21698
rect 11566 21634 11618 21646
rect 16718 21634 16770 21646
rect 32510 21634 32562 21646
rect 35870 21698 35922 21710
rect 35870 21634 35922 21646
rect 43710 21698 43762 21710
rect 43710 21634 43762 21646
rect 5406 21586 5458 21598
rect 12126 21586 12178 21598
rect 23886 21586 23938 21598
rect 25342 21586 25394 21598
rect 33182 21586 33234 21598
rect 36990 21586 37042 21598
rect 40798 21586 40850 21598
rect 4722 21534 4734 21586
rect 4786 21534 4798 21586
rect 5842 21534 5854 21586
rect 5906 21534 5918 21586
rect 8530 21534 8542 21586
rect 8594 21534 8606 21586
rect 9874 21534 9886 21586
rect 9938 21534 9950 21586
rect 12674 21534 12686 21586
rect 12738 21534 12750 21586
rect 17938 21534 17950 21586
rect 18002 21534 18014 21586
rect 23426 21534 23438 21586
rect 23490 21534 23502 21586
rect 24546 21534 24558 21586
rect 24610 21534 24622 21586
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 31266 21534 31278 21586
rect 31330 21534 31342 21586
rect 33618 21534 33630 21586
rect 33682 21534 33694 21586
rect 37314 21534 37326 21586
rect 37378 21534 37390 21586
rect 41458 21534 41470 21586
rect 41522 21534 41534 21586
rect 45042 21534 45054 21586
rect 45106 21534 45118 21586
rect 45602 21534 45614 21586
rect 45666 21534 45678 21586
rect 5406 21522 5458 21534
rect 12126 21522 12178 21534
rect 23886 21522 23938 21534
rect 25342 21522 25394 21534
rect 33182 21522 33234 21534
rect 36990 21522 37042 21534
rect 40798 21522 40850 21534
rect 10558 21474 10610 21486
rect 6626 21422 6638 21474
rect 6690 21422 6702 21474
rect 9650 21422 9662 21474
rect 9714 21422 9726 21474
rect 10882 21422 10894 21474
rect 10946 21422 10958 21474
rect 18498 21422 18510 21474
rect 18562 21422 18574 21474
rect 29474 21422 29486 21474
rect 29538 21422 29550 21474
rect 45714 21422 45726 21474
rect 45778 21422 45790 21474
rect 10558 21410 10610 21422
rect 1710 21362 1762 21374
rect 1710 21298 1762 21310
rect 15822 21362 15874 21374
rect 15822 21298 15874 21310
rect 20414 21362 20466 21374
rect 20414 21298 20466 21310
rect 29038 21362 29090 21374
rect 29038 21298 29090 21310
rect 36654 21362 36706 21374
rect 36654 21298 36706 21310
rect 40462 21362 40514 21374
rect 40462 21298 40514 21310
rect 44494 21362 44546 21374
rect 44706 21310 44718 21362
rect 44770 21310 44782 21362
rect 44494 21298 44546 21310
rect 1344 21194 46592 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 46592 21194
rect 1344 21108 46592 21142
rect 28590 20914 28642 20926
rect 3826 20862 3838 20914
rect 3890 20862 3902 20914
rect 21522 20862 21534 20914
rect 21586 20862 21598 20914
rect 33954 20862 33966 20914
rect 34018 20862 34030 20914
rect 28590 20850 28642 20862
rect 5518 20802 5570 20814
rect 13022 20802 13074 20814
rect 2034 20750 2046 20802
rect 2098 20750 2110 20802
rect 6178 20750 6190 20802
rect 6242 20750 6254 20802
rect 12450 20750 12462 20802
rect 12514 20750 12526 20802
rect 5518 20738 5570 20750
rect 13022 20738 13074 20750
rect 13358 20802 13410 20814
rect 20862 20802 20914 20814
rect 24446 20802 24498 20814
rect 29262 20802 29314 20814
rect 37102 20802 37154 20814
rect 40686 20802 40738 20814
rect 14018 20750 14030 20802
rect 14082 20750 14094 20802
rect 20178 20750 20190 20802
rect 20242 20750 20254 20802
rect 23650 20750 23662 20802
rect 23714 20750 23726 20802
rect 25106 20750 25118 20802
rect 25170 20750 25182 20802
rect 29698 20750 29710 20802
rect 29762 20750 29774 20802
rect 37426 20750 37438 20802
rect 37490 20750 37502 20802
rect 41234 20750 41246 20802
rect 41298 20750 41310 20802
rect 45042 20750 45054 20802
rect 45106 20750 45118 20802
rect 13358 20738 13410 20750
rect 20862 20738 20914 20750
rect 24446 20738 24498 20750
rect 29262 20738 29314 20750
rect 37102 20738 37154 20750
rect 40686 20738 40738 20750
rect 9326 20690 9378 20702
rect 2258 20638 2270 20690
rect 2322 20638 2334 20690
rect 3042 20638 3054 20690
rect 3106 20638 3118 20690
rect 9326 20626 9378 20638
rect 10110 20690 10162 20702
rect 36094 20690 36146 20702
rect 34962 20638 34974 20690
rect 35026 20638 35038 20690
rect 10110 20626 10162 20638
rect 36094 20626 36146 20638
rect 46174 20690 46226 20702
rect 46174 20626 46226 20638
rect 9214 20578 9266 20590
rect 17054 20578 17106 20590
rect 8642 20526 8654 20578
rect 8706 20526 8718 20578
rect 16370 20526 16382 20578
rect 16434 20526 16446 20578
rect 9214 20514 9266 20526
rect 17054 20514 17106 20526
rect 17166 20578 17218 20590
rect 28142 20578 28194 20590
rect 32734 20578 32786 20590
rect 17938 20526 17950 20578
rect 18002 20526 18014 20578
rect 27570 20526 27582 20578
rect 27634 20526 27646 20578
rect 32162 20526 32174 20578
rect 32226 20526 32238 20578
rect 17166 20514 17218 20526
rect 28142 20514 28194 20526
rect 32734 20514 32786 20526
rect 33630 20578 33682 20590
rect 33630 20514 33682 20526
rect 35982 20578 36034 20590
rect 40574 20578 40626 20590
rect 44382 20578 44434 20590
rect 45838 20578 45890 20590
rect 40002 20526 40014 20578
rect 40066 20526 40078 20578
rect 43810 20526 43822 20578
rect 43874 20526 43886 20578
rect 44818 20526 44830 20578
rect 44882 20526 44894 20578
rect 35982 20514 36034 20526
rect 40574 20514 40626 20526
rect 44382 20514 44434 20526
rect 45838 20514 45890 20526
rect 1344 20410 46592 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 46592 20410
rect 1344 20324 46592 20358
rect 2482 20190 2494 20242
rect 2546 20190 2558 20242
rect 40338 20190 40350 20242
rect 40402 20190 40414 20242
rect 10222 20130 10274 20142
rect 10222 20066 10274 20078
rect 16158 20130 16210 20142
rect 16158 20066 16210 20078
rect 20414 20130 20466 20142
rect 20414 20066 20466 20078
rect 23998 20130 24050 20142
rect 23998 20066 24050 20078
rect 26910 20130 26962 20142
rect 39230 20130 39282 20142
rect 32050 20078 32062 20130
rect 32114 20078 32126 20130
rect 38882 20078 38894 20130
rect 38946 20078 38958 20130
rect 42914 20078 42926 20130
rect 42978 20078 42990 20130
rect 45714 20078 45726 20130
rect 45778 20078 45790 20130
rect 26910 20066 26962 20078
rect 39230 20066 39282 20078
rect 5406 20018 5458 20030
rect 13246 20018 13298 20030
rect 21086 20018 21138 20030
rect 29598 20018 29650 20030
rect 4946 19966 4958 20018
rect 5010 19966 5022 20018
rect 8530 19966 8542 20018
rect 8594 19966 8606 20018
rect 12450 19966 12462 20018
rect 12514 19966 12526 20018
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 13906 19966 13918 20018
rect 13970 19966 13982 20018
rect 17826 19966 17838 20018
rect 17890 19966 17902 20018
rect 21746 19966 21758 20018
rect 21810 19966 21822 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 29138 19966 29150 20018
rect 29202 19966 29214 20018
rect 33058 19966 33070 20018
rect 33122 19966 33134 20018
rect 33282 19966 33294 20018
rect 33346 19966 33358 20018
rect 33954 19966 33966 20018
rect 34018 19966 34030 20018
rect 34626 19966 34638 20018
rect 34690 19966 34702 20018
rect 39778 19966 39790 20018
rect 39842 19966 39854 20018
rect 5406 19954 5458 19966
rect 13246 19954 13298 19966
rect 21086 19954 21138 19966
rect 29598 19954 29650 19966
rect 20862 19906 20914 19918
rect 43822 19906 43874 19918
rect 44494 19906 44546 19918
rect 7858 19854 7870 19906
rect 7922 19854 7934 19906
rect 18610 19854 18622 19906
rect 18674 19854 18686 19906
rect 25218 19854 25230 19906
rect 25282 19854 25294 19906
rect 31042 19854 31054 19906
rect 31106 19854 31118 19906
rect 33730 19854 33742 19906
rect 33794 19854 33806 19906
rect 41906 19854 41918 19906
rect 41970 19854 41982 19906
rect 44146 19854 44158 19906
rect 44210 19854 44222 19906
rect 44930 19854 44942 19906
rect 44994 19854 45006 19906
rect 20862 19842 20914 19854
rect 43822 19842 43874 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 9438 19794 9490 19806
rect 9438 19730 9490 19742
rect 16942 19794 16994 19806
rect 16942 19730 16994 19742
rect 24782 19794 24834 19806
rect 24782 19730 24834 19742
rect 26126 19794 26178 19806
rect 26126 19730 26178 19742
rect 38334 19794 38386 19806
rect 43810 19742 43822 19794
rect 43874 19791 43886 19794
rect 44161 19791 44207 19854
rect 44494 19842 44546 19854
rect 43874 19745 44207 19791
rect 43874 19742 43886 19745
rect 38334 19730 38386 19742
rect 1344 19626 46592 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 46592 19626
rect 1344 19540 46592 19574
rect 43474 19406 43486 19458
rect 43538 19406 43550 19458
rect 7646 19346 7698 19358
rect 3826 19294 3838 19346
rect 3890 19294 3902 19346
rect 6850 19294 6862 19346
rect 6914 19294 6926 19346
rect 7646 19282 7698 19294
rect 8094 19346 8146 19358
rect 21758 19346 21810 19358
rect 19170 19294 19182 19346
rect 19234 19294 19246 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 8094 19282 8146 19294
rect 21758 19282 21810 19294
rect 27806 19346 27858 19358
rect 27806 19282 27858 19294
rect 35982 19346 36034 19358
rect 44158 19346 44210 19358
rect 38546 19294 38558 19346
rect 38610 19294 38622 19346
rect 41122 19294 41134 19346
rect 41186 19294 41198 19346
rect 43810 19294 43822 19346
rect 43874 19294 43886 19346
rect 35982 19282 36034 19294
rect 44158 19282 44210 19294
rect 8542 19234 8594 19246
rect 14926 19234 14978 19246
rect 18846 19234 18898 19246
rect 2034 19182 2046 19234
rect 2098 19182 2110 19234
rect 8978 19182 8990 19234
rect 9042 19182 9054 19234
rect 13682 19182 13694 19234
rect 13746 19182 13758 19234
rect 14354 19182 14366 19234
rect 14418 19182 14430 19234
rect 18274 19182 18286 19234
rect 18338 19182 18350 19234
rect 8542 19170 8594 19182
rect 14926 19170 14978 19182
rect 18846 19170 18898 19182
rect 19406 19234 19458 19246
rect 25790 19234 25842 19246
rect 25442 19182 25454 19234
rect 25506 19182 25518 19234
rect 19406 19170 19458 19182
rect 25790 19170 25842 19182
rect 29374 19234 29426 19246
rect 29810 19182 29822 19234
rect 29874 19182 29886 19234
rect 33506 19182 33518 19234
rect 33570 19182 33582 19234
rect 39442 19182 39454 19234
rect 39506 19182 39518 19234
rect 42914 19182 42926 19234
rect 42978 19182 42990 19234
rect 44930 19182 44942 19234
rect 44994 19182 45006 19234
rect 29374 19170 29426 19182
rect 12574 19122 12626 19134
rect 19742 19122 19794 19134
rect 2258 19070 2270 19122
rect 2322 19070 2334 19122
rect 2818 19070 2830 19122
rect 2882 19070 2894 19122
rect 6066 19070 6078 19122
rect 6130 19070 6142 19122
rect 12226 19070 12238 19122
rect 12290 19070 12302 19122
rect 13458 19070 13470 19122
rect 13522 19070 13534 19122
rect 14130 19070 14142 19122
rect 14194 19070 14206 19122
rect 12574 19058 12626 19070
rect 19742 19058 19794 19070
rect 23102 19122 23154 19134
rect 42130 19070 42142 19122
rect 42194 19070 42206 19122
rect 46050 19070 46062 19122
rect 46114 19070 46126 19122
rect 23102 19058 23154 19070
rect 12014 19010 12066 19022
rect 11442 18958 11454 19010
rect 11506 18958 11518 19010
rect 12014 18946 12066 18958
rect 15150 19010 15202 19022
rect 19854 19010 19906 19022
rect 15922 18958 15934 19010
rect 15986 18958 15998 19010
rect 15150 18946 15202 18958
rect 19854 18946 19906 18958
rect 22318 19010 22370 19022
rect 32846 19010 32898 19022
rect 32274 18958 32286 19010
rect 32338 18958 32350 19010
rect 22318 18946 22370 18958
rect 32846 18946 32898 18958
rect 34078 19010 34130 19022
rect 34078 18946 34130 18958
rect 36094 19010 36146 19022
rect 36094 18946 36146 18958
rect 1344 18842 46592 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 46592 18842
rect 1344 18756 46592 18790
rect 32510 18674 32562 18686
rect 2146 18622 2158 18674
rect 2210 18622 2222 18674
rect 5954 18622 5966 18674
rect 6018 18622 6030 18674
rect 16370 18622 16382 18674
rect 16434 18622 16446 18674
rect 32510 18610 32562 18622
rect 10222 18562 10274 18574
rect 10222 18498 10274 18510
rect 18622 18562 18674 18574
rect 18622 18498 18674 18510
rect 22094 18562 22146 18574
rect 35870 18562 35922 18574
rect 23986 18510 23998 18562
rect 24050 18510 24062 18562
rect 31042 18510 31054 18562
rect 31106 18510 31118 18562
rect 22094 18498 22146 18510
rect 35870 18498 35922 18510
rect 41582 18562 41634 18574
rect 41582 18498 41634 18510
rect 5294 18450 5346 18462
rect 8878 18450 8930 18462
rect 13246 18450 13298 18462
rect 18174 18450 18226 18462
rect 4722 18398 4734 18450
rect 4786 18398 4798 18450
rect 8418 18398 8430 18450
rect 8482 18398 8494 18450
rect 12562 18398 12574 18450
rect 12626 18398 12638 18450
rect 13010 18398 13022 18450
rect 13074 18398 13086 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 17826 18398 17838 18450
rect 17890 18398 17902 18450
rect 5294 18386 5346 18398
rect 8878 18386 8930 18398
rect 13246 18386 13298 18398
rect 18174 18386 18226 18398
rect 19182 18450 19234 18462
rect 23662 18450 23714 18462
rect 19730 18398 19742 18450
rect 19794 18398 19806 18450
rect 19182 18386 19234 18398
rect 23662 18386 23714 18398
rect 24334 18450 24386 18462
rect 33182 18450 33234 18462
rect 36990 18450 37042 18462
rect 40350 18450 40402 18462
rect 25666 18398 25678 18450
rect 25730 18398 25742 18450
rect 30258 18398 30270 18450
rect 30322 18398 30334 18450
rect 31714 18398 31726 18450
rect 31778 18398 31790 18450
rect 31938 18398 31950 18450
rect 32002 18398 32014 18450
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 39442 18398 39454 18450
rect 39506 18398 39518 18450
rect 43810 18398 43822 18450
rect 43874 18398 43886 18450
rect 44370 18398 44382 18450
rect 44434 18398 44446 18450
rect 44930 18398 44942 18450
rect 44994 18398 45006 18450
rect 24334 18386 24386 18398
rect 33182 18386 33234 18398
rect 36990 18386 37042 18398
rect 40350 18386 40402 18398
rect 31390 18338 31442 18350
rect 18946 18286 18958 18338
rect 19010 18286 19022 18338
rect 23314 18286 23326 18338
rect 23378 18286 23390 18338
rect 28578 18286 28590 18338
rect 28642 18286 28654 18338
rect 37538 18286 37550 18338
rect 37602 18286 37614 18338
rect 46050 18286 46062 18338
rect 46114 18286 46126 18338
rect 31390 18274 31442 18286
rect 1598 18226 1650 18238
rect 1598 18162 1650 18174
rect 5406 18226 5458 18238
rect 5406 18162 5458 18174
rect 9438 18226 9490 18238
rect 9438 18162 9490 18174
rect 16942 18226 16994 18238
rect 16942 18162 16994 18174
rect 22878 18226 22930 18238
rect 22878 18162 22930 18174
rect 27582 18226 27634 18238
rect 27582 18162 27634 18174
rect 36654 18226 36706 18238
rect 36654 18162 36706 18174
rect 40798 18226 40850 18238
rect 40798 18162 40850 18174
rect 1344 18058 46592 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 46592 18058
rect 1344 17972 46592 18006
rect 21870 17778 21922 17790
rect 3938 17726 3950 17778
rect 4002 17726 4014 17778
rect 8306 17726 8318 17778
rect 8370 17726 8382 17778
rect 15250 17726 15262 17778
rect 15314 17726 15326 17778
rect 21634 17726 21646 17778
rect 21698 17726 21710 17778
rect 21870 17714 21922 17726
rect 22542 17778 22594 17790
rect 22542 17714 22594 17726
rect 28254 17778 28306 17790
rect 28254 17714 28306 17726
rect 30270 17778 30322 17790
rect 36094 17778 36146 17790
rect 34402 17726 34414 17778
rect 34466 17726 34478 17778
rect 35746 17726 35758 17778
rect 35810 17726 35822 17778
rect 42242 17726 42254 17778
rect 42306 17726 42318 17778
rect 30270 17714 30322 17726
rect 36094 17714 36146 17726
rect 9214 17666 9266 17678
rect 16942 17666 16994 17678
rect 22766 17666 22818 17678
rect 30494 17666 30546 17678
rect 37326 17666 37378 17678
rect 2034 17614 2046 17666
rect 2098 17614 2110 17666
rect 6626 17614 6638 17666
rect 6690 17614 6702 17666
rect 9650 17614 9662 17666
rect 9714 17614 9726 17666
rect 13794 17614 13806 17666
rect 13858 17614 13870 17666
rect 17490 17614 17502 17666
rect 17554 17614 17566 17666
rect 23426 17614 23438 17666
rect 23490 17614 23502 17666
rect 27570 17614 27582 17666
rect 27634 17614 27646 17666
rect 31154 17614 31166 17666
rect 31218 17614 31230 17666
rect 34626 17614 34638 17666
rect 34690 17614 34702 17666
rect 35298 17614 35310 17666
rect 35362 17614 35374 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 45154 17614 45166 17666
rect 45218 17614 45230 17666
rect 9214 17602 9266 17614
rect 16942 17602 16994 17614
rect 22766 17602 22818 17614
rect 30494 17602 30546 17614
rect 37326 17602 37378 17614
rect 19854 17554 19906 17566
rect 27022 17554 27074 17566
rect 44270 17554 44322 17566
rect 2258 17502 2270 17554
rect 2322 17502 2334 17554
rect 3042 17502 3054 17554
rect 3106 17502 3118 17554
rect 13570 17502 13582 17554
rect 13634 17502 13646 17554
rect 16482 17502 16494 17554
rect 16546 17502 16558 17554
rect 22194 17502 22206 17554
rect 22258 17502 22270 17554
rect 26674 17502 26686 17554
rect 26738 17502 26750 17554
rect 27794 17502 27806 17554
rect 27858 17502 27870 17554
rect 35074 17502 35086 17554
rect 35138 17502 35150 17554
rect 43250 17502 43262 17554
rect 43314 17502 43326 17554
rect 46050 17502 46062 17554
rect 46114 17502 46126 17554
rect 19854 17490 19906 17502
rect 27022 17490 27074 17502
rect 44270 17490 44322 17502
rect 5070 17442 5122 17454
rect 5070 17378 5122 17390
rect 5854 17442 5906 17454
rect 12686 17442 12738 17454
rect 12114 17390 12126 17442
rect 12178 17390 12190 17442
rect 5854 17378 5906 17390
rect 12686 17378 12738 17390
rect 14366 17442 14418 17454
rect 14366 17378 14418 17390
rect 14814 17442 14866 17454
rect 14814 17378 14866 17390
rect 20638 17442 20690 17454
rect 26462 17442 26514 17454
rect 25890 17390 25902 17442
rect 25954 17390 25966 17442
rect 20638 17378 20690 17390
rect 26462 17378 26514 17390
rect 30158 17442 30210 17454
rect 34190 17442 34242 17454
rect 40798 17442 40850 17454
rect 33618 17390 33630 17442
rect 33682 17390 33694 17442
rect 40002 17390 40014 17442
rect 40066 17390 40078 17442
rect 30158 17378 30210 17390
rect 34190 17378 34242 17390
rect 40798 17378 40850 17390
rect 1344 17274 46592 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 46592 17274
rect 1344 17188 46592 17222
rect 2146 17054 2158 17106
rect 2210 17054 2222 17106
rect 24098 17054 24110 17106
rect 24162 17054 24174 17106
rect 36082 17054 36094 17106
rect 36146 17054 36158 17106
rect 8318 16994 8370 17006
rect 8318 16930 8370 16942
rect 10222 16994 10274 17006
rect 18062 16994 18114 17006
rect 25902 16994 25954 17006
rect 13458 16942 13470 16994
rect 13522 16942 13534 16994
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 17714 16942 17726 16994
rect 17778 16942 17790 16994
rect 18834 16942 18846 16994
rect 18898 16942 18910 16994
rect 10222 16930 10274 16942
rect 18062 16930 18114 16942
rect 25902 16930 25954 16942
rect 31838 16994 31890 17006
rect 31838 16930 31890 16942
rect 36654 16994 36706 17006
rect 36654 16930 36706 16942
rect 39678 16994 39730 17006
rect 39678 16930 39730 16942
rect 43710 16994 43762 17006
rect 43710 16930 43762 16942
rect 5070 16882 5122 16894
rect 4610 16830 4622 16882
rect 4674 16830 4686 16882
rect 5070 16818 5122 16830
rect 5406 16882 5458 16894
rect 21086 16882 21138 16894
rect 28814 16882 28866 16894
rect 6066 16830 6078 16882
rect 6130 16830 6142 16882
rect 12450 16830 12462 16882
rect 12514 16830 12526 16882
rect 13010 16830 13022 16882
rect 13074 16830 13086 16882
rect 13682 16830 13694 16882
rect 13746 16830 13758 16882
rect 21746 16830 21758 16882
rect 21810 16830 21822 16882
rect 28242 16830 28254 16882
rect 28306 16830 28318 16882
rect 5406 16818 5458 16830
rect 21086 16818 21138 16830
rect 28814 16818 28866 16830
rect 28926 16882 28978 16894
rect 33182 16882 33234 16894
rect 36990 16882 37042 16894
rect 41022 16882 41074 16894
rect 44494 16882 44546 16894
rect 46062 16882 46114 16894
rect 29474 16830 29486 16882
rect 29538 16830 29550 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 37314 16830 37326 16882
rect 37378 16830 37390 16882
rect 41458 16830 41470 16882
rect 41522 16830 41534 16882
rect 44930 16830 44942 16882
rect 44994 16830 45006 16882
rect 28926 16818 28978 16830
rect 33182 16818 33234 16830
rect 36990 16818 37042 16830
rect 41022 16818 41074 16830
rect 44494 16818 44546 16830
rect 46062 16818 46114 16830
rect 15810 16718 15822 16770
rect 15874 16718 15886 16770
rect 19618 16718 19630 16770
rect 19682 16718 19694 16770
rect 1598 16658 1650 16670
rect 1598 16594 1650 16606
rect 9102 16658 9154 16670
rect 9102 16594 9154 16606
rect 9438 16658 9490 16670
rect 9438 16594 9490 16606
rect 24782 16658 24834 16670
rect 24782 16594 24834 16606
rect 25118 16658 25170 16670
rect 25118 16594 25170 16606
rect 32622 16658 32674 16670
rect 32622 16594 32674 16606
rect 40462 16658 40514 16670
rect 40462 16594 40514 16606
rect 1344 16490 46592 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 46592 16490
rect 1344 16404 46592 16438
rect 1934 16210 1986 16222
rect 13582 16210 13634 16222
rect 4050 16158 4062 16210
rect 4114 16158 4126 16210
rect 6626 16158 6638 16210
rect 6690 16158 6702 16210
rect 1934 16146 1986 16158
rect 13582 16146 13634 16158
rect 18958 16210 19010 16222
rect 45490 16158 45502 16210
rect 45554 16158 45566 16210
rect 18958 16146 19010 16158
rect 8542 16098 8594 16110
rect 14926 16098 14978 16110
rect 24894 16098 24946 16110
rect 29038 16098 29090 16110
rect 33070 16098 33122 16110
rect 40574 16098 40626 16110
rect 8866 16046 8878 16098
rect 8930 16046 8942 16098
rect 15250 16046 15262 16098
rect 15314 16046 15326 16098
rect 24210 16046 24222 16098
rect 24274 16046 24286 16098
rect 25106 16046 25118 16098
rect 25170 16046 25182 16098
rect 25666 16046 25678 16098
rect 25730 16046 25742 16098
rect 29698 16046 29710 16098
rect 29762 16046 29774 16098
rect 33506 16046 33518 16098
rect 33570 16046 33582 16098
rect 39890 16046 39902 16098
rect 39954 16046 39966 16098
rect 8542 16034 8594 16046
rect 14926 16034 14978 16046
rect 24894 16034 24946 16046
rect 29038 16034 29090 16046
rect 33070 16034 33122 16046
rect 40574 16034 40626 16046
rect 40910 16098 40962 16110
rect 41346 16046 41358 16098
rect 41410 16046 41422 16098
rect 45938 16046 45950 16098
rect 46002 16046 46014 16098
rect 40910 16034 40962 16046
rect 21982 15986 22034 15998
rect 2258 15934 2270 15986
rect 2322 15934 2334 15986
rect 2706 15934 2718 15986
rect 2770 15934 2782 15986
rect 7746 15934 7758 15986
rect 7810 15934 7822 15986
rect 18610 15934 18622 15986
rect 18674 15934 18686 15986
rect 21982 15922 22034 15934
rect 27918 15986 27970 15998
rect 27918 15922 27970 15934
rect 43598 15986 43650 15998
rect 43598 15922 43650 15934
rect 5742 15874 5794 15886
rect 5742 15810 5794 15822
rect 6302 15874 6354 15886
rect 12014 15874 12066 15886
rect 11442 15822 11454 15874
rect 11506 15822 11518 15874
rect 6302 15810 6354 15822
rect 12014 15810 12066 15822
rect 12350 15874 12402 15886
rect 12350 15810 12402 15822
rect 12910 15874 12962 15886
rect 12910 15810 12962 15822
rect 14030 15874 14082 15886
rect 18398 15874 18450 15886
rect 17826 15822 17838 15874
rect 17890 15822 17902 15874
rect 14030 15810 14082 15822
rect 18398 15810 18450 15822
rect 21198 15874 21250 15886
rect 21198 15810 21250 15822
rect 28702 15874 28754 15886
rect 32734 15874 32786 15886
rect 36542 15874 36594 15886
rect 32162 15822 32174 15874
rect 32226 15822 32238 15874
rect 35746 15822 35758 15874
rect 35810 15822 35822 15874
rect 28702 15810 28754 15822
rect 32734 15810 32786 15822
rect 36542 15810 36594 15822
rect 36878 15874 36930 15886
rect 44382 15874 44434 15886
rect 37538 15822 37550 15874
rect 37602 15822 37614 15874
rect 36878 15810 36930 15822
rect 44382 15810 44434 15822
rect 1344 15706 46592 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 46592 15706
rect 1344 15620 46592 15654
rect 1934 15538 1986 15550
rect 10334 15538 10386 15550
rect 28142 15538 28194 15550
rect 41022 15538 41074 15550
rect 45726 15538 45778 15550
rect 8194 15486 8206 15538
rect 8258 15486 8270 15538
rect 23202 15486 23214 15538
rect 23266 15486 23278 15538
rect 31602 15486 31614 15538
rect 31666 15486 31678 15538
rect 44818 15486 44830 15538
rect 44882 15486 44894 15538
rect 1934 15474 1986 15486
rect 10334 15474 10386 15486
rect 28142 15474 28194 15486
rect 41022 15474 41074 15486
rect 45726 15474 45778 15486
rect 24334 15426 24386 15438
rect 28030 15426 28082 15438
rect 3378 15374 3390 15426
rect 3442 15374 3454 15426
rect 9538 15374 9550 15426
rect 9602 15374 9614 15426
rect 11890 15374 11902 15426
rect 11954 15374 11966 15426
rect 15698 15374 15710 15426
rect 15762 15374 15774 15426
rect 17490 15374 17502 15426
rect 17554 15374 17566 15426
rect 24658 15374 24670 15426
rect 24722 15374 24734 15426
rect 27346 15374 27358 15426
rect 27410 15374 27422 15426
rect 24334 15362 24386 15374
rect 28030 15362 28082 15374
rect 33742 15426 33794 15438
rect 45390 15426 45442 15438
rect 39442 15374 39454 15426
rect 39506 15374 39518 15426
rect 33742 15362 33794 15374
rect 45390 15362 45442 15374
rect 5070 15314 5122 15326
rect 20190 15314 20242 15326
rect 28926 15314 28978 15326
rect 36654 15314 36706 15326
rect 41694 15314 41746 15326
rect 1922 15262 1934 15314
rect 1986 15262 1998 15314
rect 5618 15262 5630 15314
rect 5682 15262 5694 15314
rect 20850 15262 20862 15314
rect 20914 15262 20926 15314
rect 29250 15262 29262 15314
rect 29314 15262 29326 15314
rect 35970 15262 35982 15314
rect 36034 15262 36046 15314
rect 41122 15262 41134 15314
rect 41186 15262 41198 15314
rect 42354 15262 42366 15314
rect 42418 15262 42430 15314
rect 45602 15262 45614 15314
rect 45666 15262 45678 15314
rect 5070 15250 5122 15262
rect 20190 15250 20242 15262
rect 28926 15250 28978 15262
rect 36654 15250 36706 15262
rect 41694 15250 41746 15262
rect 9886 15202 9938 15214
rect 2594 15150 2606 15202
rect 2658 15150 2670 15202
rect 9886 15138 9938 15150
rect 10782 15202 10834 15214
rect 12786 15150 12798 15202
rect 12850 15150 12862 15202
rect 14578 15150 14590 15202
rect 14642 15150 14654 15202
rect 18722 15150 18734 15202
rect 18786 15150 18798 15202
rect 26226 15150 26238 15202
rect 26290 15150 26302 15202
rect 38322 15150 38334 15202
rect 38386 15150 38398 15202
rect 10782 15138 10834 15150
rect 8766 15090 8818 15102
rect 8766 15026 8818 15038
rect 23886 15090 23938 15102
rect 23886 15026 23938 15038
rect 32398 15090 32450 15102
rect 32398 15026 32450 15038
rect 32958 15090 33010 15102
rect 32958 15026 33010 15038
rect 1344 14922 46592 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 46592 14922
rect 1344 14836 46592 14870
rect 9662 14642 9714 14654
rect 3826 14590 3838 14642
rect 3890 14590 3902 14642
rect 9662 14578 9714 14590
rect 9998 14642 10050 14654
rect 10434 14590 10446 14642
rect 10498 14590 10510 14642
rect 16258 14590 16270 14642
rect 16322 14590 16334 14642
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 34626 14590 34638 14642
rect 34690 14590 34702 14642
rect 37986 14590 37998 14642
rect 38050 14590 38062 14642
rect 40002 14590 40014 14642
rect 40066 14590 40078 14642
rect 42802 14590 42814 14642
rect 42866 14590 42878 14642
rect 9998 14578 10050 14590
rect 9214 14530 9266 14542
rect 8642 14478 8654 14530
rect 8706 14478 8718 14530
rect 9214 14466 9266 14478
rect 23998 14530 24050 14542
rect 29710 14530 29762 14542
rect 24434 14478 24446 14530
rect 24498 14478 24510 14530
rect 30370 14478 30382 14530
rect 30434 14478 30446 14530
rect 39778 14478 39790 14530
rect 39842 14478 39854 14530
rect 44818 14478 44830 14530
rect 44882 14478 44894 14530
rect 23998 14466 24050 14478
rect 29710 14466 29762 14478
rect 1934 14418 1986 14430
rect 26686 14418 26738 14430
rect 4946 14366 4958 14418
rect 5010 14366 5022 14418
rect 11666 14366 11678 14418
rect 11730 14366 11742 14418
rect 15026 14366 15038 14418
rect 15090 14366 15102 14418
rect 19730 14366 19742 14418
rect 19794 14366 19806 14418
rect 35634 14366 35646 14418
rect 35698 14366 35710 14418
rect 38994 14366 39006 14418
rect 39058 14366 39070 14418
rect 43922 14366 43934 14418
rect 43986 14366 43998 14418
rect 45938 14366 45950 14418
rect 46002 14366 46014 14418
rect 1934 14354 1986 14366
rect 26686 14354 26738 14366
rect 2046 14306 2098 14318
rect 2046 14242 2098 14254
rect 2718 14306 2770 14318
rect 2718 14242 2770 14254
rect 3166 14306 3218 14318
rect 3166 14242 3218 14254
rect 5518 14306 5570 14318
rect 27470 14306 27522 14318
rect 33406 14306 33458 14318
rect 6178 14254 6190 14306
rect 6242 14254 6254 14306
rect 32834 14254 32846 14306
rect 32898 14254 32910 14306
rect 5518 14242 5570 14254
rect 27470 14242 27522 14254
rect 33406 14242 33458 14254
rect 1344 14138 46592 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 46592 14138
rect 1344 14052 46592 14086
rect 8878 13970 8930 13982
rect 4834 13918 4846 13970
rect 4898 13918 4910 13970
rect 8878 13906 8930 13918
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 32510 13858 32562 13870
rect 33406 13858 33458 13870
rect 34078 13858 34130 13870
rect 6178 13806 6190 13858
rect 6242 13806 6254 13858
rect 6962 13806 6974 13858
rect 7026 13806 7038 13858
rect 13570 13806 13582 13858
rect 13634 13806 13646 13858
rect 16370 13806 16382 13858
rect 16434 13806 16446 13858
rect 20626 13806 20638 13858
rect 20690 13806 20702 13858
rect 21298 13806 21310 13858
rect 21362 13806 21374 13858
rect 24322 13806 24334 13858
rect 24386 13806 24398 13858
rect 28018 13806 28030 13858
rect 28082 13806 28094 13858
rect 29474 13806 29486 13858
rect 29538 13806 29550 13858
rect 32162 13806 32174 13858
rect 32226 13806 32238 13858
rect 33058 13806 33070 13858
rect 33122 13806 33134 13858
rect 33730 13806 33742 13858
rect 33794 13806 33806 13858
rect 32510 13794 32562 13806
rect 33406 13794 33458 13806
rect 34078 13794 34130 13806
rect 34526 13858 34578 13870
rect 42478 13858 42530 13870
rect 34850 13806 34862 13858
rect 34914 13806 34926 13858
rect 37426 13806 37438 13858
rect 37490 13806 37502 13858
rect 45378 13806 45390 13858
rect 45442 13806 45454 13858
rect 34526 13794 34578 13806
rect 42478 13794 42530 13806
rect 1934 13746 1986 13758
rect 42814 13746 42866 13758
rect 2594 13694 2606 13746
rect 2658 13694 2670 13746
rect 24546 13694 24558 13746
rect 24610 13694 24622 13746
rect 38434 13694 38446 13746
rect 38498 13694 38510 13746
rect 1934 13682 1986 13694
rect 42814 13682 42866 13694
rect 5854 13634 5906 13646
rect 8430 13634 8482 13646
rect 43262 13634 43314 13646
rect 7970 13582 7982 13634
rect 8034 13582 8046 13634
rect 12562 13582 12574 13634
rect 12626 13582 12638 13634
rect 15362 13582 15374 13634
rect 15426 13582 15438 13634
rect 19618 13582 19630 13634
rect 19682 13582 19694 13634
rect 22418 13582 22430 13634
rect 22482 13582 22494 13634
rect 27122 13582 27134 13634
rect 27186 13582 27198 13634
rect 30594 13582 30606 13634
rect 30658 13582 30670 13634
rect 36194 13582 36206 13634
rect 36258 13582 36270 13634
rect 38546 13582 38558 13634
rect 38610 13582 38622 13634
rect 5854 13570 5906 13582
rect 8430 13570 8482 13582
rect 43262 13570 43314 13582
rect 43822 13634 43874 13646
rect 44258 13582 44270 13634
rect 44322 13582 44334 13634
rect 43822 13570 43874 13582
rect 5630 13522 5682 13534
rect 5630 13458 5682 13470
rect 1344 13354 46592 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 46592 13354
rect 1344 13268 46592 13302
rect 34862 13074 34914 13086
rect 35870 13074 35922 13086
rect 3714 13022 3726 13074
rect 3778 13022 3790 13074
rect 7858 13022 7870 13074
rect 7922 13022 7934 13074
rect 10210 13022 10222 13074
rect 10274 13022 10286 13074
rect 15474 13022 15486 13074
rect 15538 13022 15550 13074
rect 19282 13022 19294 13074
rect 19346 13022 19358 13074
rect 23874 13022 23886 13074
rect 23938 13022 23950 13074
rect 26226 13022 26238 13074
rect 26290 13022 26302 13074
rect 30258 13022 30270 13074
rect 30322 13022 30334 13074
rect 33282 13022 33294 13074
rect 33346 13022 33358 13074
rect 35074 13022 35086 13074
rect 35138 13022 35150 13074
rect 36194 13022 36206 13074
rect 36258 13022 36270 13074
rect 38098 13022 38110 13074
rect 38162 13022 38174 13074
rect 41010 13022 41022 13074
rect 41074 13022 41086 13074
rect 43586 13022 43598 13074
rect 43650 13022 43662 13074
rect 45490 13022 45502 13074
rect 45554 13022 45566 13074
rect 34862 13010 34914 13022
rect 35870 13010 35922 13022
rect 46174 12962 46226 12974
rect 45042 12910 45054 12962
rect 45106 12910 45118 12962
rect 46174 12898 46226 12910
rect 2370 12798 2382 12850
rect 2434 12798 2446 12850
rect 6514 12798 6526 12850
rect 6578 12798 6590 12850
rect 11218 12798 11230 12850
rect 11282 12798 11294 12850
rect 16706 12798 16718 12850
rect 16770 12798 16782 12850
rect 20514 12798 20526 12850
rect 20578 12798 20590 12850
rect 22866 12798 22878 12850
rect 22930 12798 22942 12850
rect 27234 12798 27246 12850
rect 27298 12798 27310 12850
rect 31266 12798 31278 12850
rect 31330 12798 31342 12850
rect 34290 12798 34302 12850
rect 34354 12798 34366 12850
rect 39106 12798 39118 12850
rect 39170 12798 39182 12850
rect 42018 12798 42030 12850
rect 42082 12798 42094 12850
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 43038 12738 43090 12750
rect 43038 12674 43090 12686
rect 44270 12738 44322 12750
rect 44270 12674 44322 12686
rect 1344 12570 46592 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 46592 12570
rect 1344 12484 46592 12518
rect 5630 12402 5682 12414
rect 2258 12350 2270 12402
rect 2322 12350 2334 12402
rect 5630 12338 5682 12350
rect 8082 12238 8094 12290
rect 8146 12238 8158 12290
rect 13010 12238 13022 12290
rect 13074 12238 13086 12290
rect 17938 12238 17950 12290
rect 18002 12238 18014 12290
rect 23986 12238 23998 12290
rect 24050 12238 24062 12290
rect 27570 12238 27582 12290
rect 27634 12238 27646 12290
rect 30370 12238 30382 12290
rect 30434 12238 30446 12290
rect 36418 12238 36430 12290
rect 36482 12238 36494 12290
rect 37314 12238 37326 12290
rect 37378 12238 37390 12290
rect 42914 12238 42926 12290
rect 42978 12238 42990 12290
rect 45938 12238 45950 12290
rect 46002 12238 46014 12290
rect 5070 12178 5122 12190
rect 4610 12126 4622 12178
rect 4674 12126 4686 12178
rect 5070 12114 5122 12126
rect 6962 12014 6974 12066
rect 7026 12014 7038 12066
rect 12002 12014 12014 12066
rect 12066 12014 12078 12066
rect 19058 12014 19070 12066
rect 19122 12014 19134 12066
rect 22978 12014 22990 12066
rect 23042 12014 23054 12066
rect 26562 12014 26574 12066
rect 26626 12014 26638 12066
rect 29362 12014 29374 12066
rect 29426 12014 29438 12066
rect 35074 12014 35086 12066
rect 35138 12014 35150 12066
rect 38658 12014 38670 12066
rect 38722 12014 38734 12066
rect 41906 12014 41918 12066
rect 41970 12014 41982 12066
rect 44706 12014 44718 12066
rect 44770 12014 44782 12066
rect 1598 11954 1650 11966
rect 1598 11890 1650 11902
rect 1344 11786 46592 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 46592 11786
rect 1344 11700 46592 11734
rect 45726 11618 45778 11630
rect 45726 11554 45778 11566
rect 35870 11506 35922 11518
rect 3490 11454 3502 11506
rect 3554 11454 3566 11506
rect 6402 11454 6414 11506
rect 6466 11454 6478 11506
rect 10434 11454 10446 11506
rect 10498 11454 10510 11506
rect 22642 11454 22654 11506
rect 22706 11454 22718 11506
rect 25218 11454 25230 11506
rect 25282 11454 25294 11506
rect 30482 11454 30494 11506
rect 30546 11454 30558 11506
rect 33394 11454 33406 11506
rect 33458 11454 33470 11506
rect 35522 11454 35534 11506
rect 35586 11454 35598 11506
rect 36194 11454 36206 11506
rect 36258 11454 36270 11506
rect 37986 11454 37998 11506
rect 38050 11454 38062 11506
rect 42242 11454 42254 11506
rect 42306 11454 42318 11506
rect 35870 11442 35922 11454
rect 35298 11342 35310 11394
rect 35362 11342 35374 11394
rect 2370 11230 2382 11282
rect 2434 11230 2446 11282
rect 7746 11230 7758 11282
rect 7810 11230 7822 11282
rect 9314 11230 9326 11282
rect 9378 11230 9390 11282
rect 21522 11230 21534 11282
rect 21586 11230 21598 11282
rect 26562 11230 26574 11282
rect 26626 11230 26638 11282
rect 29362 11230 29374 11282
rect 29426 11230 29438 11282
rect 34402 11230 34414 11282
rect 34466 11230 34478 11282
rect 39218 11230 39230 11282
rect 39282 11230 39294 11282
rect 43250 11230 43262 11282
rect 43314 11230 43326 11282
rect 44942 11170 44994 11182
rect 44942 11106 44994 11118
rect 1344 11002 46592 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 46592 11002
rect 1344 10916 46592 10950
rect 44830 10834 44882 10846
rect 4498 10782 4510 10834
rect 4562 10782 4574 10834
rect 44830 10770 44882 10782
rect 45726 10722 45778 10734
rect 6738 10670 6750 10722
rect 6802 10670 6814 10722
rect 11778 10670 11790 10722
rect 11842 10670 11854 10722
rect 27906 10670 27918 10722
rect 27970 10670 27982 10722
rect 35410 10670 35422 10722
rect 35474 10670 35486 10722
rect 38658 10670 38670 10722
rect 38722 10670 38734 10722
rect 43922 10670 43934 10722
rect 43986 10670 43998 10722
rect 45726 10658 45778 10670
rect 1822 10610 1874 10622
rect 46062 10610 46114 10622
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 1822 10546 1874 10558
rect 46062 10546 46114 10558
rect 45502 10498 45554 10510
rect 5954 10446 5966 10498
rect 6018 10446 6030 10498
rect 10546 10446 10558 10498
rect 10610 10446 10622 10498
rect 26562 10446 26574 10498
rect 26626 10446 26638 10498
rect 34402 10446 34414 10498
rect 34466 10446 34478 10498
rect 37426 10446 37438 10498
rect 37490 10446 37502 10498
rect 42914 10446 42926 10498
rect 42978 10446 42990 10498
rect 45502 10434 45554 10446
rect 5294 10386 5346 10398
rect 5294 10322 5346 10334
rect 1344 10218 46592 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 46592 10218
rect 1344 10132 46592 10166
rect 5854 9938 5906 9950
rect 10546 9886 10558 9938
rect 10610 9886 10622 9938
rect 32722 9886 32734 9938
rect 32786 9886 32798 9938
rect 38322 9886 38334 9938
rect 38386 9886 38398 9938
rect 41122 9886 41134 9938
rect 41186 9886 41198 9938
rect 45378 9886 45390 9938
rect 45442 9886 45454 9938
rect 5854 9874 5906 9886
rect 44034 9774 44046 9826
rect 44098 9774 44110 9826
rect 43598 9714 43650 9726
rect 9202 9662 9214 9714
rect 9266 9662 9278 9714
rect 33954 9662 33966 9714
rect 34018 9662 34030 9714
rect 39330 9662 39342 9714
rect 39394 9662 39406 9714
rect 42130 9662 42142 9714
rect 42194 9662 42206 9714
rect 43598 9650 43650 9662
rect 43262 9602 43314 9614
rect 43262 9538 43314 9550
rect 44270 9602 44322 9614
rect 44270 9538 44322 9550
rect 44942 9602 44994 9614
rect 44942 9538 44994 9550
rect 1344 9434 46592 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 46592 9434
rect 1344 9348 46592 9382
rect 43934 9266 43986 9278
rect 43934 9202 43986 9214
rect 35634 9102 35646 9154
rect 35698 9102 35710 9154
rect 41010 9102 41022 9154
rect 41074 9102 41086 9154
rect 46050 9102 46062 9154
rect 46114 9102 46126 9154
rect 34738 8878 34750 8930
rect 34802 8878 34814 8930
rect 42130 8878 42142 8930
rect 42194 8878 42206 8930
rect 44706 8878 44718 8930
rect 44770 8878 44782 8930
rect 1344 8650 46592 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 46592 8650
rect 1344 8564 46592 8598
rect 40226 8318 40238 8370
rect 40290 8318 40302 8370
rect 45602 8318 45614 8370
rect 45666 8318 45678 8370
rect 2818 8206 2830 8258
rect 2882 8206 2894 8258
rect 44270 8146 44322 8158
rect 2034 8094 2046 8146
rect 2098 8094 2110 8146
rect 41234 8094 41246 8146
rect 41298 8094 41310 8146
rect 44270 8082 44322 8094
rect 3390 8034 3442 8046
rect 3390 7970 3442 7982
rect 43934 8034 43986 8046
rect 43934 7970 43986 7982
rect 44942 8034 44994 8046
rect 44942 7970 44994 7982
rect 1344 7866 46592 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 46592 7866
rect 1344 7780 46592 7814
rect 44606 7698 44658 7710
rect 44606 7634 44658 7646
rect 42354 7534 42366 7586
rect 42418 7534 42430 7586
rect 46050 7534 46062 7586
rect 46114 7534 46126 7586
rect 2930 7422 2942 7474
rect 2994 7422 3006 7474
rect 44930 7422 44942 7474
rect 44994 7422 45006 7474
rect 3502 7362 3554 7374
rect 1922 7310 1934 7362
rect 1986 7310 1998 7362
rect 41458 7310 41470 7362
rect 41522 7310 41534 7362
rect 3502 7298 3554 7310
rect 1344 7082 46592 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 46592 7082
rect 1344 6996 46592 7030
rect 41906 6750 41918 6802
rect 41970 6750 41982 6802
rect 45726 6690 45778 6702
rect 2930 6638 2942 6690
rect 2994 6638 3006 6690
rect 45726 6626 45778 6638
rect 2034 6526 2046 6578
rect 2098 6526 2110 6578
rect 42802 6526 42814 6578
rect 42866 6526 42878 6578
rect 44942 6466 44994 6478
rect 44942 6402 44994 6414
rect 1344 6298 46592 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 46592 6298
rect 1344 6212 46592 6246
rect 22206 6130 22258 6142
rect 22206 6066 22258 6078
rect 24446 6130 24498 6142
rect 24446 6066 24498 6078
rect 33406 6130 33458 6142
rect 33406 6066 33458 6078
rect 33854 6130 33906 6142
rect 33854 6066 33906 6078
rect 20750 6018 20802 6030
rect 20750 5954 20802 5966
rect 22990 6018 23042 6030
rect 22990 5954 23042 5966
rect 23662 6018 23714 6030
rect 23662 5954 23714 5966
rect 26462 6018 26514 6030
rect 45938 5966 45950 6018
rect 46002 5966 46014 6018
rect 26462 5954 26514 5966
rect 23998 5906 24050 5918
rect 33070 5906 33122 5918
rect 2930 5854 2942 5906
rect 2994 5854 3006 5906
rect 20962 5854 20974 5906
rect 21026 5854 21038 5906
rect 22418 5854 22430 5906
rect 22482 5854 22494 5906
rect 23202 5854 23214 5906
rect 23266 5854 23278 5906
rect 26226 5854 26238 5906
rect 26290 5854 26302 5906
rect 23998 5842 24050 5854
rect 33070 5842 33122 5854
rect 20414 5794 20466 5806
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 20414 5730 20466 5742
rect 28814 5794 28866 5806
rect 44930 5742 44942 5794
rect 44994 5742 45006 5794
rect 28814 5730 28866 5742
rect 1344 5514 46592 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 46592 5514
rect 1344 5428 46592 5462
rect 46174 5234 46226 5246
rect 24882 5182 24894 5234
rect 24946 5182 24958 5234
rect 45602 5182 45614 5234
rect 45666 5182 45678 5234
rect 46174 5170 46226 5182
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 2494 5122 2546 5134
rect 14702 5122 14754 5134
rect 13682 5070 13694 5122
rect 13746 5070 13758 5122
rect 2494 5058 2546 5070
rect 14702 5058 14754 5070
rect 15598 5122 15650 5134
rect 15598 5058 15650 5070
rect 16942 5122 16994 5134
rect 18062 5122 18114 5134
rect 19742 5122 19794 5134
rect 17490 5070 17502 5122
rect 17554 5070 17566 5122
rect 18610 5070 18622 5122
rect 18674 5070 18686 5122
rect 16942 5058 16994 5070
rect 18062 5058 18114 5070
rect 19742 5058 19794 5070
rect 22766 5122 22818 5134
rect 22766 5058 22818 5070
rect 23102 5122 23154 5134
rect 24446 5122 24498 5134
rect 41694 5122 41746 5134
rect 44942 5122 44994 5134
rect 23874 5070 23886 5122
rect 23938 5070 23950 5122
rect 26114 5070 26126 5122
rect 26178 5070 26190 5122
rect 28242 5070 28254 5122
rect 28306 5070 28318 5122
rect 29362 5070 29374 5122
rect 29426 5070 29438 5122
rect 30034 5070 30046 5122
rect 30098 5070 30110 5122
rect 31266 5070 31278 5122
rect 31330 5070 31342 5122
rect 31938 5070 31950 5122
rect 32002 5070 32014 5122
rect 32610 5070 32622 5122
rect 32674 5070 32686 5122
rect 33282 5070 33294 5122
rect 33346 5070 33358 5122
rect 33954 5070 33966 5122
rect 34018 5070 34030 5122
rect 37650 5070 37662 5122
rect 37714 5070 37726 5122
rect 38322 5070 38334 5122
rect 38386 5070 38398 5122
rect 39106 5070 39118 5122
rect 39170 5070 39182 5122
rect 40114 5070 40126 5122
rect 40178 5070 40190 5122
rect 44034 5070 44046 5122
rect 44098 5070 44110 5122
rect 23102 5058 23154 5070
rect 24446 5058 24498 5070
rect 41694 5058 41746 5070
rect 44942 5058 44994 5070
rect 2046 5010 2098 5022
rect 2046 4946 2098 4958
rect 12238 5010 12290 5022
rect 12238 4946 12290 4958
rect 16606 5010 16658 5022
rect 16606 4946 16658 4958
rect 17278 5010 17330 5022
rect 17278 4946 17330 4958
rect 18398 5010 18450 5022
rect 18398 4946 18450 4958
rect 20414 5010 20466 5022
rect 20414 4946 20466 4958
rect 21758 5010 21810 5022
rect 21758 4946 21810 4958
rect 22430 5010 22482 5022
rect 22430 4946 22482 4958
rect 23438 5010 23490 5022
rect 23438 4946 23490 4958
rect 24110 5010 24162 5022
rect 24110 4946 24162 4958
rect 26686 5010 26738 5022
rect 26686 4946 26738 4958
rect 27022 5010 27074 5022
rect 27022 4946 27074 4958
rect 28478 5010 28530 5022
rect 28478 4946 28530 4958
rect 30270 5010 30322 5022
rect 30270 4946 30322 4958
rect 32846 5010 32898 5022
rect 32846 4946 32898 4958
rect 38558 5010 38610 5022
rect 38558 4946 38610 4958
rect 40350 5010 40402 5022
rect 40350 4946 40402 4958
rect 44270 5010 44322 5022
rect 44270 4946 44322 4958
rect 9438 4898 9490 4910
rect 9438 4834 9490 4846
rect 12574 4898 12626 4910
rect 12574 4834 12626 4846
rect 13470 4898 13522 4910
rect 13470 4834 13522 4846
rect 15038 4898 15090 4910
rect 15038 4834 15090 4846
rect 15934 4898 15986 4910
rect 15934 4834 15986 4846
rect 19518 4898 19570 4910
rect 19518 4834 19570 4846
rect 20078 4898 20130 4910
rect 20078 4834 20130 4846
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 22094 4898 22146 4910
rect 22094 4834 22146 4846
rect 26350 4898 26402 4910
rect 26350 4834 26402 4846
rect 29598 4898 29650 4910
rect 29598 4834 29650 4846
rect 30942 4898 30994 4910
rect 30942 4834 30994 4846
rect 31502 4898 31554 4910
rect 31502 4834 31554 4846
rect 32174 4898 32226 4910
rect 32174 4834 32226 4846
rect 33518 4898 33570 4910
rect 33518 4834 33570 4846
rect 34190 4898 34242 4910
rect 34190 4834 34242 4846
rect 34750 4898 34802 4910
rect 34750 4834 34802 4846
rect 35646 4898 35698 4910
rect 35646 4834 35698 4846
rect 37886 4898 37938 4910
rect 37886 4834 37938 4846
rect 39342 4898 39394 4910
rect 39342 4834 39394 4846
rect 40910 4898 40962 4910
rect 40910 4834 40962 4846
rect 43598 4898 43650 4910
rect 43598 4834 43650 4846
rect 1344 4730 46592 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 46592 4730
rect 1344 4644 46592 4678
rect 2046 4562 2098 4574
rect 2046 4498 2098 4510
rect 8878 4562 8930 4574
rect 8878 4498 8930 4510
rect 9998 4562 10050 4574
rect 9998 4498 10050 4510
rect 14702 4562 14754 4574
rect 14702 4498 14754 4510
rect 15038 4562 15090 4574
rect 15038 4498 15090 4510
rect 17726 4562 17778 4574
rect 17726 4498 17778 4510
rect 19406 4562 19458 4574
rect 19406 4498 19458 4510
rect 21086 4562 21138 4574
rect 21086 4498 21138 4510
rect 22654 4562 22706 4574
rect 22654 4498 22706 4510
rect 26462 4562 26514 4574
rect 26462 4498 26514 4510
rect 28030 4562 28082 4574
rect 28030 4498 28082 4510
rect 30494 4562 30546 4574
rect 30494 4498 30546 4510
rect 32174 4562 32226 4574
rect 32174 4498 32226 4510
rect 33406 4562 33458 4574
rect 33406 4498 33458 4510
rect 34078 4562 34130 4574
rect 34078 4498 34130 4510
rect 35422 4562 35474 4574
rect 35422 4498 35474 4510
rect 37214 4562 37266 4574
rect 37214 4498 37266 4510
rect 39902 4562 39954 4574
rect 39902 4498 39954 4510
rect 40910 4562 40962 4574
rect 40910 4498 40962 4510
rect 44718 4562 44770 4574
rect 44718 4498 44770 4510
rect 46174 4562 46226 4574
rect 46174 4498 46226 4510
rect 10334 4450 10386 4462
rect 10334 4386 10386 4398
rect 18398 4450 18450 4462
rect 18398 4386 18450 4398
rect 19742 4450 19794 4462
rect 19742 4386 19794 4398
rect 20078 4450 20130 4462
rect 20078 4386 20130 4398
rect 23326 4450 23378 4462
rect 23326 4386 23378 4398
rect 24446 4450 24498 4462
rect 24446 4386 24498 4398
rect 29150 4450 29202 4462
rect 29150 4386 29202 4398
rect 31166 4450 31218 4462
rect 31166 4386 31218 4398
rect 34526 4450 34578 4462
rect 34526 4386 34578 4398
rect 35870 4450 35922 4462
rect 35870 4386 35922 4398
rect 41918 4450 41970 4462
rect 41918 4386 41970 4398
rect 43598 4450 43650 4462
rect 43598 4386 43650 4398
rect 44046 4450 44098 4462
rect 44046 4386 44098 4398
rect 45166 4450 45218 4462
rect 45166 4386 45218 4398
rect 45502 4450 45554 4462
rect 45502 4386 45554 4398
rect 45838 4450 45890 4462
rect 45838 4386 45890 4398
rect 1710 4338 1762 4350
rect 1710 4274 1762 4286
rect 9662 4338 9714 4350
rect 14366 4338 14418 4350
rect 13010 4286 13022 4338
rect 13074 4286 13086 4338
rect 9662 4274 9714 4286
rect 14366 4274 14418 4286
rect 17390 4338 17442 4350
rect 17390 4274 17442 4286
rect 19070 4338 19122 4350
rect 31838 4338 31890 4350
rect 34862 4338 34914 4350
rect 22866 4286 22878 4338
rect 22930 4286 22942 4338
rect 23538 4286 23550 4338
rect 23602 4286 23614 4338
rect 24210 4286 24222 4338
rect 24274 4286 24286 4338
rect 28242 4286 28254 4338
rect 28306 4286 28318 4338
rect 30706 4286 30718 4338
rect 30770 4286 30782 4338
rect 31378 4286 31390 4338
rect 31442 4286 31454 4338
rect 33170 4286 33182 4338
rect 33234 4286 33246 4338
rect 33842 4286 33854 4338
rect 33906 4286 33918 4338
rect 36082 4286 36094 4338
rect 36146 4286 36158 4338
rect 40114 4286 40126 4338
rect 40178 4286 40190 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 42130 4286 42142 4338
rect 42194 4286 42206 4338
rect 44482 4286 44494 4338
rect 44546 4286 44558 4338
rect 19070 4274 19122 4286
rect 31838 4274 31890 4286
rect 34862 4274 34914 4286
rect 2494 4226 2546 4238
rect 2494 4162 2546 4174
rect 11454 4226 11506 4238
rect 11454 4162 11506 4174
rect 12014 4226 12066 4238
rect 12014 4162 12066 4174
rect 13582 4226 13634 4238
rect 13582 4162 13634 4174
rect 14142 4226 14194 4238
rect 16830 4226 16882 4238
rect 22318 4226 22370 4238
rect 15474 4174 15486 4226
rect 15538 4174 15550 4226
rect 21522 4174 21534 4226
rect 21586 4174 21598 4226
rect 14142 4162 14194 4174
rect 16830 4162 16882 4174
rect 22318 4162 22370 4174
rect 26238 4226 26290 4238
rect 26238 4162 26290 4174
rect 27694 4226 27746 4238
rect 27694 4162 27746 4174
rect 30270 4226 30322 4238
rect 30270 4162 30322 4174
rect 36654 4226 36706 4238
rect 38558 4226 38610 4238
rect 37650 4174 37662 4226
rect 37714 4174 37726 4226
rect 36654 4162 36706 4174
rect 38558 4162 38610 4174
rect 39678 4226 39730 4238
rect 39678 4162 39730 4174
rect 8094 4114 8146 4126
rect 12350 4114 12402 4126
rect 11554 4062 11566 4114
rect 11618 4111 11630 4114
rect 12002 4111 12014 4114
rect 11618 4065 12014 4111
rect 11618 4062 11630 4065
rect 12002 4062 12014 4065
rect 12066 4062 12078 4114
rect 8094 4050 8146 4062
rect 12350 4050 12402 4062
rect 27246 4114 27298 4126
rect 27246 4050 27298 4062
rect 1344 3946 46592 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 46592 3946
rect 1344 3860 46592 3894
rect 19070 3666 19122 3678
rect 23214 3666 23266 3678
rect 42702 3666 42754 3678
rect 19730 3614 19742 3666
rect 19794 3614 19806 3666
rect 25554 3614 25566 3666
rect 25618 3614 25630 3666
rect 30482 3614 30494 3666
rect 30546 3614 30558 3666
rect 32946 3614 32958 3666
rect 33010 3614 33022 3666
rect 36978 3614 36990 3666
rect 37042 3614 37054 3666
rect 40226 3614 40238 3666
rect 40290 3614 40302 3666
rect 41794 3614 41806 3666
rect 41858 3614 41870 3666
rect 19070 3602 19122 3614
rect 23214 3602 23266 3614
rect 42702 3602 42754 3614
rect 8766 3554 8818 3566
rect 8766 3490 8818 3502
rect 10558 3554 10610 3566
rect 10558 3490 10610 3502
rect 12238 3554 12290 3566
rect 20190 3554 20242 3566
rect 25118 3554 25170 3566
rect 13794 3502 13806 3554
rect 13858 3502 13870 3554
rect 16258 3502 16270 3554
rect 16322 3502 16334 3554
rect 18498 3502 18510 3554
rect 18562 3502 18574 3554
rect 21186 3502 21198 3554
rect 21250 3502 21262 3554
rect 22418 3502 22430 3554
rect 22482 3502 22494 3554
rect 12238 3490 12290 3502
rect 20190 3490 20242 3502
rect 25118 3490 25170 3502
rect 26462 3554 26514 3566
rect 27694 3554 27746 3566
rect 30046 3554 30098 3566
rect 26898 3502 26910 3554
rect 26962 3502 26974 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 26462 3490 26514 3502
rect 27694 3490 27746 3502
rect 30046 3490 30098 3502
rect 32510 3554 32562 3566
rect 36542 3554 36594 3566
rect 34290 3502 34302 3554
rect 34354 3502 34366 3554
rect 34962 3502 34974 3554
rect 35026 3502 35038 3554
rect 32510 3490 32562 3502
rect 36542 3490 36594 3502
rect 39790 3554 39842 3566
rect 39790 3490 39842 3502
rect 41358 3554 41410 3566
rect 46050 3502 46062 3554
rect 46114 3502 46126 3554
rect 41358 3490 41410 3502
rect 1710 3442 1762 3454
rect 1710 3378 1762 3390
rect 2046 3442 2098 3454
rect 2046 3378 2098 3390
rect 2942 3442 2994 3454
rect 2942 3378 2994 3390
rect 6862 3442 6914 3454
rect 6862 3378 6914 3390
rect 7198 3442 7250 3454
rect 7198 3378 7250 3390
rect 7646 3442 7698 3454
rect 7646 3378 7698 3390
rect 10894 3442 10946 3454
rect 10894 3378 10946 3390
rect 11566 3442 11618 3454
rect 11566 3378 11618 3390
rect 12574 3442 12626 3454
rect 12574 3378 12626 3390
rect 21422 3442 21474 3454
rect 21422 3378 21474 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 24670 3442 24722 3454
rect 24670 3378 24722 3390
rect 26686 3442 26738 3454
rect 26686 3378 26738 3390
rect 27358 3442 27410 3454
rect 27358 3378 27410 3390
rect 29262 3442 29314 3454
rect 29262 3378 29314 3390
rect 31614 3442 31666 3454
rect 31614 3378 31666 3390
rect 33854 3442 33906 3454
rect 33854 3378 33906 3390
rect 34078 3442 34130 3454
rect 34078 3378 34130 3390
rect 34750 3442 34802 3454
rect 34750 3378 34802 3390
rect 37886 3442 37938 3454
rect 37886 3378 37938 3390
rect 38110 3442 38162 3454
rect 38110 3378 38162 3390
rect 38446 3442 38498 3454
rect 38446 3378 38498 3390
rect 38782 3442 38834 3454
rect 38782 3378 38834 3390
rect 39118 3442 39170 3454
rect 39118 3378 39170 3390
rect 45838 3442 45890 3454
rect 45838 3378 45890 3390
rect 2382 3330 2434 3342
rect 2382 3266 2434 3278
rect 7982 3330 8034 3342
rect 7982 3266 8034 3278
rect 9774 3330 9826 3342
rect 9774 3266 9826 3278
rect 11230 3330 11282 3342
rect 11230 3266 11282 3278
rect 11902 3330 11954 3342
rect 11902 3266 11954 3278
rect 13134 3330 13186 3342
rect 13134 3266 13186 3278
rect 15598 3330 15650 3342
rect 15598 3266 15650 3278
rect 17838 3330 17890 3342
rect 17838 3266 17890 3278
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 43038 3330 43090 3342
rect 43038 3266 43090 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 44382 3330 44434 3342
rect 44382 3266 44434 3278
rect 44830 3330 44882 3342
rect 44830 3266 44882 3278
rect 45278 3330 45330 3342
rect 45278 3266 45330 3278
rect 1344 3162 46592 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 46592 3162
rect 1344 3076 46592 3110
rect 43922 2382 43934 2434
rect 43986 2431 43998 2434
rect 45266 2431 45278 2434
rect 43986 2385 45278 2431
rect 43986 2382 43998 2385
rect 45266 2382 45278 2385
rect 45330 2382 45342 2434
rect 8866 926 8878 978
rect 8930 975 8942 978
rect 9762 975 9774 978
rect 8930 929 9774 975
rect 8930 926 8942 929
rect 9762 926 9774 929
rect 9826 926 9838 978
<< via1 >>
rect 32286 45166 32338 45218
rect 33406 45166 33458 45218
rect 14142 44830 14194 44882
rect 14926 44830 14978 44882
rect 16830 44830 16882 44882
rect 17502 44830 17554 44882
rect 20190 44830 20242 44882
rect 20974 44830 21026 44882
rect 26910 44830 26962 44882
rect 27582 44830 27634 44882
rect 28926 44830 28978 44882
rect 30046 44830 30098 44882
rect 36990 44830 37042 44882
rect 38110 44830 38162 44882
rect 40350 44830 40402 44882
rect 41918 44830 41970 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 17502 44494 17554 44546
rect 25566 44494 25618 44546
rect 7422 44382 7474 44434
rect 9774 44382 9826 44434
rect 13470 44382 13522 44434
rect 14926 44382 14978 44434
rect 19518 44382 19570 44434
rect 20974 44382 21026 44434
rect 23438 44382 23490 44434
rect 25342 44382 25394 44434
rect 28814 44382 28866 44434
rect 30382 44382 30434 44434
rect 32622 44382 32674 44434
rect 33406 44382 33458 44434
rect 36766 44382 36818 44434
rect 37102 44382 37154 44434
rect 40350 44382 40402 44434
rect 41918 44382 41970 44434
rect 44046 44382 44098 44434
rect 7870 44270 7922 44322
rect 13694 44270 13746 44322
rect 20190 44270 20242 44322
rect 21982 44270 22034 44322
rect 23886 44270 23938 44322
rect 26238 44270 26290 44322
rect 26910 44270 26962 44322
rect 27582 44270 27634 44322
rect 33966 44270 34018 44322
rect 34526 44270 34578 44322
rect 37662 44270 37714 44322
rect 38110 44270 38162 44322
rect 38782 44270 38834 44322
rect 43710 44270 43762 44322
rect 15934 44158 15986 44210
rect 35982 44158 36034 44210
rect 46174 44158 46226 44210
rect 7646 44046 7698 44098
rect 9326 44046 9378 44098
rect 14030 44046 14082 44098
rect 14366 44046 14418 44098
rect 18286 44046 18338 44098
rect 26686 44046 26738 44098
rect 27358 44046 27410 44098
rect 28366 44046 28418 44098
rect 29934 44046 29986 44098
rect 32174 44046 32226 44098
rect 33742 44046 33794 44098
rect 34862 44046 34914 44098
rect 38446 44046 38498 44098
rect 39118 44046 39170 44098
rect 39790 44046 39842 44098
rect 41358 44046 41410 44098
rect 45614 44046 45666 44098
rect 45838 44046 45890 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 17726 43710 17778 43762
rect 27694 43710 27746 43762
rect 30046 43710 30098 43762
rect 34302 43710 34354 43762
rect 37886 43710 37938 43762
rect 18734 43598 18786 43650
rect 19070 43598 19122 43650
rect 20414 43598 20466 43650
rect 21086 43598 21138 43650
rect 21422 43598 21474 43650
rect 21758 43598 21810 43650
rect 23998 43598 24050 43650
rect 25230 43598 25282 43650
rect 25566 43598 25618 43650
rect 30494 43598 30546 43650
rect 31614 43598 31666 43650
rect 31838 43598 31890 43650
rect 34974 43598 35026 43650
rect 35198 43598 35250 43650
rect 35534 43598 35586 43650
rect 38334 43598 38386 43650
rect 39678 43598 39730 43650
rect 39902 43598 39954 43650
rect 40238 43598 40290 43650
rect 42590 43598 42642 43650
rect 42814 43598 42866 43650
rect 18398 43486 18450 43538
rect 19294 43486 19346 43538
rect 19854 43486 19906 43538
rect 20862 43486 20914 43538
rect 22094 43486 22146 43538
rect 22430 43486 22482 43538
rect 23774 43486 23826 43538
rect 24334 43486 24386 43538
rect 26462 43486 26514 43538
rect 28478 43486 28530 43538
rect 29822 43486 29874 43538
rect 30718 43486 30770 43538
rect 32062 43486 32114 43538
rect 39006 43486 39058 43538
rect 41246 43486 41298 43538
rect 43038 43486 43090 43538
rect 45054 43486 45106 43538
rect 22878 43374 22930 43426
rect 26910 43374 26962 43426
rect 28926 43374 28978 43426
rect 41694 43374 41746 43426
rect 46062 43374 46114 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 45726 42926 45778 42978
rect 18174 42814 18226 42866
rect 25006 42814 25058 42866
rect 7534 42702 7586 42754
rect 13918 42702 13970 42754
rect 19070 42702 19122 42754
rect 20638 42702 20690 42754
rect 21646 42702 21698 42754
rect 22430 42702 22482 42754
rect 23326 42702 23378 42754
rect 25566 42702 25618 42754
rect 26574 42702 26626 42754
rect 38222 42702 38274 42754
rect 39006 42702 39058 42754
rect 39678 42702 39730 42754
rect 40238 42702 40290 42754
rect 44046 42702 44098 42754
rect 7758 42590 7810 42642
rect 14142 42590 14194 42642
rect 18846 42590 18898 42642
rect 20414 42590 20466 42642
rect 22206 42590 22258 42642
rect 23550 42590 23602 42642
rect 25902 42590 25954 42642
rect 26238 42590 26290 42642
rect 38558 42590 38610 42642
rect 39230 42590 39282 42642
rect 39902 42590 39954 42642
rect 40574 42590 40626 42642
rect 1710 42478 1762 42530
rect 21870 42478 21922 42530
rect 44270 42478 44322 42530
rect 44942 42478 44994 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 27134 42142 27186 42194
rect 27806 42142 27858 42194
rect 28142 42142 28194 42194
rect 30494 42142 30546 42194
rect 37438 42142 37490 42194
rect 38782 42142 38834 42194
rect 28478 42030 28530 42082
rect 38446 42030 38498 42082
rect 44158 42030 44210 42082
rect 26910 41918 26962 41970
rect 27582 41918 27634 41970
rect 30270 41918 30322 41970
rect 37102 41918 37154 41970
rect 44942 41806 44994 41858
rect 46286 41806 46338 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 44830 41022 44882 41074
rect 45166 41022 45218 41074
rect 45838 41022 45890 41074
rect 46174 41022 46226 41074
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 46062 40574 46114 40626
rect 45390 40462 45442 40514
rect 44158 40238 44210 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 43038 39678 43090 39730
rect 42254 39454 42306 39506
rect 46174 39454 46226 39506
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 43262 38894 43314 38946
rect 45726 38894 45778 38946
rect 41918 38670 41970 38722
rect 44718 38670 44770 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 17838 38110 17890 38162
rect 41358 38110 41410 38162
rect 18846 37886 18898 37938
rect 42366 37886 42418 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 13806 37326 13858 37378
rect 17502 37326 17554 37378
rect 38110 37326 38162 37378
rect 43822 37326 43874 37378
rect 15150 37102 15202 37154
rect 18622 37102 18674 37154
rect 39230 37102 39282 37154
rect 42478 37102 42530 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 14814 36542 14866 36594
rect 18734 36542 18786 36594
rect 22430 36542 22482 36594
rect 38558 36542 38610 36594
rect 40910 36542 40962 36594
rect 15822 36318 15874 36370
rect 19742 36318 19794 36370
rect 23550 36318 23602 36370
rect 37438 36318 37490 36370
rect 41918 36318 41970 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 42478 35870 42530 35922
rect 6190 35758 6242 35810
rect 16046 35758 16098 35810
rect 19518 35758 19570 35810
rect 22654 35758 22706 35810
rect 39902 35758 39954 35810
rect 41694 35646 41746 35698
rect 44942 35646 44994 35698
rect 45390 35646 45442 35698
rect 5182 35534 5234 35586
rect 14702 35534 14754 35586
rect 16494 35534 16546 35586
rect 16830 35534 16882 35586
rect 20638 35534 20690 35586
rect 23662 35534 23714 35586
rect 38894 35534 38946 35586
rect 41806 35422 41858 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 8654 34974 8706 35026
rect 11454 34974 11506 35026
rect 14702 34974 14754 35026
rect 17614 34974 17666 35026
rect 22318 34974 22370 35026
rect 25118 34974 25170 35026
rect 32622 34974 32674 35026
rect 38110 34974 38162 35026
rect 40798 34974 40850 35026
rect 7310 34750 7362 34802
rect 12686 34750 12738 34802
rect 15934 34750 15986 34802
rect 18510 34750 18562 34802
rect 23550 34750 23602 34802
rect 26126 34750 26178 34802
rect 31502 34750 31554 34802
rect 39006 34750 39058 34802
rect 42142 34750 42194 34802
rect 16606 34638 16658 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 1710 34302 1762 34354
rect 2270 34302 2322 34354
rect 44942 34302 44994 34354
rect 45502 34302 45554 34354
rect 8542 34190 8594 34242
rect 13582 34190 13634 34242
rect 15710 34190 15762 34242
rect 19742 34190 19794 34242
rect 21534 34190 21586 34242
rect 27246 34190 27298 34242
rect 30270 34190 30322 34242
rect 33406 34190 33458 34242
rect 37326 34190 37378 34242
rect 4846 34078 4898 34130
rect 5406 34078 5458 34130
rect 41806 34078 41858 34130
rect 42366 34078 42418 34130
rect 5854 33966 5906 34018
rect 7534 33966 7586 34018
rect 11342 33966 11394 34018
rect 12350 33966 12402 34018
rect 12574 33966 12626 34018
rect 14366 33966 14418 34018
rect 17502 33966 17554 34018
rect 17950 33966 18002 34018
rect 18398 33966 18450 34018
rect 22654 33966 22706 34018
rect 26238 33966 26290 34018
rect 29038 33966 29090 34018
rect 30830 33966 30882 34018
rect 31054 33966 31106 34018
rect 34526 33966 34578 34018
rect 38670 33966 38722 34018
rect 40350 33966 40402 34018
rect 41246 33966 41298 34018
rect 41246 33854 41298 33906
rect 41694 33854 41746 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 12350 33518 12402 33570
rect 12910 33518 12962 33570
rect 17054 33518 17106 33570
rect 44382 33518 44434 33570
rect 3614 33406 3666 33458
rect 8878 33406 8930 33458
rect 11902 33406 11954 33458
rect 19518 33406 19570 33458
rect 24670 33406 24722 33458
rect 30158 33406 30210 33458
rect 33182 33406 33234 33458
rect 37998 33406 38050 33458
rect 13358 33294 13410 33346
rect 14030 33294 14082 33346
rect 40686 33294 40738 33346
rect 41358 33294 41410 33346
rect 4958 33182 5010 33234
rect 9662 33182 9714 33234
rect 10894 33182 10946 33234
rect 17390 33182 17442 33234
rect 17726 33182 17778 33234
rect 18398 33182 18450 33234
rect 21646 33182 21698 33234
rect 22990 33182 23042 33234
rect 23326 33182 23378 33234
rect 25678 33182 25730 33234
rect 28254 33182 28306 33234
rect 31166 33182 31218 33234
rect 34078 33182 34130 33234
rect 39006 33182 39058 33234
rect 6190 33070 6242 33122
rect 12350 33070 12402 33122
rect 12910 33070 12962 33122
rect 16494 33070 16546 33122
rect 21534 33070 21586 33122
rect 28366 33070 28418 33122
rect 40014 33070 40066 33122
rect 40462 33070 40514 33122
rect 43598 33070 43650 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 5518 32734 5570 32786
rect 6078 32734 6130 32786
rect 13246 32734 13298 32786
rect 17502 32734 17554 32786
rect 23774 32734 23826 32786
rect 24334 32734 24386 32786
rect 29710 32734 29762 32786
rect 30270 32734 30322 32786
rect 44494 32734 44546 32786
rect 45166 32734 45218 32786
rect 6974 32622 7026 32674
rect 9438 32622 9490 32674
rect 10222 32622 10274 32674
rect 14030 32622 14082 32674
rect 18174 32622 18226 32674
rect 30494 32622 30546 32674
rect 33854 32622 33906 32674
rect 38782 32622 38834 32674
rect 2382 32510 2434 32562
rect 2942 32510 2994 32562
rect 12462 32510 12514 32562
rect 13134 32510 13186 32562
rect 16382 32510 16434 32562
rect 16942 32510 16994 32562
rect 20638 32510 20690 32562
rect 21310 32510 21362 32562
rect 26574 32510 26626 32562
rect 27246 32510 27298 32562
rect 30718 32510 30770 32562
rect 31390 32510 31442 32562
rect 31838 32510 31890 32562
rect 33294 32510 33346 32562
rect 41022 32510 41074 32562
rect 41694 32510 41746 32562
rect 42030 32510 42082 32562
rect 7982 32398 8034 32450
rect 8990 32398 9042 32450
rect 19182 32398 19234 32450
rect 31166 32398 31218 32450
rect 32174 32398 32226 32450
rect 33070 32398 33122 32450
rect 35198 32398 35250 32450
rect 37662 32398 37714 32450
rect 39678 32398 39730 32450
rect 40014 32398 40066 32450
rect 40238 32398 40290 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 17054 31950 17106 32002
rect 3502 31838 3554 31890
rect 5518 31838 5570 31890
rect 13022 31838 13074 31890
rect 20862 31838 20914 31890
rect 21198 31838 21250 31890
rect 28702 31838 28754 31890
rect 29038 31838 29090 31890
rect 33966 31838 34018 31890
rect 35758 31838 35810 31890
rect 42590 31838 42642 31890
rect 8654 31726 8706 31778
rect 9214 31726 9266 31778
rect 9550 31726 9602 31778
rect 9998 31726 10050 31778
rect 13358 31726 13410 31778
rect 13918 31726 13970 31778
rect 17166 31726 17218 31778
rect 17838 31726 17890 31778
rect 24222 31726 24274 31778
rect 24782 31726 24834 31778
rect 25230 31726 25282 31778
rect 25678 31726 25730 31778
rect 32062 31726 32114 31778
rect 32510 31726 32562 31778
rect 39118 31726 39170 31778
rect 39454 31726 39506 31778
rect 43038 31726 43090 31778
rect 2382 31614 2434 31666
rect 21982 31614 22034 31666
rect 29822 31614 29874 31666
rect 34974 31614 35026 31666
rect 42814 31614 42866 31666
rect 43710 31614 43762 31666
rect 6078 31502 6130 31554
rect 12350 31502 12402 31554
rect 16494 31502 16546 31554
rect 20302 31502 20354 31554
rect 28142 31502 28194 31554
rect 35870 31502 35922 31554
rect 37102 31502 37154 31554
rect 38782 31502 38834 31554
rect 42030 31502 42082 31554
rect 43822 31502 43874 31554
rect 44942 31502 44994 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 5742 31166 5794 31218
rect 15710 31166 15762 31218
rect 17278 31166 17330 31218
rect 18062 31166 18114 31218
rect 24222 31166 24274 31218
rect 24782 31166 24834 31218
rect 28926 31166 28978 31218
rect 30046 31166 30098 31218
rect 35870 31166 35922 31218
rect 36654 31166 36706 31218
rect 43822 31166 43874 31218
rect 44606 31166 44658 31218
rect 4958 31054 5010 31106
rect 8542 31054 8594 31106
rect 10782 31054 10834 31106
rect 14926 31054 14978 31106
rect 25230 31054 25282 31106
rect 29710 31054 29762 31106
rect 31950 31054 32002 31106
rect 38894 31054 38946 31106
rect 39678 31054 39730 31106
rect 2270 30942 2322 30994
rect 2718 30942 2770 30994
rect 6078 30942 6130 30994
rect 9998 30942 10050 30994
rect 11006 30942 11058 30994
rect 12126 30942 12178 30994
rect 12574 30942 12626 30994
rect 20302 30942 20354 30994
rect 20750 30942 20802 30994
rect 21086 30942 21138 30994
rect 21758 30942 21810 30994
rect 26014 30942 26066 30994
rect 26686 30942 26738 30994
rect 33070 30942 33122 30994
rect 33630 30942 33682 30994
rect 41134 30942 41186 30994
rect 41582 30942 41634 30994
rect 45054 30942 45106 30994
rect 7198 30830 7250 30882
rect 7534 30830 7586 30882
rect 10446 30830 10498 30882
rect 11454 30830 11506 30882
rect 11678 30830 11730 30882
rect 16158 30830 16210 30882
rect 16494 30830 16546 30882
rect 16830 30830 16882 30882
rect 25566 30830 25618 30882
rect 30942 30830 30994 30882
rect 36990 30830 37042 30882
rect 37438 30830 37490 30882
rect 37886 30830 37938 30882
rect 39902 30830 39954 30882
rect 44830 30830 44882 30882
rect 45614 30830 45666 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 4062 30270 4114 30322
rect 14926 30270 14978 30322
rect 26910 30270 26962 30322
rect 42142 30270 42194 30322
rect 45726 30270 45778 30322
rect 5630 30158 5682 30210
rect 6078 30158 6130 30210
rect 9214 30158 9266 30210
rect 9550 30158 9602 30210
rect 9886 30158 9938 30210
rect 13022 30158 13074 30210
rect 13694 30158 13746 30210
rect 14254 30158 14306 30210
rect 15598 30158 15650 30210
rect 18622 30158 18674 30210
rect 19070 30158 19122 30210
rect 20414 30158 20466 30210
rect 21534 30158 21586 30210
rect 25118 30158 25170 30210
rect 25678 30158 25730 30210
rect 29262 30158 29314 30210
rect 29710 30158 29762 30210
rect 32734 30158 32786 30210
rect 32846 30158 32898 30210
rect 35982 30158 36034 30210
rect 36542 30158 36594 30210
rect 37326 30158 37378 30210
rect 37774 30158 37826 30210
rect 40910 30158 40962 30210
rect 41694 30158 41746 30210
rect 44270 30158 44322 30210
rect 45054 30158 45106 30210
rect 1934 30046 1986 30098
rect 3054 30046 3106 30098
rect 13470 30046 13522 30098
rect 14590 30046 14642 30098
rect 15262 30046 15314 30098
rect 16382 30046 16434 30098
rect 20750 30046 20802 30098
rect 21758 30046 21810 30098
rect 27918 30046 27970 30098
rect 43150 30046 43202 30098
rect 43934 30046 43986 30098
rect 44830 30046 44882 30098
rect 45502 30046 45554 30098
rect 2046 29934 2098 29986
rect 8654 29934 8706 29986
rect 12462 29934 12514 29986
rect 21982 29934 22034 29986
rect 22766 29934 22818 29986
rect 32174 29934 32226 29986
rect 33518 29934 33570 29986
rect 40238 29934 40290 29986
rect 41246 29934 41298 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 7534 29598 7586 29650
rect 8206 29598 8258 29650
rect 8654 29598 8706 29650
rect 12350 29598 12402 29650
rect 13134 29598 13186 29650
rect 16382 29598 16434 29650
rect 16942 29598 16994 29650
rect 21982 29598 22034 29650
rect 26014 29598 26066 29650
rect 30942 29598 30994 29650
rect 31502 29598 31554 29650
rect 38782 29598 38834 29650
rect 40798 29598 40850 29650
rect 41582 29598 41634 29650
rect 44942 29598 44994 29650
rect 2270 29486 2322 29538
rect 17390 29486 17442 29538
rect 21198 29486 21250 29538
rect 22654 29486 22706 29538
rect 25230 29486 25282 29538
rect 27582 29486 27634 29538
rect 32062 29486 32114 29538
rect 33182 29486 33234 29538
rect 33518 29486 33570 29538
rect 37998 29486 38050 29538
rect 45838 29486 45890 29538
rect 4734 29374 4786 29426
rect 5070 29374 5122 29426
rect 9662 29374 9714 29426
rect 10110 29374 10162 29426
rect 13358 29374 13410 29426
rect 13918 29374 13970 29426
rect 17614 29374 17666 29426
rect 18398 29374 18450 29426
rect 18846 29374 18898 29426
rect 25454 29374 25506 29426
rect 25902 29374 25954 29426
rect 27918 29374 27970 29426
rect 28478 29374 28530 29426
rect 35310 29374 35362 29426
rect 35758 29374 35810 29426
rect 39118 29374 39170 29426
rect 43822 29374 43874 29426
rect 44382 29374 44434 29426
rect 3278 29262 3330 29314
rect 8766 29262 8818 29314
rect 23662 29262 23714 29314
rect 27022 29262 27074 29314
rect 27358 29262 27410 29314
rect 31726 29262 31778 29314
rect 40014 29262 40066 29314
rect 45054 29262 45106 29314
rect 45502 29262 45554 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 11790 28814 11842 28866
rect 18846 28814 18898 28866
rect 29038 28814 29090 28866
rect 36542 28814 36594 28866
rect 40574 28814 40626 28866
rect 44942 28814 44994 28866
rect 45390 28814 45442 28866
rect 1934 28702 1986 28754
rect 2158 28702 2210 28754
rect 4062 28702 4114 28754
rect 5630 28702 5682 28754
rect 7534 28702 7586 28754
rect 14030 28702 14082 28754
rect 14478 28702 14530 28754
rect 19070 28702 19122 28754
rect 21646 28702 21698 28754
rect 24222 28702 24274 28754
rect 28142 28702 28194 28754
rect 44942 28702 44994 28754
rect 45390 28702 45442 28754
rect 6302 28590 6354 28642
rect 6638 28590 6690 28642
rect 7422 28590 7474 28642
rect 8318 28590 8370 28642
rect 8766 28590 8818 28642
rect 12014 28590 12066 28642
rect 12238 28590 12290 28642
rect 12910 28590 12962 28642
rect 13582 28590 13634 28642
rect 14926 28590 14978 28642
rect 15150 28590 15202 28642
rect 15822 28590 15874 28642
rect 19294 28590 19346 28642
rect 20750 28590 20802 28642
rect 23774 28590 23826 28642
rect 24446 28590 24498 28642
rect 25006 28590 25058 28642
rect 26574 28590 26626 28642
rect 32174 28590 32226 28642
rect 32510 28590 32562 28642
rect 32846 28590 32898 28642
rect 33406 28590 33458 28642
rect 36990 28590 37042 28642
rect 37550 28590 37602 28642
rect 40798 28590 40850 28642
rect 41358 28590 41410 28642
rect 3054 28478 3106 28530
rect 5966 28478 6018 28530
rect 29822 28478 29874 28530
rect 11230 28366 11282 28418
rect 18062 28366 18114 28418
rect 35982 28366 36034 28418
rect 39902 28366 39954 28418
rect 43598 28366 43650 28418
rect 44382 28366 44434 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 3502 28030 3554 28082
rect 4286 28030 4338 28082
rect 8318 28030 8370 28082
rect 16382 28030 16434 28082
rect 16942 28030 16994 28082
rect 17502 28030 17554 28082
rect 20750 28030 20802 28082
rect 21534 28030 21586 28082
rect 29822 28030 29874 28082
rect 30606 28030 30658 28082
rect 31502 28030 31554 28082
rect 37326 28030 37378 28082
rect 44606 28030 44658 28082
rect 3278 27918 3330 27970
rect 36542 27918 36594 27970
rect 40910 27918 40962 27970
rect 41246 27918 41298 27970
rect 45838 27918 45890 27970
rect 6526 27806 6578 27858
rect 7198 27806 7250 27858
rect 10110 27806 10162 27858
rect 13358 27806 13410 27858
rect 13918 27806 13970 27858
rect 18286 27806 18338 27858
rect 23886 27806 23938 27858
rect 24446 27806 24498 27858
rect 25454 27806 25506 27858
rect 27134 27806 27186 27858
rect 27470 27806 27522 27858
rect 31838 27806 31890 27858
rect 33854 27806 33906 27858
rect 34302 27806 34354 27858
rect 37550 27806 37602 27858
rect 41470 27806 41522 27858
rect 42142 27806 42194 27858
rect 46062 27806 46114 27858
rect 2942 27694 2994 27746
rect 9886 27694 9938 27746
rect 11790 27694 11842 27746
rect 19070 27694 19122 27746
rect 25230 27694 25282 27746
rect 38670 27694 38722 27746
rect 45614 27694 45666 27746
rect 45166 27582 45218 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 16270 27246 16322 27298
rect 24894 27246 24946 27298
rect 25006 27246 25058 27298
rect 40574 27246 40626 27298
rect 44382 27246 44434 27298
rect 4062 27134 4114 27186
rect 5630 27134 5682 27186
rect 5966 27134 6018 27186
rect 12126 27134 12178 27186
rect 14926 27134 14978 27186
rect 20302 27134 20354 27186
rect 20526 27134 20578 27186
rect 34526 27134 34578 27186
rect 46174 27134 46226 27186
rect 6974 27022 7026 27074
rect 7982 27022 8034 27074
rect 8542 27022 8594 27074
rect 13470 27022 13522 27074
rect 19406 27022 19458 27074
rect 19742 27022 19794 27074
rect 21198 27022 21250 27074
rect 21870 27022 21922 27074
rect 28142 27022 28194 27074
rect 28702 27022 28754 27074
rect 30158 27022 30210 27074
rect 31838 27022 31890 27074
rect 36990 27022 37042 27074
rect 37438 27022 37490 27074
rect 40686 27022 40738 27074
rect 41358 27022 41410 27074
rect 44942 27022 44994 27074
rect 3054 26910 3106 26962
rect 6414 26910 6466 26962
rect 6750 26910 6802 26962
rect 11678 26910 11730 26962
rect 12574 26910 12626 26962
rect 12910 26910 12962 26962
rect 24110 26910 24162 26962
rect 35534 26910 35586 26962
rect 36430 26910 36482 26962
rect 39790 26910 39842 26962
rect 45726 26910 45778 26962
rect 11118 26798 11170 26850
rect 17054 26798 17106 26850
rect 25790 26798 25842 26850
rect 43822 26798 43874 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 1598 26462 1650 26514
rect 2382 26462 2434 26514
rect 8542 26462 8594 26514
rect 9102 26462 9154 26514
rect 9662 26462 9714 26514
rect 14926 26462 14978 26514
rect 17502 26462 17554 26514
rect 18062 26462 18114 26514
rect 22430 26462 22482 26514
rect 23214 26462 23266 26514
rect 28254 26462 28306 26514
rect 32958 26462 33010 26514
rect 36766 26462 36818 26514
rect 43822 26462 43874 26514
rect 11230 26350 11282 26402
rect 16494 26350 16546 26402
rect 18846 26350 18898 26402
rect 33742 26350 33794 26402
rect 37550 26350 37602 26402
rect 45390 26350 45442 26402
rect 4734 26238 4786 26290
rect 5182 26238 5234 26290
rect 5630 26238 5682 26290
rect 6078 26238 6130 26290
rect 11790 26238 11842 26290
rect 12350 26238 12402 26290
rect 19070 26238 19122 26290
rect 19630 26238 19682 26290
rect 20190 26238 20242 26290
rect 23886 26238 23938 26290
rect 25118 26238 25170 26290
rect 25678 26238 25730 26290
rect 29038 26238 29090 26290
rect 36094 26238 36146 26290
rect 36654 26238 36706 26290
rect 39902 26238 39954 26290
rect 40462 26238 40514 26290
rect 41022 26238 41074 26290
rect 41470 26238 41522 26290
rect 46174 26238 46226 26290
rect 9550 26126 9602 26178
rect 11566 26126 11618 26178
rect 15822 26126 15874 26178
rect 16046 26126 16098 26178
rect 16830 26126 16882 26178
rect 17950 26126 18002 26178
rect 23998 26126 24050 26178
rect 31390 26126 31442 26178
rect 44718 26126 44770 26178
rect 45054 26126 45106 26178
rect 45726 26126 45778 26178
rect 15486 26014 15538 26066
rect 28814 26014 28866 26066
rect 44494 26014 44546 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 13022 25678 13074 25730
rect 35310 25678 35362 25730
rect 4062 25566 4114 25618
rect 6974 25566 7026 25618
rect 16382 25566 16434 25618
rect 18958 25566 19010 25618
rect 23102 25566 23154 25618
rect 28254 25566 28306 25618
rect 37998 25566 38050 25618
rect 43822 25566 43874 25618
rect 44830 25566 44882 25618
rect 45502 25566 45554 25618
rect 8542 25454 8594 25506
rect 9550 25454 9602 25506
rect 9886 25454 9938 25506
rect 13694 25454 13746 25506
rect 14366 25454 14418 25506
rect 20302 25454 20354 25506
rect 24558 25454 24610 25506
rect 25006 25454 25058 25506
rect 31054 25454 31106 25506
rect 31614 25454 31666 25506
rect 32286 25454 32338 25506
rect 37774 25454 37826 25506
rect 38446 25454 38498 25506
rect 39006 25454 39058 25506
rect 43150 25454 43202 25506
rect 3054 25342 3106 25394
rect 13470 25342 13522 25394
rect 14142 25342 14194 25394
rect 15374 25342 15426 25394
rect 22094 25342 22146 25394
rect 28590 25342 28642 25394
rect 29598 25342 29650 25394
rect 30382 25342 30434 25394
rect 30830 25342 30882 25394
rect 35870 25342 35922 25394
rect 37326 25342 37378 25394
rect 42254 25342 42306 25394
rect 42926 25342 42978 25394
rect 43598 25342 43650 25394
rect 45166 25342 45218 25394
rect 8990 25230 9042 25282
rect 12462 25230 12514 25282
rect 20750 25230 20802 25282
rect 27246 25230 27298 25282
rect 28030 25230 28082 25282
rect 34750 25230 34802 25282
rect 35758 25230 35810 25282
rect 37214 25230 37266 25282
rect 41470 25230 41522 25282
rect 42030 25230 42082 25282
rect 42366 25230 42418 25282
rect 45614 25230 45666 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 3950 24894 4002 24946
rect 4734 24894 4786 24946
rect 12574 24894 12626 24946
rect 16158 24894 16210 24946
rect 20414 24894 20466 24946
rect 20974 24894 21026 24946
rect 23998 24894 24050 24946
rect 24782 24894 24834 24946
rect 29374 24894 29426 24946
rect 35982 24894 36034 24946
rect 44494 24894 44546 24946
rect 45054 24894 45106 24946
rect 2046 24782 2098 24834
rect 28590 24782 28642 24834
rect 41022 24782 41074 24834
rect 45502 24782 45554 24834
rect 1822 24670 1874 24722
rect 3502 24670 3554 24722
rect 6974 24670 7026 24722
rect 7646 24670 7698 24722
rect 9662 24670 9714 24722
rect 10110 24670 10162 24722
rect 13246 24670 13298 24722
rect 13918 24670 13970 24722
rect 17502 24670 17554 24722
rect 17838 24670 17890 24722
rect 21198 24670 21250 24722
rect 21646 24670 21698 24722
rect 25678 24670 25730 24722
rect 26350 24670 26402 24722
rect 32174 24670 32226 24722
rect 32958 24670 33010 24722
rect 33630 24670 33682 24722
rect 39454 24670 39506 24722
rect 41358 24670 41410 24722
rect 42030 24670 42082 24722
rect 2494 24558 2546 24610
rect 3614 24558 3666 24610
rect 31054 24558 31106 24610
rect 37102 24558 37154 24610
rect 38558 24558 38610 24610
rect 45726 24558 45778 24610
rect 13134 24446 13186 24498
rect 16942 24446 16994 24498
rect 36654 24446 36706 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 4062 23998 4114 24050
rect 7870 23998 7922 24050
rect 8430 23998 8482 24050
rect 14926 23998 14978 24050
rect 20414 23998 20466 24050
rect 22206 23998 22258 24050
rect 30158 23998 30210 24050
rect 32958 23998 33010 24050
rect 36206 23998 36258 24050
rect 36990 23998 37042 24050
rect 42478 23998 42530 24050
rect 42814 23998 42866 24050
rect 2046 23886 2098 23938
rect 9326 23886 9378 23938
rect 9662 23886 9714 23938
rect 19294 23886 19346 23938
rect 19966 23886 20018 23938
rect 23326 23886 23378 23938
rect 29262 23886 29314 23938
rect 35422 23886 35474 23938
rect 37886 23886 37938 23938
rect 38558 23886 38610 23938
rect 41582 23886 41634 23938
rect 45054 23886 45106 23938
rect 2270 23774 2322 23826
rect 3054 23774 3106 23826
rect 5630 23774 5682 23826
rect 5966 23774 6018 23826
rect 6638 23774 6690 23826
rect 14030 23774 14082 23826
rect 20750 23774 20802 23826
rect 21310 23774 21362 23826
rect 21646 23774 21698 23826
rect 22430 23774 22482 23826
rect 26798 23774 26850 23826
rect 31166 23774 31218 23826
rect 33966 23774 34018 23826
rect 43822 23774 43874 23826
rect 44830 23774 44882 23826
rect 8878 23662 8930 23714
rect 12238 23662 12290 23714
rect 12798 23662 12850 23714
rect 16270 23662 16322 23714
rect 17054 23662 17106 23714
rect 22542 23662 22594 23714
rect 37102 23662 37154 23714
rect 40798 23662 40850 23714
rect 45614 23662 45666 23714
rect 46062 23662 46114 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 5518 23326 5570 23378
rect 17502 23326 17554 23378
rect 22542 23326 22594 23378
rect 23326 23326 23378 23378
rect 24334 23326 24386 23378
rect 26574 23326 26626 23378
rect 30046 23326 30098 23378
rect 30606 23326 30658 23378
rect 37102 23326 37154 23378
rect 45166 23326 45218 23378
rect 46062 23326 46114 23378
rect 13918 23214 13970 23266
rect 19406 23214 19458 23266
rect 23886 23214 23938 23266
rect 26014 23214 26066 23266
rect 32062 23214 32114 23266
rect 33070 23214 33122 23266
rect 38110 23214 38162 23266
rect 39678 23214 39730 23266
rect 40910 23214 40962 23266
rect 2046 23102 2098 23154
rect 2606 23102 2658 23154
rect 2942 23102 2994 23154
rect 8878 23102 8930 23154
rect 12574 23102 12626 23154
rect 16158 23102 16210 23154
rect 16830 23102 16882 23154
rect 19630 23102 19682 23154
rect 20190 23102 20242 23154
rect 26686 23102 26738 23154
rect 26910 23102 26962 23154
rect 27582 23102 27634 23154
rect 33294 23102 33346 23154
rect 34414 23102 34466 23154
rect 34862 23102 34914 23154
rect 40014 23102 40066 23154
rect 41134 23102 41186 23154
rect 42030 23102 42082 23154
rect 42590 23102 42642 23154
rect 1934 22990 1986 23042
rect 6526 22990 6578 23042
rect 9662 22990 9714 23042
rect 10222 22990 10274 23042
rect 17390 22990 17442 23042
rect 18174 22990 18226 23042
rect 19070 22990 19122 23042
rect 23550 22990 23602 23042
rect 25790 22990 25842 23042
rect 31054 22990 31106 23042
rect 39118 22990 39170 23042
rect 6078 22878 6130 22930
rect 13134 22878 13186 22930
rect 37886 22878 37938 22930
rect 45726 22878 45778 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 2158 22430 2210 22482
rect 4062 22430 4114 22482
rect 16718 22430 16770 22482
rect 40574 22430 40626 22482
rect 2046 22318 2098 22370
rect 5518 22318 5570 22370
rect 6078 22318 6130 22370
rect 9550 22318 9602 22370
rect 9886 22318 9938 22370
rect 13806 22318 13858 22370
rect 17166 22318 17218 22370
rect 17838 22318 17890 22370
rect 21422 22318 21474 22370
rect 21870 22318 21922 22370
rect 25006 22318 25058 22370
rect 25678 22318 25730 22370
rect 32174 22318 32226 22370
rect 32734 22318 32786 22370
rect 33070 22318 33122 22370
rect 33518 22318 33570 22370
rect 37102 22318 37154 22370
rect 37550 22318 37602 22370
rect 40798 22318 40850 22370
rect 41358 22318 41410 22370
rect 45054 22318 45106 22370
rect 3054 22206 3106 22258
rect 13022 22206 13074 22258
rect 16382 22206 16434 22258
rect 8430 22094 8482 22146
rect 9214 22094 9266 22146
rect 12238 22094 12290 22146
rect 14478 22094 14530 22146
rect 20302 22094 20354 22146
rect 20862 22094 20914 22146
rect 24334 22094 24386 22146
rect 24894 22094 24946 22146
rect 28030 22094 28082 22146
rect 28702 22094 28754 22146
rect 29038 22094 29090 22146
rect 29822 22094 29874 22146
rect 35758 22094 35810 22146
rect 36542 22094 36594 22146
rect 39902 22094 39954 22146
rect 43822 22094 43874 22146
rect 44382 22094 44434 22146
rect 44830 22094 44882 22146
rect 46286 22094 46338 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2494 21758 2546 21810
rect 15038 21758 15090 21810
rect 21198 21758 21250 21810
rect 28478 21758 28530 21810
rect 39902 21758 39954 21810
rect 6078 21646 6130 21698
rect 11230 21646 11282 21698
rect 11566 21646 11618 21698
rect 11902 21646 11954 21698
rect 16382 21646 16434 21698
rect 16718 21646 16770 21698
rect 24334 21646 24386 21698
rect 32174 21646 32226 21698
rect 32510 21646 32562 21698
rect 35870 21646 35922 21698
rect 43710 21646 43762 21698
rect 4734 21534 4786 21586
rect 5406 21534 5458 21586
rect 5854 21534 5906 21586
rect 8542 21534 8594 21586
rect 9886 21534 9938 21586
rect 12126 21534 12178 21586
rect 12686 21534 12738 21586
rect 17950 21534 18002 21586
rect 23438 21534 23490 21586
rect 23886 21534 23938 21586
rect 24558 21534 24610 21586
rect 25342 21534 25394 21586
rect 26014 21534 26066 21586
rect 31278 21534 31330 21586
rect 33182 21534 33234 21586
rect 33630 21534 33682 21586
rect 36990 21534 37042 21586
rect 37326 21534 37378 21586
rect 40798 21534 40850 21586
rect 41470 21534 41522 21586
rect 45054 21534 45106 21586
rect 45614 21534 45666 21586
rect 6638 21422 6690 21474
rect 9662 21422 9714 21474
rect 10558 21422 10610 21474
rect 10894 21422 10946 21474
rect 18510 21422 18562 21474
rect 29486 21422 29538 21474
rect 45726 21422 45778 21474
rect 1710 21310 1762 21362
rect 15822 21310 15874 21362
rect 20414 21310 20466 21362
rect 29038 21310 29090 21362
rect 36654 21310 36706 21362
rect 40462 21310 40514 21362
rect 44494 21310 44546 21362
rect 44718 21310 44770 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 3838 20862 3890 20914
rect 21534 20862 21586 20914
rect 28590 20862 28642 20914
rect 33966 20862 34018 20914
rect 2046 20750 2098 20802
rect 5518 20750 5570 20802
rect 6190 20750 6242 20802
rect 12462 20750 12514 20802
rect 13022 20750 13074 20802
rect 13358 20750 13410 20802
rect 14030 20750 14082 20802
rect 20190 20750 20242 20802
rect 20862 20750 20914 20802
rect 23662 20750 23714 20802
rect 24446 20750 24498 20802
rect 25118 20750 25170 20802
rect 29262 20750 29314 20802
rect 29710 20750 29762 20802
rect 37102 20750 37154 20802
rect 37438 20750 37490 20802
rect 40686 20750 40738 20802
rect 41246 20750 41298 20802
rect 45054 20750 45106 20802
rect 2270 20638 2322 20690
rect 3054 20638 3106 20690
rect 9326 20638 9378 20690
rect 10110 20638 10162 20690
rect 34974 20638 35026 20690
rect 36094 20638 36146 20690
rect 46174 20638 46226 20690
rect 8654 20526 8706 20578
rect 9214 20526 9266 20578
rect 16382 20526 16434 20578
rect 17054 20526 17106 20578
rect 17166 20526 17218 20578
rect 17950 20526 18002 20578
rect 27582 20526 27634 20578
rect 28142 20526 28194 20578
rect 32174 20526 32226 20578
rect 32734 20526 32786 20578
rect 33630 20526 33682 20578
rect 35982 20526 36034 20578
rect 40014 20526 40066 20578
rect 40574 20526 40626 20578
rect 43822 20526 43874 20578
rect 44382 20526 44434 20578
rect 44830 20526 44882 20578
rect 45838 20526 45890 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 2494 20190 2546 20242
rect 40350 20190 40402 20242
rect 10222 20078 10274 20130
rect 16158 20078 16210 20130
rect 20414 20078 20466 20130
rect 23998 20078 24050 20130
rect 26910 20078 26962 20130
rect 32062 20078 32114 20130
rect 38894 20078 38946 20130
rect 39230 20078 39282 20130
rect 42926 20078 42978 20130
rect 45726 20078 45778 20130
rect 4958 19966 5010 20018
rect 5406 19966 5458 20018
rect 8542 19966 8594 20018
rect 12462 19966 12514 20018
rect 13022 19966 13074 20018
rect 13246 19966 13298 20018
rect 13918 19966 13970 20018
rect 17838 19966 17890 20018
rect 21086 19966 21138 20018
rect 21758 19966 21810 20018
rect 25454 19966 25506 20018
rect 29150 19966 29202 20018
rect 29598 19966 29650 20018
rect 33070 19966 33122 20018
rect 33294 19966 33346 20018
rect 33966 19966 34018 20018
rect 34638 19966 34690 20018
rect 39790 19966 39842 20018
rect 7870 19854 7922 19906
rect 18622 19854 18674 19906
rect 20862 19854 20914 19906
rect 25230 19854 25282 19906
rect 31054 19854 31106 19906
rect 33742 19854 33794 19906
rect 41918 19854 41970 19906
rect 43822 19854 43874 19906
rect 44158 19854 44210 19906
rect 44494 19854 44546 19906
rect 44942 19854 44994 19906
rect 1934 19742 1986 19794
rect 9438 19742 9490 19794
rect 16942 19742 16994 19794
rect 24782 19742 24834 19794
rect 26126 19742 26178 19794
rect 38334 19742 38386 19794
rect 43822 19742 43874 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 43486 19406 43538 19458
rect 3838 19294 3890 19346
rect 6862 19294 6914 19346
rect 7646 19294 7698 19346
rect 8094 19294 8146 19346
rect 19182 19294 19234 19346
rect 21422 19294 21474 19346
rect 21758 19294 21810 19346
rect 27806 19294 27858 19346
rect 35982 19294 36034 19346
rect 38558 19294 38610 19346
rect 41134 19294 41186 19346
rect 43822 19294 43874 19346
rect 44158 19294 44210 19346
rect 2046 19182 2098 19234
rect 8542 19182 8594 19234
rect 8990 19182 9042 19234
rect 13694 19182 13746 19234
rect 14366 19182 14418 19234
rect 14926 19182 14978 19234
rect 18286 19182 18338 19234
rect 18846 19182 18898 19234
rect 19406 19182 19458 19234
rect 25454 19182 25506 19234
rect 25790 19182 25842 19234
rect 29374 19182 29426 19234
rect 29822 19182 29874 19234
rect 33518 19182 33570 19234
rect 39454 19182 39506 19234
rect 42926 19182 42978 19234
rect 44942 19182 44994 19234
rect 2270 19070 2322 19122
rect 2830 19070 2882 19122
rect 6078 19070 6130 19122
rect 12238 19070 12290 19122
rect 12574 19070 12626 19122
rect 13470 19070 13522 19122
rect 14142 19070 14194 19122
rect 19742 19070 19794 19122
rect 23102 19070 23154 19122
rect 42142 19070 42194 19122
rect 46062 19070 46114 19122
rect 11454 18958 11506 19010
rect 12014 18958 12066 19010
rect 15150 18958 15202 19010
rect 15934 18958 15986 19010
rect 19854 18958 19906 19010
rect 22318 18958 22370 19010
rect 32286 18958 32338 19010
rect 32846 18958 32898 19010
rect 34078 18958 34130 19010
rect 36094 18958 36146 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 2158 18622 2210 18674
rect 5966 18622 6018 18674
rect 16382 18622 16434 18674
rect 32510 18622 32562 18674
rect 10222 18510 10274 18562
rect 18622 18510 18674 18562
rect 22094 18510 22146 18562
rect 23998 18510 24050 18562
rect 31054 18510 31106 18562
rect 35870 18510 35922 18562
rect 41582 18510 41634 18562
rect 4734 18398 4786 18450
rect 5294 18398 5346 18450
rect 8430 18398 8482 18450
rect 8878 18398 8930 18450
rect 12574 18398 12626 18450
rect 13022 18398 13074 18450
rect 13246 18398 13298 18450
rect 13918 18398 13970 18450
rect 17838 18398 17890 18450
rect 18174 18398 18226 18450
rect 19182 18398 19234 18450
rect 19742 18398 19794 18450
rect 23662 18398 23714 18450
rect 24334 18398 24386 18450
rect 25678 18398 25730 18450
rect 30270 18398 30322 18450
rect 31726 18398 31778 18450
rect 31950 18398 32002 18450
rect 33182 18398 33234 18450
rect 33630 18398 33682 18450
rect 36990 18398 37042 18450
rect 39454 18398 39506 18450
rect 40350 18398 40402 18450
rect 43822 18398 43874 18450
rect 44382 18398 44434 18450
rect 44942 18398 44994 18450
rect 18958 18286 19010 18338
rect 23326 18286 23378 18338
rect 28590 18286 28642 18338
rect 31390 18286 31442 18338
rect 37550 18286 37602 18338
rect 46062 18286 46114 18338
rect 1598 18174 1650 18226
rect 5406 18174 5458 18226
rect 9438 18174 9490 18226
rect 16942 18174 16994 18226
rect 22878 18174 22930 18226
rect 27582 18174 27634 18226
rect 36654 18174 36706 18226
rect 40798 18174 40850 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 3950 17726 4002 17778
rect 8318 17726 8370 17778
rect 15262 17726 15314 17778
rect 21646 17726 21698 17778
rect 21870 17726 21922 17778
rect 22542 17726 22594 17778
rect 28254 17726 28306 17778
rect 30270 17726 30322 17778
rect 34414 17726 34466 17778
rect 35758 17726 35810 17778
rect 36094 17726 36146 17778
rect 42254 17726 42306 17778
rect 2046 17614 2098 17666
rect 6638 17614 6690 17666
rect 9214 17614 9266 17666
rect 9662 17614 9714 17666
rect 13806 17614 13858 17666
rect 16942 17614 16994 17666
rect 17502 17614 17554 17666
rect 22766 17614 22818 17666
rect 23438 17614 23490 17666
rect 27582 17614 27634 17666
rect 30494 17614 30546 17666
rect 31166 17614 31218 17666
rect 34638 17614 34690 17666
rect 35310 17614 35362 17666
rect 37326 17614 37378 17666
rect 37662 17614 37714 17666
rect 45166 17614 45218 17666
rect 2270 17502 2322 17554
rect 3054 17502 3106 17554
rect 13582 17502 13634 17554
rect 16494 17502 16546 17554
rect 19854 17502 19906 17554
rect 22206 17502 22258 17554
rect 26686 17502 26738 17554
rect 27022 17502 27074 17554
rect 27806 17502 27858 17554
rect 35086 17502 35138 17554
rect 43262 17502 43314 17554
rect 44270 17502 44322 17554
rect 46062 17502 46114 17554
rect 5070 17390 5122 17442
rect 5854 17390 5906 17442
rect 12126 17390 12178 17442
rect 12686 17390 12738 17442
rect 14366 17390 14418 17442
rect 14814 17390 14866 17442
rect 20638 17390 20690 17442
rect 25902 17390 25954 17442
rect 26462 17390 26514 17442
rect 30158 17390 30210 17442
rect 33630 17390 33682 17442
rect 34190 17390 34242 17442
rect 40014 17390 40066 17442
rect 40798 17390 40850 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 2158 17054 2210 17106
rect 24110 17054 24162 17106
rect 36094 17054 36146 17106
rect 8318 16942 8370 16994
rect 10222 16942 10274 16994
rect 13470 16942 13522 16994
rect 14702 16942 14754 16994
rect 17726 16942 17778 16994
rect 18062 16942 18114 16994
rect 18846 16942 18898 16994
rect 25902 16942 25954 16994
rect 31838 16942 31890 16994
rect 36654 16942 36706 16994
rect 39678 16942 39730 16994
rect 43710 16942 43762 16994
rect 4622 16830 4674 16882
rect 5070 16830 5122 16882
rect 5406 16830 5458 16882
rect 6078 16830 6130 16882
rect 12462 16830 12514 16882
rect 13022 16830 13074 16882
rect 13694 16830 13746 16882
rect 21086 16830 21138 16882
rect 21758 16830 21810 16882
rect 28254 16830 28306 16882
rect 28814 16830 28866 16882
rect 28926 16830 28978 16882
rect 29486 16830 29538 16882
rect 33182 16830 33234 16882
rect 33630 16830 33682 16882
rect 36990 16830 37042 16882
rect 37326 16830 37378 16882
rect 41022 16830 41074 16882
rect 41470 16830 41522 16882
rect 44494 16830 44546 16882
rect 44942 16830 44994 16882
rect 46062 16830 46114 16882
rect 15822 16718 15874 16770
rect 19630 16718 19682 16770
rect 1598 16606 1650 16658
rect 9102 16606 9154 16658
rect 9438 16606 9490 16658
rect 24782 16606 24834 16658
rect 25118 16606 25170 16658
rect 32622 16606 32674 16658
rect 40462 16606 40514 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 1934 16158 1986 16210
rect 4062 16158 4114 16210
rect 6638 16158 6690 16210
rect 13582 16158 13634 16210
rect 18958 16158 19010 16210
rect 45502 16158 45554 16210
rect 8542 16046 8594 16098
rect 8878 16046 8930 16098
rect 14926 16046 14978 16098
rect 15262 16046 15314 16098
rect 24222 16046 24274 16098
rect 24894 16046 24946 16098
rect 25118 16046 25170 16098
rect 25678 16046 25730 16098
rect 29038 16046 29090 16098
rect 29710 16046 29762 16098
rect 33070 16046 33122 16098
rect 33518 16046 33570 16098
rect 39902 16046 39954 16098
rect 40574 16046 40626 16098
rect 40910 16046 40962 16098
rect 41358 16046 41410 16098
rect 45950 16046 46002 16098
rect 2270 15934 2322 15986
rect 2718 15934 2770 15986
rect 7758 15934 7810 15986
rect 18622 15934 18674 15986
rect 21982 15934 22034 15986
rect 27918 15934 27970 15986
rect 43598 15934 43650 15986
rect 5742 15822 5794 15874
rect 6302 15822 6354 15874
rect 11454 15822 11506 15874
rect 12014 15822 12066 15874
rect 12350 15822 12402 15874
rect 12910 15822 12962 15874
rect 14030 15822 14082 15874
rect 17838 15822 17890 15874
rect 18398 15822 18450 15874
rect 21198 15822 21250 15874
rect 28702 15822 28754 15874
rect 32174 15822 32226 15874
rect 32734 15822 32786 15874
rect 35758 15822 35810 15874
rect 36542 15822 36594 15874
rect 36878 15822 36930 15874
rect 37550 15822 37602 15874
rect 44382 15822 44434 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 1934 15486 1986 15538
rect 8206 15486 8258 15538
rect 10334 15486 10386 15538
rect 23214 15486 23266 15538
rect 28142 15486 28194 15538
rect 31614 15486 31666 15538
rect 41022 15486 41074 15538
rect 44830 15486 44882 15538
rect 45726 15486 45778 15538
rect 3390 15374 3442 15426
rect 9550 15374 9602 15426
rect 11902 15374 11954 15426
rect 15710 15374 15762 15426
rect 17502 15374 17554 15426
rect 24334 15374 24386 15426
rect 24670 15374 24722 15426
rect 27358 15374 27410 15426
rect 28030 15374 28082 15426
rect 33742 15374 33794 15426
rect 39454 15374 39506 15426
rect 45390 15374 45442 15426
rect 1934 15262 1986 15314
rect 5070 15262 5122 15314
rect 5630 15262 5682 15314
rect 20190 15262 20242 15314
rect 20862 15262 20914 15314
rect 28926 15262 28978 15314
rect 29262 15262 29314 15314
rect 35982 15262 36034 15314
rect 36654 15262 36706 15314
rect 41134 15262 41186 15314
rect 41694 15262 41746 15314
rect 42366 15262 42418 15314
rect 45614 15262 45666 15314
rect 2606 15150 2658 15202
rect 9886 15150 9938 15202
rect 10782 15150 10834 15202
rect 12798 15150 12850 15202
rect 14590 15150 14642 15202
rect 18734 15150 18786 15202
rect 26238 15150 26290 15202
rect 38334 15150 38386 15202
rect 8766 15038 8818 15090
rect 23886 15038 23938 15090
rect 32398 15038 32450 15090
rect 32958 15038 33010 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 3838 14590 3890 14642
rect 9662 14590 9714 14642
rect 9998 14590 10050 14642
rect 10446 14590 10498 14642
rect 16270 14590 16322 14642
rect 18622 14590 18674 14642
rect 34638 14590 34690 14642
rect 37998 14590 38050 14642
rect 40014 14590 40066 14642
rect 42814 14590 42866 14642
rect 8654 14478 8706 14530
rect 9214 14478 9266 14530
rect 23998 14478 24050 14530
rect 24446 14478 24498 14530
rect 29710 14478 29762 14530
rect 30382 14478 30434 14530
rect 39790 14478 39842 14530
rect 44830 14478 44882 14530
rect 1934 14366 1986 14418
rect 4958 14366 5010 14418
rect 11678 14366 11730 14418
rect 15038 14366 15090 14418
rect 19742 14366 19794 14418
rect 26686 14366 26738 14418
rect 35646 14366 35698 14418
rect 39006 14366 39058 14418
rect 43934 14366 43986 14418
rect 45950 14366 46002 14418
rect 2046 14254 2098 14306
rect 2718 14254 2770 14306
rect 3166 14254 3218 14306
rect 5518 14254 5570 14306
rect 6190 14254 6242 14306
rect 27470 14254 27522 14306
rect 32846 14254 32898 14306
rect 33406 14254 33458 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4846 13918 4898 13970
rect 8878 13918 8930 13970
rect 9662 13918 9714 13970
rect 6190 13806 6242 13858
rect 6974 13806 7026 13858
rect 13582 13806 13634 13858
rect 16382 13806 16434 13858
rect 20638 13806 20690 13858
rect 21310 13806 21362 13858
rect 24334 13806 24386 13858
rect 28030 13806 28082 13858
rect 29486 13806 29538 13858
rect 32174 13806 32226 13858
rect 32510 13806 32562 13858
rect 33070 13806 33122 13858
rect 33406 13806 33458 13858
rect 33742 13806 33794 13858
rect 34078 13806 34130 13858
rect 34526 13806 34578 13858
rect 34862 13806 34914 13858
rect 37438 13806 37490 13858
rect 42478 13806 42530 13858
rect 45390 13806 45442 13858
rect 1934 13694 1986 13746
rect 2606 13694 2658 13746
rect 24558 13694 24610 13746
rect 38446 13694 38498 13746
rect 42814 13694 42866 13746
rect 5854 13582 5906 13634
rect 7982 13582 8034 13634
rect 8430 13582 8482 13634
rect 12574 13582 12626 13634
rect 15374 13582 15426 13634
rect 19630 13582 19682 13634
rect 22430 13582 22482 13634
rect 27134 13582 27186 13634
rect 30606 13582 30658 13634
rect 36206 13582 36258 13634
rect 38558 13582 38610 13634
rect 43262 13582 43314 13634
rect 43822 13582 43874 13634
rect 44270 13582 44322 13634
rect 5630 13470 5682 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 3726 13022 3778 13074
rect 7870 13022 7922 13074
rect 10222 13022 10274 13074
rect 15486 13022 15538 13074
rect 19294 13022 19346 13074
rect 23886 13022 23938 13074
rect 26238 13022 26290 13074
rect 30270 13022 30322 13074
rect 33294 13022 33346 13074
rect 34862 13022 34914 13074
rect 35086 13022 35138 13074
rect 35870 13022 35922 13074
rect 36206 13022 36258 13074
rect 38110 13022 38162 13074
rect 41022 13022 41074 13074
rect 43598 13022 43650 13074
rect 45502 13022 45554 13074
rect 45054 12910 45106 12962
rect 46174 12910 46226 12962
rect 2382 12798 2434 12850
rect 6526 12798 6578 12850
rect 11230 12798 11282 12850
rect 16718 12798 16770 12850
rect 20526 12798 20578 12850
rect 22878 12798 22930 12850
rect 27246 12798 27298 12850
rect 31278 12798 31330 12850
rect 34302 12798 34354 12850
rect 39118 12798 39170 12850
rect 42030 12798 42082 12850
rect 5742 12686 5794 12738
rect 43038 12686 43090 12738
rect 44270 12686 44322 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 2270 12350 2322 12402
rect 5630 12350 5682 12402
rect 8094 12238 8146 12290
rect 13022 12238 13074 12290
rect 17950 12238 18002 12290
rect 23998 12238 24050 12290
rect 27582 12238 27634 12290
rect 30382 12238 30434 12290
rect 36430 12238 36482 12290
rect 37326 12238 37378 12290
rect 42926 12238 42978 12290
rect 45950 12238 46002 12290
rect 4622 12126 4674 12178
rect 5070 12126 5122 12178
rect 6974 12014 7026 12066
rect 12014 12014 12066 12066
rect 19070 12014 19122 12066
rect 22990 12014 23042 12066
rect 26574 12014 26626 12066
rect 29374 12014 29426 12066
rect 35086 12014 35138 12066
rect 38670 12014 38722 12066
rect 41918 12014 41970 12066
rect 44718 12014 44770 12066
rect 1598 11902 1650 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 45726 11566 45778 11618
rect 3502 11454 3554 11506
rect 6414 11454 6466 11506
rect 10446 11454 10498 11506
rect 22654 11454 22706 11506
rect 25230 11454 25282 11506
rect 30494 11454 30546 11506
rect 33406 11454 33458 11506
rect 35534 11454 35586 11506
rect 35870 11454 35922 11506
rect 36206 11454 36258 11506
rect 37998 11454 38050 11506
rect 42254 11454 42306 11506
rect 35310 11342 35362 11394
rect 2382 11230 2434 11282
rect 7758 11230 7810 11282
rect 9326 11230 9378 11282
rect 21534 11230 21586 11282
rect 26574 11230 26626 11282
rect 29374 11230 29426 11282
rect 34414 11230 34466 11282
rect 39230 11230 39282 11282
rect 43262 11230 43314 11282
rect 44942 11118 44994 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4510 10782 4562 10834
rect 44830 10782 44882 10834
rect 6750 10670 6802 10722
rect 11790 10670 11842 10722
rect 27918 10670 27970 10722
rect 35422 10670 35474 10722
rect 38670 10670 38722 10722
rect 43934 10670 43986 10722
rect 45726 10670 45778 10722
rect 1822 10558 1874 10610
rect 2270 10558 2322 10610
rect 46062 10558 46114 10610
rect 5966 10446 6018 10498
rect 10558 10446 10610 10498
rect 26574 10446 26626 10498
rect 34414 10446 34466 10498
rect 37438 10446 37490 10498
rect 42926 10446 42978 10498
rect 45502 10446 45554 10498
rect 5294 10334 5346 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 5854 9886 5906 9938
rect 10558 9886 10610 9938
rect 32734 9886 32786 9938
rect 38334 9886 38386 9938
rect 41134 9886 41186 9938
rect 45390 9886 45442 9938
rect 44046 9774 44098 9826
rect 9214 9662 9266 9714
rect 33966 9662 34018 9714
rect 39342 9662 39394 9714
rect 42142 9662 42194 9714
rect 43598 9662 43650 9714
rect 43262 9550 43314 9602
rect 44270 9550 44322 9602
rect 44942 9550 44994 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 43934 9214 43986 9266
rect 35646 9102 35698 9154
rect 41022 9102 41074 9154
rect 46062 9102 46114 9154
rect 34750 8878 34802 8930
rect 42142 8878 42194 8930
rect 44718 8878 44770 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 40238 8318 40290 8370
rect 45614 8318 45666 8370
rect 2830 8206 2882 8258
rect 2046 8094 2098 8146
rect 41246 8094 41298 8146
rect 44270 8094 44322 8146
rect 3390 7982 3442 8034
rect 43934 7982 43986 8034
rect 44942 7982 44994 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 44606 7646 44658 7698
rect 42366 7534 42418 7586
rect 46062 7534 46114 7586
rect 2942 7422 2994 7474
rect 44942 7422 44994 7474
rect 1934 7310 1986 7362
rect 3502 7310 3554 7362
rect 41470 7310 41522 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 41918 6750 41970 6802
rect 2942 6638 2994 6690
rect 45726 6638 45778 6690
rect 2046 6526 2098 6578
rect 42814 6526 42866 6578
rect 44942 6414 44994 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 22206 6078 22258 6130
rect 24446 6078 24498 6130
rect 33406 6078 33458 6130
rect 33854 6078 33906 6130
rect 20750 5966 20802 6018
rect 22990 5966 23042 6018
rect 23662 5966 23714 6018
rect 26462 5966 26514 6018
rect 45950 5966 46002 6018
rect 2942 5854 2994 5906
rect 20974 5854 21026 5906
rect 22430 5854 22482 5906
rect 23214 5854 23266 5906
rect 23998 5854 24050 5906
rect 26238 5854 26290 5906
rect 33070 5854 33122 5906
rect 1934 5742 1986 5794
rect 20414 5742 20466 5794
rect 28814 5742 28866 5794
rect 44942 5742 44994 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 24894 5182 24946 5234
rect 45614 5182 45666 5234
rect 46174 5182 46226 5234
rect 1710 5070 1762 5122
rect 2494 5070 2546 5122
rect 13694 5070 13746 5122
rect 14702 5070 14754 5122
rect 15598 5070 15650 5122
rect 16942 5070 16994 5122
rect 17502 5070 17554 5122
rect 18062 5070 18114 5122
rect 18622 5070 18674 5122
rect 19742 5070 19794 5122
rect 22766 5070 22818 5122
rect 23102 5070 23154 5122
rect 23886 5070 23938 5122
rect 24446 5070 24498 5122
rect 26126 5070 26178 5122
rect 28254 5070 28306 5122
rect 29374 5070 29426 5122
rect 30046 5070 30098 5122
rect 31278 5070 31330 5122
rect 31950 5070 32002 5122
rect 32622 5070 32674 5122
rect 33294 5070 33346 5122
rect 33966 5070 34018 5122
rect 37662 5070 37714 5122
rect 38334 5070 38386 5122
rect 39118 5070 39170 5122
rect 40126 5070 40178 5122
rect 41694 5070 41746 5122
rect 44046 5070 44098 5122
rect 44942 5070 44994 5122
rect 2046 4958 2098 5010
rect 12238 4958 12290 5010
rect 16606 4958 16658 5010
rect 17278 4958 17330 5010
rect 18398 4958 18450 5010
rect 20414 4958 20466 5010
rect 21758 4958 21810 5010
rect 22430 4958 22482 5010
rect 23438 4958 23490 5010
rect 24110 4958 24162 5010
rect 26686 4958 26738 5010
rect 27022 4958 27074 5010
rect 28478 4958 28530 5010
rect 30270 4958 30322 5010
rect 32846 4958 32898 5010
rect 38558 4958 38610 5010
rect 40350 4958 40402 5010
rect 44270 4958 44322 5010
rect 9438 4846 9490 4898
rect 12574 4846 12626 4898
rect 13470 4846 13522 4898
rect 15038 4846 15090 4898
rect 15934 4846 15986 4898
rect 19518 4846 19570 4898
rect 20078 4846 20130 4898
rect 20750 4846 20802 4898
rect 22094 4846 22146 4898
rect 26350 4846 26402 4898
rect 29598 4846 29650 4898
rect 30942 4846 30994 4898
rect 31502 4846 31554 4898
rect 32174 4846 32226 4898
rect 33518 4846 33570 4898
rect 34190 4846 34242 4898
rect 34750 4846 34802 4898
rect 35646 4846 35698 4898
rect 37886 4846 37938 4898
rect 39342 4846 39394 4898
rect 40910 4846 40962 4898
rect 43598 4846 43650 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 2046 4510 2098 4562
rect 8878 4510 8930 4562
rect 9998 4510 10050 4562
rect 14702 4510 14754 4562
rect 15038 4510 15090 4562
rect 17726 4510 17778 4562
rect 19406 4510 19458 4562
rect 21086 4510 21138 4562
rect 22654 4510 22706 4562
rect 26462 4510 26514 4562
rect 28030 4510 28082 4562
rect 30494 4510 30546 4562
rect 32174 4510 32226 4562
rect 33406 4510 33458 4562
rect 34078 4510 34130 4562
rect 35422 4510 35474 4562
rect 37214 4510 37266 4562
rect 39902 4510 39954 4562
rect 40910 4510 40962 4562
rect 44718 4510 44770 4562
rect 46174 4510 46226 4562
rect 10334 4398 10386 4450
rect 18398 4398 18450 4450
rect 19742 4398 19794 4450
rect 20078 4398 20130 4450
rect 23326 4398 23378 4450
rect 24446 4398 24498 4450
rect 29150 4398 29202 4450
rect 31166 4398 31218 4450
rect 34526 4398 34578 4450
rect 35870 4398 35922 4450
rect 41918 4398 41970 4450
rect 43598 4398 43650 4450
rect 44046 4398 44098 4450
rect 45166 4398 45218 4450
rect 45502 4398 45554 4450
rect 45838 4398 45890 4450
rect 1710 4286 1762 4338
rect 9662 4286 9714 4338
rect 13022 4286 13074 4338
rect 14366 4286 14418 4338
rect 17390 4286 17442 4338
rect 19070 4286 19122 4338
rect 22878 4286 22930 4338
rect 23550 4286 23602 4338
rect 24222 4286 24274 4338
rect 28254 4286 28306 4338
rect 30718 4286 30770 4338
rect 31390 4286 31442 4338
rect 31838 4286 31890 4338
rect 33182 4286 33234 4338
rect 33854 4286 33906 4338
rect 34862 4286 34914 4338
rect 36094 4286 36146 4338
rect 40126 4286 40178 4338
rect 41134 4286 41186 4338
rect 42142 4286 42194 4338
rect 44494 4286 44546 4338
rect 2494 4174 2546 4226
rect 11454 4174 11506 4226
rect 12014 4174 12066 4226
rect 13582 4174 13634 4226
rect 14142 4174 14194 4226
rect 15486 4174 15538 4226
rect 16830 4174 16882 4226
rect 21534 4174 21586 4226
rect 22318 4174 22370 4226
rect 26238 4174 26290 4226
rect 27694 4174 27746 4226
rect 30270 4174 30322 4226
rect 36654 4174 36706 4226
rect 37662 4174 37714 4226
rect 38558 4174 38610 4226
rect 39678 4174 39730 4226
rect 8094 4062 8146 4114
rect 11566 4062 11618 4114
rect 12014 4062 12066 4114
rect 12350 4062 12402 4114
rect 27246 4062 27298 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19070 3614 19122 3666
rect 19742 3614 19794 3666
rect 23214 3614 23266 3666
rect 25566 3614 25618 3666
rect 30494 3614 30546 3666
rect 32958 3614 33010 3666
rect 36990 3614 37042 3666
rect 40238 3614 40290 3666
rect 41806 3614 41858 3666
rect 42702 3614 42754 3666
rect 8766 3502 8818 3554
rect 10558 3502 10610 3554
rect 12238 3502 12290 3554
rect 13806 3502 13858 3554
rect 16270 3502 16322 3554
rect 18510 3502 18562 3554
rect 20190 3502 20242 3554
rect 21198 3502 21250 3554
rect 22430 3502 22482 3554
rect 25118 3502 25170 3554
rect 26462 3502 26514 3554
rect 26910 3502 26962 3554
rect 27694 3502 27746 3554
rect 28590 3502 28642 3554
rect 30046 3502 30098 3554
rect 32510 3502 32562 3554
rect 34302 3502 34354 3554
rect 34974 3502 35026 3554
rect 36542 3502 36594 3554
rect 39790 3502 39842 3554
rect 41358 3502 41410 3554
rect 46062 3502 46114 3554
rect 1710 3390 1762 3442
rect 2046 3390 2098 3442
rect 2942 3390 2994 3442
rect 6862 3390 6914 3442
rect 7198 3390 7250 3442
rect 7646 3390 7698 3442
rect 10894 3390 10946 3442
rect 11566 3390 11618 3442
rect 12574 3390 12626 3442
rect 21422 3390 21474 3442
rect 23662 3390 23714 3442
rect 23998 3390 24050 3442
rect 24670 3390 24722 3442
rect 26686 3390 26738 3442
rect 27358 3390 27410 3442
rect 29262 3390 29314 3442
rect 31614 3390 31666 3442
rect 33854 3390 33906 3442
rect 34078 3390 34130 3442
rect 34750 3390 34802 3442
rect 37886 3390 37938 3442
rect 38110 3390 38162 3442
rect 38446 3390 38498 3442
rect 38782 3390 38834 3442
rect 39118 3390 39170 3442
rect 45838 3390 45890 3442
rect 2382 3278 2434 3330
rect 7982 3278 8034 3330
rect 9774 3278 9826 3330
rect 11230 3278 11282 3330
rect 11902 3278 11954 3330
rect 13134 3278 13186 3330
rect 15598 3278 15650 3330
rect 17838 3278 17890 3330
rect 21758 3278 21810 3330
rect 35982 3278 36034 3330
rect 43038 3278 43090 3330
rect 43934 3278 43986 3330
rect 44382 3278 44434 3330
rect 44830 3278 44882 3330
rect 45278 3278 45330 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 43934 2382 43986 2434
rect 45278 2382 45330 2434
rect 8878 926 8930 978
rect 9774 926 9826 978
<< metal2 >>
rect 7392 47200 7504 48000
rect 8064 47200 8176 48000
rect 13440 47200 13552 48000
rect 14112 47200 14224 48000
rect 14784 47200 14896 48000
rect 16800 47200 16912 48000
rect 17472 47200 17584 48000
rect 18144 47200 18256 48000
rect 18816 47200 18928 48000
rect 19488 47200 19600 48000
rect 20160 47200 20272 48000
rect 20832 47200 20944 48000
rect 21504 47200 21616 48000
rect 22176 47200 22288 48000
rect 22848 47200 22960 48000
rect 23520 47200 23632 48000
rect 24192 47200 24304 48000
rect 24864 47200 24976 48000
rect 25536 47200 25648 48000
rect 26208 47200 26320 48000
rect 26880 47200 26992 48000
rect 27552 47200 27664 48000
rect 28224 47200 28336 48000
rect 28896 47200 29008 48000
rect 29568 47200 29680 48000
rect 30240 47200 30352 48000
rect 30912 47200 31024 48000
rect 31584 47200 31696 48000
rect 32256 47200 32368 48000
rect 34272 47200 34384 48000
rect 34944 47200 35056 48000
rect 35616 47200 35728 48000
rect 36288 47200 36400 48000
rect 36960 47200 37072 48000
rect 37632 47200 37744 48000
rect 38304 47200 38416 48000
rect 38976 47200 39088 48000
rect 39648 47200 39760 48000
rect 40320 47200 40432 48000
rect 40992 47200 41104 48000
rect 41664 47200 41776 48000
rect 42336 47200 42448 48000
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 7420 44436 7476 47200
rect 8092 44548 8148 47200
rect 8092 44482 8148 44492
rect 9772 44548 9828 44558
rect 7420 44434 7924 44436
rect 7420 44382 7422 44434
rect 7474 44382 7924 44434
rect 7420 44380 7924 44382
rect 7420 44370 7476 44380
rect 7868 44322 7924 44380
rect 9772 44434 9828 44492
rect 9772 44382 9774 44434
rect 9826 44382 9828 44434
rect 9772 44370 9828 44382
rect 13468 44436 13524 47200
rect 14140 44882 14196 47200
rect 14140 44830 14142 44882
rect 14194 44830 14196 44882
rect 14140 44818 14196 44830
rect 13468 44434 13748 44436
rect 13468 44382 13470 44434
rect 13522 44382 13748 44434
rect 13468 44380 13748 44382
rect 13468 44370 13524 44380
rect 7868 44270 7870 44322
rect 7922 44270 7924 44322
rect 7868 44258 7924 44270
rect 13692 44322 13748 44380
rect 13692 44270 13694 44322
rect 13746 44270 13748 44322
rect 13692 44258 13748 44270
rect 14812 44212 14868 47200
rect 14924 44882 14980 44894
rect 14924 44830 14926 44882
rect 14978 44830 14980 44882
rect 14924 44434 14980 44830
rect 16828 44882 16884 47200
rect 17500 45556 17556 47200
rect 17500 45500 17780 45556
rect 16828 44830 16830 44882
rect 16882 44830 16884 44882
rect 16828 44818 16884 44830
rect 17500 44882 17556 44894
rect 17500 44830 17502 44882
rect 17554 44830 17556 44882
rect 17500 44546 17556 44830
rect 17500 44494 17502 44546
rect 17554 44494 17556 44546
rect 17500 44482 17556 44494
rect 14924 44382 14926 44434
rect 14978 44382 14980 44434
rect 14924 44370 14980 44382
rect 14812 44146 14868 44156
rect 15932 44212 15988 44222
rect 15932 44118 15988 44156
rect 7644 44098 7700 44110
rect 7644 44046 7646 44098
rect 7698 44046 7700 44098
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 7532 42756 7588 42766
rect 7644 42756 7700 44046
rect 7532 42754 7700 42756
rect 7532 42702 7534 42754
rect 7586 42702 7700 42754
rect 7532 42700 7700 42702
rect 7756 44100 7812 44110
rect 7532 42690 7588 42700
rect 7756 42642 7812 44044
rect 9324 44100 9380 44110
rect 9324 44006 9380 44044
rect 14028 44098 14084 44110
rect 14028 44046 14030 44098
rect 14082 44046 14084 44098
rect 13916 42756 13972 42766
rect 14028 42756 14084 44046
rect 14364 44098 14420 44110
rect 14364 44046 14366 44098
rect 14418 44046 14420 44098
rect 14364 43708 14420 44046
rect 13916 42754 14084 42756
rect 13916 42702 13918 42754
rect 13970 42702 14084 42754
rect 13916 42700 14084 42702
rect 14140 43652 14420 43708
rect 17724 43762 17780 45500
rect 17724 43710 17726 43762
rect 17778 43710 17780 43762
rect 17724 43698 17780 43710
rect 13916 42690 13972 42700
rect 7756 42590 7758 42642
rect 7810 42590 7812 42642
rect 7756 42578 7812 42590
rect 14140 42642 14196 43652
rect 18172 43540 18228 47200
rect 18844 45556 18900 47200
rect 18844 45500 19348 45556
rect 18284 44100 18340 44110
rect 18284 44098 18900 44100
rect 18284 44046 18286 44098
rect 18338 44046 18900 44098
rect 18284 44044 18900 44046
rect 18284 44034 18340 44044
rect 18732 43650 18788 43662
rect 18732 43598 18734 43650
rect 18786 43598 18788 43650
rect 18396 43540 18452 43550
rect 18172 43538 18452 43540
rect 18172 43486 18398 43538
rect 18450 43486 18452 43538
rect 18172 43484 18452 43486
rect 18172 42866 18228 43484
rect 18396 43474 18452 43484
rect 18172 42814 18174 42866
rect 18226 42814 18228 42866
rect 18172 42802 18228 42814
rect 18732 42756 18788 43598
rect 18732 42690 18788 42700
rect 14140 42590 14142 42642
rect 14194 42590 14196 42642
rect 14140 42578 14196 42590
rect 18844 42642 18900 44044
rect 19068 43650 19124 43662
rect 19068 43598 19070 43650
rect 19122 43598 19124 43650
rect 19068 42754 19124 43598
rect 19292 43540 19348 45500
rect 19516 44434 19572 47200
rect 20188 44882 20244 47200
rect 20188 44830 20190 44882
rect 20242 44830 20244 44882
rect 20188 44818 20244 44830
rect 19516 44382 19518 44434
rect 19570 44382 19572 44434
rect 19516 44370 19572 44382
rect 20188 44322 20244 44334
rect 20188 44270 20190 44322
rect 20242 44270 20244 44322
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43708 20244 44270
rect 20860 43708 20916 47200
rect 20972 44882 21028 44894
rect 20972 44830 20974 44882
rect 21026 44830 21028 44882
rect 20972 44434 21028 44830
rect 20972 44382 20974 44434
rect 21026 44382 21028 44434
rect 20972 44370 21028 44382
rect 20188 43652 20356 43708
rect 19852 43540 19908 43550
rect 19292 43538 19908 43540
rect 19292 43486 19294 43538
rect 19346 43486 19854 43538
rect 19906 43486 19908 43538
rect 19292 43484 19908 43486
rect 19292 43474 19348 43484
rect 19852 43474 19908 43484
rect 19068 42702 19070 42754
rect 19122 42702 19124 42754
rect 19068 42690 19124 42702
rect 18844 42590 18846 42642
rect 18898 42590 18900 42642
rect 18844 42578 18900 42590
rect 20300 42644 20356 43652
rect 20412 43652 21140 43708
rect 20412 43650 20468 43652
rect 20412 43598 20414 43650
rect 20466 43598 20468 43650
rect 20412 43586 20468 43598
rect 21084 43650 21140 43652
rect 21084 43598 21086 43650
rect 21138 43598 21140 43650
rect 21084 43586 21140 43598
rect 21420 43650 21476 43662
rect 21420 43598 21422 43650
rect 21474 43598 21476 43650
rect 20860 43540 20916 43550
rect 20860 43446 20916 43484
rect 20636 42756 20692 42766
rect 20636 42662 20692 42700
rect 21420 42756 21476 43598
rect 21532 43540 21588 47200
rect 21980 44322 22036 44334
rect 21980 44270 21982 44322
rect 22034 44270 22036 44322
rect 21532 43474 21588 43484
rect 21756 43650 21812 43662
rect 21756 43598 21758 43650
rect 21810 43598 21812 43650
rect 21420 42690 21476 42700
rect 21644 42756 21700 42766
rect 21756 42756 21812 43598
rect 21644 42754 21812 42756
rect 21644 42702 21646 42754
rect 21698 42702 21812 42754
rect 21644 42700 21812 42702
rect 21644 42690 21700 42700
rect 20412 42644 20468 42654
rect 20300 42642 20468 42644
rect 20300 42590 20414 42642
rect 20466 42590 20468 42642
rect 20300 42588 20468 42590
rect 21980 42644 22036 44270
rect 22204 43708 22260 47200
rect 22876 43708 22932 47200
rect 23436 44436 23492 44446
rect 23548 44436 23604 47200
rect 23436 44434 23604 44436
rect 23436 44382 23438 44434
rect 23490 44382 23604 44434
rect 23436 44380 23604 44382
rect 23436 44370 23492 44380
rect 23884 44324 23940 44334
rect 23660 44322 23940 44324
rect 23660 44270 23886 44322
rect 23938 44270 23940 44322
rect 23660 44268 23940 44270
rect 22204 43652 22820 43708
rect 22876 43652 23044 43708
rect 22092 43540 22148 43550
rect 22428 43540 22484 43550
rect 22092 43446 22148 43484
rect 22316 43538 22484 43540
rect 22316 43486 22430 43538
rect 22482 43486 22484 43538
rect 22316 43484 22484 43486
rect 22204 42644 22260 42654
rect 21980 42642 22260 42644
rect 21980 42590 22206 42642
rect 22258 42590 22260 42642
rect 21980 42588 22260 42590
rect 20412 42578 20468 42588
rect 22204 42578 22260 42588
rect 1708 42532 1764 42542
rect 1708 42438 1764 42476
rect 21868 42530 21924 42542
rect 21868 42478 21870 42530
rect 21922 42478 21924 42530
rect 21868 42420 21924 42478
rect 22316 42420 22372 43484
rect 22428 43474 22484 43484
rect 22764 43428 22820 43652
rect 22988 43540 23044 43652
rect 22988 43474 23044 43484
rect 23324 43652 23380 43662
rect 22876 43428 22932 43438
rect 22764 43426 22932 43428
rect 22764 43374 22878 43426
rect 22930 43374 22932 43426
rect 22764 43372 22932 43374
rect 22876 43362 22932 43372
rect 22428 42756 22484 42766
rect 22428 42662 22484 42700
rect 23324 42754 23380 43596
rect 23324 42702 23326 42754
rect 23378 42702 23380 42754
rect 23324 42690 23380 42702
rect 23548 42644 23604 42654
rect 23660 42644 23716 44268
rect 23884 44258 23940 44268
rect 23996 43652 24052 43662
rect 23996 43558 24052 43596
rect 24220 43652 24276 47200
rect 24892 44548 24948 47200
rect 25564 45108 25620 47200
rect 26236 45556 26292 47200
rect 26236 45500 26852 45556
rect 24892 44482 24948 44492
rect 25340 45052 25620 45108
rect 25340 44436 25396 45052
rect 25564 44548 25620 44558
rect 25564 44454 25620 44492
rect 25340 44342 25396 44380
rect 26236 44324 26292 44334
rect 25900 44322 26292 44324
rect 25900 44270 26238 44322
rect 26290 44270 26292 44322
rect 25900 44268 26292 44270
rect 25228 43652 25284 43662
rect 24220 43586 24276 43596
rect 25004 43596 25228 43652
rect 23772 43540 23828 43550
rect 23772 43446 23828 43484
rect 24332 43540 24388 43550
rect 24332 43446 24388 43484
rect 25004 42866 25060 43596
rect 25228 43558 25284 43596
rect 25564 43650 25620 43662
rect 25564 43598 25566 43650
rect 25618 43598 25620 43650
rect 25004 42814 25006 42866
rect 25058 42814 25060 42866
rect 25004 42802 25060 42814
rect 25564 42754 25620 43598
rect 25564 42702 25566 42754
rect 25618 42702 25620 42754
rect 25564 42690 25620 42702
rect 23548 42642 23716 42644
rect 23548 42590 23550 42642
rect 23602 42590 23716 42642
rect 23548 42588 23716 42590
rect 25900 42642 25956 44268
rect 26236 44258 26292 44268
rect 26684 44098 26740 44110
rect 26684 44046 26686 44098
rect 26738 44046 26740 44098
rect 26460 43540 26516 43550
rect 25900 42590 25902 42642
rect 25954 42590 25956 42642
rect 23548 42578 23604 42588
rect 25900 42578 25956 42590
rect 26236 43538 26516 43540
rect 26236 43486 26462 43538
rect 26514 43486 26516 43538
rect 26236 43484 26516 43486
rect 26236 42642 26292 43484
rect 26460 43474 26516 43484
rect 26572 42756 26628 42766
rect 26684 42756 26740 44046
rect 26796 43708 26852 45500
rect 26908 44882 26964 47200
rect 27580 45332 27636 47200
rect 27580 45266 27636 45276
rect 26908 44830 26910 44882
rect 26962 44830 26964 44882
rect 26908 44818 26964 44830
rect 27580 44882 27636 44894
rect 27580 44830 27582 44882
rect 27634 44830 27636 44882
rect 26908 44436 26964 44446
rect 26908 44322 26964 44380
rect 26908 44270 26910 44322
rect 26962 44270 26964 44322
rect 26908 44258 26964 44270
rect 27580 44322 27636 44830
rect 27580 44270 27582 44322
rect 27634 44270 27636 44322
rect 27356 44098 27412 44110
rect 27356 44046 27358 44098
rect 27410 44046 27412 44098
rect 27356 43708 27412 44046
rect 27580 43764 27636 44270
rect 28252 44324 28308 47200
rect 28812 45332 28868 45342
rect 28812 44434 28868 45276
rect 28924 44882 28980 47200
rect 28924 44830 28926 44882
rect 28978 44830 28980 44882
rect 28924 44818 28980 44830
rect 29596 44548 29652 47200
rect 29596 44482 29652 44492
rect 30044 44882 30100 44894
rect 30044 44830 30046 44882
rect 30098 44830 30100 44882
rect 28812 44382 28814 44434
rect 28866 44382 28868 44434
rect 28812 44370 28868 44382
rect 28252 44268 28532 44324
rect 28364 44098 28420 44110
rect 28364 44046 28366 44098
rect 28418 44046 28420 44098
rect 27692 43764 27748 43774
rect 27580 43762 27748 43764
rect 27580 43710 27694 43762
rect 27746 43710 27748 43762
rect 27580 43708 27748 43710
rect 28364 43708 28420 44046
rect 26796 43652 26964 43708
rect 26908 43426 26964 43652
rect 26908 43374 26910 43426
rect 26962 43374 26964 43426
rect 26908 43362 26964 43374
rect 27020 43652 27412 43708
rect 27692 43698 27748 43708
rect 28140 43652 28420 43708
rect 28476 43708 28532 44268
rect 29932 44098 29988 44110
rect 29932 44046 29934 44098
rect 29986 44046 29988 44098
rect 28476 43652 28980 43708
rect 26572 42754 26740 42756
rect 26572 42702 26574 42754
rect 26626 42702 26740 42754
rect 26572 42700 26740 42702
rect 26572 42690 26628 42700
rect 26236 42590 26238 42642
rect 26290 42590 26292 42642
rect 26236 42578 26292 42590
rect 19836 42364 20100 42374
rect 21868 42364 22372 42420
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 26908 41972 26964 41982
rect 27020 41972 27076 43652
rect 27804 43540 27860 43550
rect 27132 42196 27188 42206
rect 27132 42102 27188 42140
rect 27804 42194 27860 43484
rect 27804 42142 27806 42194
rect 27858 42142 27860 42194
rect 27804 42130 27860 42142
rect 28140 42194 28196 43652
rect 28476 43540 28532 43550
rect 28476 43446 28532 43484
rect 28924 43426 28980 43652
rect 29820 43540 29876 43550
rect 29820 43446 29876 43484
rect 28924 43374 28926 43426
rect 28978 43374 28980 43426
rect 28924 43362 28980 43374
rect 28140 42142 28142 42194
rect 28194 42142 28196 42194
rect 28140 42130 28196 42142
rect 28476 42980 28532 42990
rect 26908 41970 27076 41972
rect 26908 41918 26910 41970
rect 26962 41918 27076 41970
rect 26908 41916 27076 41918
rect 27580 42084 27636 42094
rect 27580 41970 27636 42028
rect 28476 42082 28532 42924
rect 29932 42196 29988 44046
rect 30044 43762 30100 44830
rect 30268 43764 30324 47200
rect 30380 44548 30436 44558
rect 30380 44434 30436 44492
rect 30940 44548 30996 47200
rect 30940 44482 30996 44492
rect 30380 44382 30382 44434
rect 30434 44382 30436 44434
rect 30380 44370 30436 44382
rect 30044 43710 30046 43762
rect 30098 43710 30100 43762
rect 30044 43698 30100 43710
rect 30156 43708 30324 43764
rect 30156 43540 30212 43708
rect 30492 43652 30548 43662
rect 30156 43474 30212 43484
rect 30268 43650 30548 43652
rect 30268 43598 30494 43650
rect 30546 43598 30548 43650
rect 30268 43596 30548 43598
rect 29932 42130 29988 42140
rect 28476 42030 28478 42082
rect 28530 42030 28532 42082
rect 28476 42018 28532 42030
rect 27580 41918 27582 41970
rect 27634 41918 27636 41970
rect 26908 41906 26964 41916
rect 27580 41906 27636 41918
rect 30268 41970 30324 43596
rect 30492 43586 30548 43596
rect 31612 43652 31668 47200
rect 32284 45218 32340 47200
rect 32284 45166 32286 45218
rect 32338 45166 32340 45218
rect 32284 45154 32340 45166
rect 33404 45218 33460 45230
rect 33404 45166 33406 45218
rect 33458 45166 33460 45218
rect 32620 44548 32676 44558
rect 32620 44434 32676 44492
rect 32620 44382 32622 44434
rect 32674 44382 32676 44434
rect 32620 44370 32676 44382
rect 33404 44436 33460 45166
rect 34300 45108 34356 47200
rect 34300 45052 34580 45108
rect 33404 44434 34020 44436
rect 33404 44382 33406 44434
rect 33458 44382 34020 44434
rect 33404 44380 34020 44382
rect 33404 44370 33460 44380
rect 33964 44322 34020 44380
rect 34524 44324 34580 45052
rect 33964 44270 33966 44322
rect 34018 44270 34020 44322
rect 33964 44258 34020 44270
rect 34300 44322 34580 44324
rect 34300 44270 34526 44322
rect 34578 44270 34580 44322
rect 34300 44268 34580 44270
rect 32172 44098 32228 44110
rect 32172 44046 32174 44098
rect 32226 44046 32228 44098
rect 31612 43558 31668 43596
rect 31836 43650 31892 43662
rect 31836 43598 31838 43650
rect 31890 43598 31892 43650
rect 30716 43540 30772 43550
rect 30716 43446 30772 43484
rect 30492 42196 30548 42206
rect 30492 42102 30548 42140
rect 31836 42084 31892 43598
rect 32060 43652 32116 43662
rect 32060 43538 32116 43596
rect 32060 43486 32062 43538
rect 32114 43486 32116 43538
rect 32060 43474 32116 43486
rect 32172 42196 32228 44046
rect 33740 44098 33796 44110
rect 33740 44046 33742 44098
rect 33794 44046 33796 44098
rect 33740 42980 33796 44046
rect 34300 43762 34356 44268
rect 34524 44258 34580 44268
rect 34300 43710 34302 43762
rect 34354 43710 34356 43762
rect 34300 43698 34356 43710
rect 34860 44098 34916 44110
rect 34860 44046 34862 44098
rect 34914 44046 34916 44098
rect 33740 42914 33796 42924
rect 34860 42756 34916 44046
rect 34972 43652 35028 47200
rect 35644 45668 35700 47200
rect 35644 45612 36036 45668
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35980 44210 36036 45612
rect 36316 44548 36372 47200
rect 36988 44882 37044 47200
rect 37660 45556 37716 47200
rect 38332 45668 38388 47200
rect 38332 45612 38612 45668
rect 37660 45500 38388 45556
rect 36988 44830 36990 44882
rect 37042 44830 37044 44882
rect 36988 44818 37044 44830
rect 38108 44882 38164 44894
rect 38108 44830 38110 44882
rect 38162 44830 38164 44882
rect 36316 44482 36372 44492
rect 37100 44548 37156 44558
rect 36764 44436 36820 44446
rect 36764 44342 36820 44380
rect 37100 44434 37156 44492
rect 37100 44382 37102 44434
rect 37154 44382 37156 44434
rect 37100 44370 37156 44382
rect 37660 44324 37716 44334
rect 38108 44324 38164 44830
rect 35980 44158 35982 44210
rect 36034 44158 36036 44210
rect 35980 44146 36036 44158
rect 37436 44322 37716 44324
rect 37436 44270 37662 44322
rect 37714 44270 37716 44322
rect 37436 44268 37716 44270
rect 35196 43652 35252 43662
rect 34972 43650 35252 43652
rect 34972 43598 34974 43650
rect 35026 43598 35198 43650
rect 35250 43598 35252 43650
rect 34972 43596 35252 43598
rect 34972 43586 35028 43596
rect 35196 43586 35252 43596
rect 35532 43650 35588 43662
rect 35532 43598 35534 43650
rect 35586 43598 35588 43650
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34860 42690 34916 42700
rect 32172 42130 32228 42140
rect 31836 42018 31892 42028
rect 30268 41918 30270 41970
rect 30322 41918 30324 41970
rect 30268 41906 30324 41918
rect 35532 41972 35588 43598
rect 37436 42194 37492 44268
rect 37660 44258 37716 44268
rect 37884 44322 38164 44324
rect 37884 44270 38110 44322
rect 38162 44270 38164 44322
rect 37884 44268 38164 44270
rect 37884 43762 37940 44268
rect 38108 44258 38164 44268
rect 37884 43710 37886 43762
rect 37938 43710 37940 43762
rect 37884 43698 37940 43710
rect 38332 43650 38388 45500
rect 38556 45220 38612 45612
rect 38556 45164 38836 45220
rect 38780 44436 38836 45164
rect 39004 44548 39060 47200
rect 39676 45556 39732 47200
rect 39676 45500 39956 45556
rect 39004 44482 39060 44492
rect 38780 44322 38836 44380
rect 38780 44270 38782 44322
rect 38834 44270 38836 44322
rect 38780 44258 38836 44270
rect 38892 44324 38948 44334
rect 38332 43598 38334 43650
rect 38386 43598 38388 43650
rect 38332 43586 38388 43598
rect 38444 44098 38500 44110
rect 38444 44046 38446 44098
rect 38498 44046 38500 44098
rect 38220 42756 38276 42766
rect 38220 42662 38276 42700
rect 37436 42142 37438 42194
rect 37490 42142 37492 42194
rect 37436 42130 37492 42142
rect 38444 42082 38500 44046
rect 38892 43708 38948 44268
rect 38780 43652 38948 43708
rect 39116 44098 39172 44110
rect 39788 44100 39844 44110
rect 39116 44046 39118 44098
rect 39170 44046 39172 44098
rect 38556 43540 38612 43550
rect 38556 42642 38612 43484
rect 38556 42590 38558 42642
rect 38610 42590 38612 42642
rect 38556 42578 38612 42590
rect 38780 42194 38836 43652
rect 39004 43540 39060 43550
rect 39004 43446 39060 43484
rect 39004 42756 39060 42766
rect 39116 42756 39172 44046
rect 39004 42754 39172 42756
rect 39004 42702 39006 42754
rect 39058 42702 39172 42754
rect 39004 42700 39172 42702
rect 39228 44098 39844 44100
rect 39228 44046 39790 44098
rect 39842 44046 39844 44098
rect 39228 44044 39844 44046
rect 39004 42690 39060 42700
rect 39228 42642 39284 44044
rect 39788 44034 39844 44044
rect 39676 43652 39732 43662
rect 39900 43652 39956 45500
rect 40348 44882 40404 47200
rect 41020 45556 41076 47200
rect 41692 45556 41748 47200
rect 41020 45500 41524 45556
rect 41692 45500 41860 45556
rect 40348 44830 40350 44882
rect 40402 44830 40404 44882
rect 40348 44818 40404 44830
rect 40236 44548 40292 44558
rect 40236 44436 40292 44492
rect 40348 44436 40404 44446
rect 40236 44434 40404 44436
rect 40236 44382 40350 44434
rect 40402 44382 40404 44434
rect 40236 44380 40404 44382
rect 40348 44370 40404 44380
rect 41356 44098 41412 44110
rect 41356 44046 41358 44098
rect 41410 44046 41412 44098
rect 41356 43708 41412 44046
rect 39676 43650 39956 43652
rect 39676 43598 39678 43650
rect 39730 43598 39902 43650
rect 39954 43598 39956 43650
rect 39676 43596 39956 43598
rect 39676 43586 39732 43596
rect 39900 43586 39956 43596
rect 40236 43650 40292 43662
rect 40236 43598 40238 43650
rect 40290 43598 40292 43650
rect 39676 42756 39732 42766
rect 39676 42662 39732 42700
rect 40236 42754 40292 43598
rect 40236 42702 40238 42754
rect 40290 42702 40292 42754
rect 40236 42690 40292 42702
rect 40572 43652 41412 43708
rect 41468 43708 41524 45500
rect 41468 43652 41748 43708
rect 39228 42590 39230 42642
rect 39282 42590 39284 42642
rect 39228 42578 39284 42590
rect 39900 42644 39956 42654
rect 39900 42550 39956 42588
rect 40572 42642 40628 43652
rect 40572 42590 40574 42642
rect 40626 42590 40628 42642
rect 40572 42578 40628 42590
rect 41244 43538 41300 43550
rect 41244 43486 41246 43538
rect 41298 43486 41300 43538
rect 41244 42644 41300 43486
rect 41692 43426 41748 43652
rect 41804 43652 41860 45500
rect 41916 44882 41972 44894
rect 41916 44830 41918 44882
rect 41970 44830 41972 44882
rect 41916 44434 41972 44830
rect 42364 44548 42420 47200
rect 42364 44482 42420 44492
rect 44044 44548 44100 44558
rect 41916 44382 41918 44434
rect 41970 44382 41972 44434
rect 41916 44370 41972 44382
rect 44044 44434 44100 44492
rect 44044 44382 44046 44434
rect 44098 44382 44100 44434
rect 44044 44370 44100 44382
rect 45724 44436 45780 44446
rect 43708 44324 43764 44334
rect 43708 44230 43764 44268
rect 44044 44100 44100 44110
rect 41804 43586 41860 43596
rect 42588 43652 42644 43662
rect 42588 43558 42644 43596
rect 42812 43650 42868 43662
rect 42812 43598 42814 43650
rect 42866 43598 42868 43650
rect 41692 43374 41694 43426
rect 41746 43374 41748 43426
rect 41692 43362 41748 43374
rect 42812 42756 42868 43598
rect 43036 43652 43092 43662
rect 43036 43538 43092 43596
rect 43036 43486 43038 43538
rect 43090 43486 43092 43538
rect 43036 43474 43092 43486
rect 42812 42690 42868 42700
rect 44044 42754 44100 44044
rect 45612 44098 45668 44110
rect 45612 44046 45614 44098
rect 45666 44046 45668 44098
rect 45612 43764 45668 44046
rect 45612 43698 45668 43708
rect 44044 42702 44046 42754
rect 44098 42702 44100 42754
rect 44044 42690 44100 42702
rect 45052 43538 45108 43550
rect 45052 43486 45054 43538
rect 45106 43486 45108 43538
rect 41244 42578 41300 42588
rect 44268 42532 44324 42542
rect 44940 42532 44996 42542
rect 44268 42530 44996 42532
rect 44268 42478 44270 42530
rect 44322 42478 44942 42530
rect 44994 42478 44996 42530
rect 44268 42476 44996 42478
rect 44268 42466 44324 42476
rect 44940 42466 44996 42476
rect 45052 42196 45108 43486
rect 45724 42978 45780 44380
rect 46172 44210 46228 44222
rect 46172 44158 46174 44210
rect 46226 44158 46228 44210
rect 45836 44100 45892 44110
rect 45836 44006 45892 44044
rect 46172 43764 46228 44158
rect 46172 43698 46228 43708
rect 46060 43426 46116 43438
rect 46060 43374 46062 43426
rect 46114 43374 46116 43426
rect 46060 43092 46116 43374
rect 46060 43026 46116 43036
rect 45724 42926 45726 42978
rect 45778 42926 45780 42978
rect 45724 42914 45780 42926
rect 38780 42142 38782 42194
rect 38834 42142 38836 42194
rect 38780 42130 38836 42142
rect 44828 42140 45108 42196
rect 46060 42420 46116 42430
rect 38444 42030 38446 42082
rect 38498 42030 38500 42082
rect 38444 42018 38500 42030
rect 44156 42084 44212 42094
rect 44156 42082 44660 42084
rect 44156 42030 44158 42082
rect 44210 42030 44660 42082
rect 44156 42028 44660 42030
rect 44156 42018 44212 42028
rect 35532 41906 35588 41916
rect 37100 41972 37156 41982
rect 37100 41878 37156 41916
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 44156 40290 44212 40302
rect 44156 40238 44158 40290
rect 44210 40238 44212 40290
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 38556 39732 38612 39742
rect 38444 39676 38556 39732
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 36316 38948 36372 38958
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 17836 38162 17892 38174
rect 17836 38110 17838 38162
rect 17890 38110 17892 38162
rect 17052 37940 17108 37950
rect 12796 37380 12852 37390
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 6188 35812 6244 35822
rect 5964 35810 6244 35812
rect 5964 35758 6190 35810
rect 6242 35758 6244 35810
rect 5964 35756 6244 35758
rect 5180 35588 5236 35598
rect 4844 35586 5236 35588
rect 4844 35534 5182 35586
rect 5234 35534 5236 35586
rect 4844 35532 5236 35534
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1708 34804 1764 34814
rect 1708 34354 1764 34748
rect 2268 34356 2324 34366
rect 1708 34302 1710 34354
rect 1762 34302 1764 34354
rect 1708 34290 1764 34302
rect 2156 34354 2324 34356
rect 2156 34302 2270 34354
rect 2322 34302 2324 34354
rect 2156 34300 2324 34302
rect 2044 31556 2100 31566
rect 1596 30436 1652 30446
rect 1596 26514 1652 30380
rect 1932 30098 1988 30110
rect 1932 30046 1934 30098
rect 1986 30046 1988 30098
rect 1932 28754 1988 30046
rect 2044 29986 2100 31500
rect 2044 29934 2046 29986
rect 2098 29934 2100 29986
rect 2044 29922 2100 29934
rect 1932 28702 1934 28754
rect 1986 28702 1988 28754
rect 1932 27972 1988 28702
rect 2156 28754 2212 34300
rect 2268 34290 2324 34300
rect 4844 34130 4900 35532
rect 5180 35522 5236 35532
rect 4844 34078 4846 34130
rect 4898 34078 4900 34130
rect 4844 34066 4900 34078
rect 5404 34130 5460 34142
rect 5404 34078 5406 34130
rect 5458 34078 5460 34130
rect 5404 34020 5460 34078
rect 5852 34020 5908 34030
rect 5404 33964 5852 34020
rect 5852 33926 5908 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 3612 33458 3668 33470
rect 3612 33406 3614 33458
rect 3666 33406 3668 33458
rect 2380 32562 2436 32574
rect 2380 32510 2382 32562
rect 2434 32510 2436 32562
rect 2380 31948 2436 32510
rect 2940 32564 2996 32574
rect 2940 32470 2996 32508
rect 3612 32564 3668 33406
rect 3612 32498 3668 32508
rect 4956 33234 5012 33246
rect 5964 33236 6020 35756
rect 6188 35746 6244 35756
rect 8652 35026 8708 35038
rect 9996 35028 10052 35038
rect 8652 34974 8654 35026
rect 8706 34974 8708 35026
rect 7308 34804 7364 34814
rect 7308 34710 7364 34748
rect 4956 33182 4958 33234
rect 5010 33182 5012 33234
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 2268 31892 2436 31948
rect 2716 31892 2772 31902
rect 2268 30994 2324 31892
rect 2268 30942 2270 30994
rect 2322 30942 2324 30994
rect 2268 30324 2324 30942
rect 2380 31666 2436 31678
rect 2380 31614 2382 31666
rect 2434 31614 2436 31666
rect 2380 30436 2436 31614
rect 2716 30994 2772 31836
rect 3500 31892 3556 31902
rect 4956 31892 5012 33182
rect 5740 33180 6020 33236
rect 6076 34244 6132 34254
rect 5516 32788 5572 32798
rect 5516 32786 5684 32788
rect 5516 32734 5518 32786
rect 5570 32734 5684 32786
rect 5516 32732 5684 32734
rect 5516 32722 5572 32732
rect 5516 31892 5572 31902
rect 4956 31890 5572 31892
rect 4956 31838 5518 31890
rect 5570 31838 5572 31890
rect 4956 31836 5572 31838
rect 3500 31798 3556 31836
rect 5516 31826 5572 31836
rect 2716 30942 2718 30994
rect 2770 30942 2772 30994
rect 2716 30930 2772 30942
rect 4956 31106 5012 31118
rect 5628 31108 5684 32732
rect 5740 31218 5796 33180
rect 6076 32786 6132 34188
rect 8540 34244 8596 34254
rect 8540 34150 8596 34188
rect 6076 32734 6078 32786
rect 6130 32734 6132 32786
rect 6076 32722 6132 32734
rect 6188 34020 6244 34030
rect 6636 34020 6692 34030
rect 6188 33122 6244 33964
rect 6188 33070 6190 33122
rect 6242 33070 6244 33122
rect 6076 31556 6132 31566
rect 6076 31462 6132 31500
rect 5740 31166 5742 31218
rect 5794 31166 5796 31218
rect 5740 31154 5796 31166
rect 4956 31054 4958 31106
rect 5010 31054 5012 31106
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 2380 30370 2436 30380
rect 2268 30258 2324 30268
rect 4060 30322 4116 30334
rect 4060 30270 4062 30322
rect 4114 30270 4116 30322
rect 3052 30098 3108 30110
rect 3052 30046 3054 30098
rect 3106 30046 3108 30098
rect 3052 29652 3108 30046
rect 4060 30100 4116 30270
rect 4060 30034 4116 30044
rect 4732 30212 4788 30222
rect 3052 29586 3108 29596
rect 2156 28702 2158 28754
rect 2210 28702 2212 28754
rect 2156 28690 2212 28702
rect 2268 29538 2324 29550
rect 2268 29486 2270 29538
rect 2322 29486 2324 29538
rect 2268 28084 2324 29486
rect 3500 29428 3556 29438
rect 3276 29316 3332 29326
rect 3500 29316 3556 29372
rect 4732 29426 4788 30156
rect 4732 29374 4734 29426
rect 4786 29374 4788 29426
rect 4732 29362 4788 29374
rect 3276 29314 3556 29316
rect 3276 29262 3278 29314
rect 3330 29262 3556 29314
rect 3276 29260 3556 29262
rect 3276 29250 3332 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4060 28754 4116 28766
rect 4060 28702 4062 28754
rect 4114 28702 4116 28754
rect 3052 28532 3108 28542
rect 3052 28530 3220 28532
rect 3052 28478 3054 28530
rect 3106 28478 3220 28530
rect 3052 28476 3220 28478
rect 3052 28466 3108 28476
rect 2268 28018 2324 28028
rect 1932 27906 1988 27916
rect 2940 27748 2996 27758
rect 1596 26462 1598 26514
rect 1650 26462 1652 26514
rect 1596 26450 1652 26462
rect 2380 27746 2996 27748
rect 2380 27694 2942 27746
rect 2994 27694 2996 27746
rect 2380 27692 2996 27694
rect 2380 26514 2436 27692
rect 2940 27682 2996 27692
rect 3052 26964 3108 26974
rect 3052 26870 3108 26908
rect 2380 26462 2382 26514
rect 2434 26462 2436 26514
rect 2380 26450 2436 26462
rect 3164 26516 3220 28476
rect 3500 28084 3556 28094
rect 3500 27990 3556 28028
rect 3276 27972 3332 27982
rect 3276 27878 3332 27916
rect 4060 27860 4116 28702
rect 4956 28756 5012 31054
rect 5516 31052 5684 31108
rect 5068 29428 5124 29438
rect 5068 29334 5124 29372
rect 4956 28690 5012 28700
rect 4284 28644 4340 28654
rect 4284 28082 4340 28588
rect 4284 28030 4286 28082
rect 4338 28030 4340 28082
rect 4284 28018 4340 28030
rect 4060 27794 4116 27804
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4060 27188 4116 27198
rect 5516 27188 5572 31052
rect 6076 30996 6132 31006
rect 6188 30996 6244 33070
rect 6076 30994 6244 30996
rect 6076 30942 6078 30994
rect 6130 30942 6244 30994
rect 6076 30940 6244 30942
rect 6076 30930 6132 30940
rect 5628 30884 5684 30894
rect 5628 30212 5684 30828
rect 6188 30884 6244 30940
rect 6188 30818 6244 30828
rect 6524 33964 6636 34020
rect 5628 30118 5684 30156
rect 6076 30210 6132 30222
rect 6076 30158 6078 30210
rect 6130 30158 6132 30210
rect 6076 30100 6132 30158
rect 6076 30034 6132 30044
rect 5628 28756 5684 28766
rect 5628 28662 5684 28700
rect 6300 28644 6356 28654
rect 6300 28550 6356 28588
rect 5964 28532 6020 28542
rect 5964 27972 6020 28476
rect 5628 27188 5684 27198
rect 5516 27186 5684 27188
rect 5516 27134 5630 27186
rect 5682 27134 5684 27186
rect 5516 27132 5684 27134
rect 4060 27094 4116 27132
rect 5628 27122 5684 27132
rect 5964 27186 6020 27916
rect 5964 27134 5966 27186
rect 6018 27134 6020 27186
rect 5964 27122 6020 27134
rect 6076 27860 6132 27870
rect 4732 26852 4788 26862
rect 3164 26450 3220 26460
rect 3948 26516 4004 26526
rect 3052 26404 3108 26414
rect 3052 25394 3108 26348
rect 3052 25342 3054 25394
rect 3106 25342 3108 25394
rect 3052 25330 3108 25342
rect 3948 24946 4004 26460
rect 4732 26290 4788 26796
rect 4732 26238 4734 26290
rect 4786 26238 4788 26290
rect 4732 26226 4788 26238
rect 5180 26292 5236 26302
rect 5180 26198 5236 26236
rect 5628 26292 5684 26302
rect 5628 26198 5684 26236
rect 6076 26290 6132 27804
rect 6524 27858 6580 33964
rect 6636 33954 6692 33964
rect 7532 34020 7588 34030
rect 7532 33926 7588 33964
rect 6748 33908 6804 33918
rect 6636 28644 6692 28654
rect 6636 28550 6692 28588
rect 6748 28420 6804 33852
rect 6972 32676 7028 32686
rect 6972 32582 7028 32620
rect 7980 32450 8036 32462
rect 7980 32398 7982 32450
rect 8034 32398 8036 32450
rect 7196 30884 7252 30894
rect 7196 29428 7252 30828
rect 7532 30882 7588 30894
rect 7532 30830 7534 30882
rect 7586 30830 7588 30882
rect 7532 29876 7588 30830
rect 7980 30884 8036 32398
rect 8652 31778 8708 34974
rect 9884 34972 9996 35028
rect 8652 31726 8654 31778
rect 8706 31726 8708 31778
rect 8652 31714 8708 31726
rect 8876 33458 8932 33470
rect 8876 33406 8878 33458
rect 8930 33406 8932 33458
rect 7980 30818 8036 30828
rect 8540 31106 8596 31118
rect 8540 31054 8542 31106
rect 8594 31054 8596 31106
rect 7532 29810 7588 29820
rect 8428 29876 8484 29886
rect 7196 29362 7252 29372
rect 7532 29650 7588 29662
rect 7532 29598 7534 29650
rect 7586 29598 7588 29650
rect 7420 29316 7476 29326
rect 6524 27806 6526 27858
rect 6578 27806 6580 27858
rect 6524 27794 6580 27806
rect 6636 28364 6804 28420
rect 6972 28644 7028 28654
rect 6412 26962 6468 26974
rect 6412 26910 6414 26962
rect 6466 26910 6468 26962
rect 6412 26908 6468 26910
rect 6636 26908 6692 28364
rect 6972 27074 7028 28588
rect 7420 28644 7476 29260
rect 7532 28754 7588 29598
rect 8204 29652 8260 29662
rect 8204 29558 8260 29596
rect 7532 28702 7534 28754
rect 7586 28702 7588 28754
rect 7532 28690 7588 28702
rect 8316 29428 8372 29438
rect 7420 28550 7476 28588
rect 8316 28642 8372 29372
rect 8316 28590 8318 28642
rect 8370 28590 8372 28642
rect 8316 28082 8372 28590
rect 8316 28030 8318 28082
rect 8370 28030 8372 28082
rect 8316 28018 8372 28030
rect 7196 27860 7252 27870
rect 7196 27858 8036 27860
rect 7196 27806 7198 27858
rect 7250 27806 8036 27858
rect 7196 27804 8036 27806
rect 7196 27794 7252 27804
rect 6972 27022 6974 27074
rect 7026 27022 7028 27074
rect 6412 26852 6692 26908
rect 6748 26962 6804 26974
rect 6748 26910 6750 26962
rect 6802 26910 6804 26962
rect 6412 26786 6468 26796
rect 6076 26238 6078 26290
rect 6130 26238 6132 26290
rect 6076 26226 6132 26238
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4732 25732 4788 25742
rect 4060 25620 4116 25630
rect 4060 25526 4116 25564
rect 3948 24894 3950 24946
rect 4002 24894 4004 24946
rect 3948 24882 4004 24894
rect 4060 25284 4116 25294
rect 2044 24836 2100 24846
rect 2044 24834 3220 24836
rect 2044 24782 2046 24834
rect 2098 24782 3220 24834
rect 2044 24780 3220 24782
rect 2044 24770 2100 24780
rect 1820 24722 1876 24734
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 24612 1876 24670
rect 2492 24612 2548 24622
rect 1820 24610 2660 24612
rect 1820 24558 2494 24610
rect 2546 24558 2660 24610
rect 1820 24556 2660 24558
rect 2492 24546 2548 24556
rect 2044 24388 2100 24398
rect 2044 23938 2100 24332
rect 2044 23886 2046 23938
rect 2098 23886 2100 23938
rect 2044 23154 2100 23886
rect 2268 23828 2324 23838
rect 2268 23826 2436 23828
rect 2268 23774 2270 23826
rect 2322 23774 2436 23826
rect 2268 23772 2436 23774
rect 2268 23762 2324 23772
rect 2044 23102 2046 23154
rect 2098 23102 2100 23154
rect 1932 23044 1988 23054
rect 1820 23042 1988 23044
rect 1820 22990 1934 23042
rect 1986 22990 1988 23042
rect 1820 22988 1988 22990
rect 1708 21362 1764 21374
rect 1708 21310 1710 21362
rect 1762 21310 1764 21362
rect 1708 18564 1764 21310
rect 1820 20244 1876 22988
rect 1932 22978 1988 22988
rect 1820 20178 1876 20188
rect 2044 22370 2100 23102
rect 2044 22318 2046 22370
rect 2098 22318 2100 22370
rect 2044 20802 2100 22318
rect 2044 20750 2046 20802
rect 2098 20750 2100 20802
rect 1932 19794 1988 19806
rect 1932 19742 1934 19794
rect 1986 19742 1988 19794
rect 1932 19572 1988 19742
rect 1932 19506 1988 19516
rect 1708 18498 1764 18508
rect 2044 19234 2100 20750
rect 2044 19182 2046 19234
rect 2098 19182 2100 19234
rect 1596 18228 1652 18238
rect 1484 18226 1652 18228
rect 1484 18174 1598 18226
rect 1650 18174 1652 18226
rect 1484 18172 1652 18174
rect 1484 12852 1540 18172
rect 1596 18162 1652 18172
rect 2044 17668 2100 19182
rect 2156 22482 2212 22494
rect 2156 22430 2158 22482
rect 2210 22430 2212 22482
rect 2156 18674 2212 22430
rect 2268 20690 2324 20702
rect 2268 20638 2270 20690
rect 2322 20638 2324 20690
rect 2268 19348 2324 20638
rect 2380 20244 2436 23772
rect 2492 23604 2548 23614
rect 2492 21810 2548 23548
rect 2604 23380 2660 24556
rect 3052 23828 3108 23838
rect 3052 23734 3108 23772
rect 2604 23314 2660 23324
rect 2604 23156 2660 23166
rect 2604 23062 2660 23100
rect 2940 23154 2996 23166
rect 2940 23102 2942 23154
rect 2994 23102 2996 23154
rect 2492 21758 2494 21810
rect 2546 21758 2548 21810
rect 2492 21746 2548 21758
rect 2828 22932 2884 22942
rect 2492 20244 2548 20254
rect 2380 20242 2548 20244
rect 2380 20190 2494 20242
rect 2546 20190 2548 20242
rect 2380 20188 2548 20190
rect 2492 20178 2548 20188
rect 2492 19572 2548 19582
rect 2548 19516 2772 19572
rect 2492 19506 2548 19516
rect 2268 19292 2436 19348
rect 2268 19124 2324 19134
rect 2268 19030 2324 19068
rect 2380 18788 2436 19292
rect 2156 18622 2158 18674
rect 2210 18622 2212 18674
rect 2156 18610 2212 18622
rect 2268 18732 2436 18788
rect 2268 18452 2324 18732
rect 1932 17666 2100 17668
rect 1932 17614 2046 17666
rect 2098 17614 2100 17666
rect 1932 17612 2100 17614
rect 1596 16658 1652 16670
rect 1596 16606 1598 16658
rect 1650 16606 1652 16658
rect 1596 14756 1652 16606
rect 1932 16210 1988 17612
rect 2044 17602 2100 17612
rect 2156 18396 2324 18452
rect 2156 17106 2212 18396
rect 2268 17556 2324 17566
rect 2268 17554 2548 17556
rect 2268 17502 2270 17554
rect 2322 17502 2548 17554
rect 2268 17500 2548 17502
rect 2268 17490 2324 17500
rect 2156 17054 2158 17106
rect 2210 17054 2212 17106
rect 2156 17042 2212 17054
rect 1932 16158 1934 16210
rect 1986 16158 1988 16210
rect 1932 16146 1988 16158
rect 2044 16996 2100 17006
rect 1932 15540 1988 15550
rect 2044 15540 2100 16940
rect 1932 15538 2100 15540
rect 1932 15486 1934 15538
rect 1986 15486 2100 15538
rect 1932 15484 2100 15486
rect 2268 15986 2324 15998
rect 2268 15934 2270 15986
rect 2322 15934 2324 15986
rect 1932 15474 1988 15484
rect 1596 14690 1652 14700
rect 1932 15314 1988 15326
rect 1932 15262 1934 15314
rect 1986 15262 1988 15314
rect 1932 14418 1988 15262
rect 1932 14366 1934 14418
rect 1986 14366 1988 14418
rect 1932 14308 1988 14366
rect 1932 14242 1988 14252
rect 2044 14306 2100 14318
rect 2044 14254 2046 14306
rect 2098 14254 2100 14306
rect 1932 13748 1988 13758
rect 1484 12786 1540 12796
rect 1820 13746 1988 13748
rect 1820 13694 1934 13746
rect 1986 13694 1988 13746
rect 1820 13692 1988 13694
rect 1820 13524 1876 13692
rect 1932 13682 1988 13692
rect 1596 11954 1652 11966
rect 1596 11902 1598 11954
rect 1650 11902 1652 11954
rect 1596 11284 1652 11902
rect 1596 11218 1652 11228
rect 1820 10610 1876 13468
rect 2044 11956 2100 14254
rect 2268 12402 2324 15934
rect 2492 15148 2548 17500
rect 2716 15986 2772 19516
rect 2828 19122 2884 22876
rect 2828 19070 2830 19122
rect 2882 19070 2884 19122
rect 2828 19058 2884 19070
rect 2716 15934 2718 15986
rect 2770 15934 2772 15986
rect 2716 15922 2772 15934
rect 2940 15764 2996 23102
rect 3052 22260 3108 22270
rect 3052 22166 3108 22204
rect 3052 20692 3108 20702
rect 3052 20598 3108 20636
rect 3052 18228 3108 18238
rect 3052 17554 3108 18172
rect 3052 17502 3054 17554
rect 3106 17502 3108 17554
rect 3052 17490 3108 17502
rect 2380 15092 2548 15148
rect 2604 15708 2996 15764
rect 2604 15202 2660 15708
rect 2604 15150 2606 15202
rect 2658 15150 2660 15202
rect 2604 15138 2660 15150
rect 3164 15148 3220 24780
rect 3500 24722 3556 24734
rect 3500 24670 3502 24722
rect 3554 24670 3556 24722
rect 3500 24612 3556 24670
rect 3500 24546 3556 24556
rect 3612 24610 3668 24622
rect 3612 24558 3614 24610
rect 3666 24558 3668 24610
rect 3612 23604 3668 24558
rect 4060 24050 4116 25228
rect 4732 24946 4788 25676
rect 6748 25732 6804 26910
rect 6748 25666 6804 25676
rect 6972 26180 7028 27022
rect 6972 25618 7028 26124
rect 6972 25566 6974 25618
rect 7026 25566 7028 25618
rect 6972 25554 7028 25566
rect 7980 27074 8036 27804
rect 7980 27022 7982 27074
rect 8034 27022 8036 27074
rect 7980 26292 8036 27022
rect 8428 27076 8484 29820
rect 8540 28420 8596 31054
rect 8652 29986 8708 29998
rect 8652 29934 8654 29986
rect 8706 29934 8708 29986
rect 8652 29650 8708 29934
rect 8652 29598 8654 29650
rect 8706 29598 8708 29650
rect 8652 29586 8708 29598
rect 8764 29316 8820 29326
rect 8764 29222 8820 29260
rect 8764 28644 8820 28654
rect 8876 28644 8932 33406
rect 9660 33236 9716 33246
rect 9324 33234 9716 33236
rect 9324 33182 9662 33234
rect 9714 33182 9716 33234
rect 9324 33180 9716 33182
rect 8988 32450 9044 32462
rect 8988 32398 8990 32450
rect 9042 32398 9044 32450
rect 8988 31780 9044 32398
rect 9212 31780 9268 31790
rect 8988 31724 9212 31780
rect 9212 31686 9268 31724
rect 9212 30212 9268 30222
rect 9324 30212 9380 33180
rect 9660 33170 9716 33180
rect 9436 32676 9492 32686
rect 9436 32582 9492 32620
rect 9212 30210 9380 30212
rect 9212 30158 9214 30210
rect 9266 30158 9380 30210
rect 9212 30156 9380 30158
rect 9548 31780 9604 31790
rect 9548 30210 9604 31724
rect 9548 30158 9550 30210
rect 9602 30158 9604 30210
rect 9212 30146 9268 30156
rect 9548 29988 9604 30158
rect 9884 30210 9940 34972
rect 9996 34962 10052 34972
rect 11452 35026 11508 35038
rect 11452 34974 11454 35026
rect 11506 34974 11508 35026
rect 11340 34018 11396 34030
rect 11340 33966 11342 34018
rect 11394 33966 11396 34018
rect 9996 33348 10052 33358
rect 9996 31778 10052 33292
rect 10892 33234 10948 33246
rect 10892 33182 10894 33234
rect 10946 33182 10948 33234
rect 10220 32676 10276 32686
rect 10220 32674 10836 32676
rect 10220 32622 10222 32674
rect 10274 32622 10836 32674
rect 10220 32620 10836 32622
rect 10220 32610 10276 32620
rect 9996 31726 9998 31778
rect 10050 31726 10052 31778
rect 9996 31714 10052 31726
rect 10780 31106 10836 32620
rect 10780 31054 10782 31106
rect 10834 31054 10836 31106
rect 10780 31042 10836 31054
rect 9884 30158 9886 30210
rect 9938 30158 9940 30210
rect 9884 30146 9940 30158
rect 9996 30996 10052 31006
rect 9996 29988 10052 30940
rect 9548 29932 10052 29988
rect 10108 30884 10164 30894
rect 9660 29428 9716 29932
rect 9660 29334 9716 29372
rect 10108 29426 10164 30828
rect 10108 29374 10110 29426
rect 10162 29374 10164 29426
rect 10108 29362 10164 29374
rect 10444 30884 10500 30894
rect 8764 28642 8932 28644
rect 8764 28590 8766 28642
rect 8818 28590 8932 28642
rect 8764 28588 8932 28590
rect 8764 28578 8820 28588
rect 9884 28420 9940 28430
rect 8540 28364 8932 28420
rect 8652 27860 8708 27870
rect 8540 27076 8596 27086
rect 8428 27074 8596 27076
rect 8428 27022 8542 27074
rect 8594 27022 8596 27074
rect 8428 27020 8596 27022
rect 8540 27010 8596 27020
rect 8540 26516 8596 26526
rect 8540 26422 8596 26460
rect 4732 24894 4734 24946
rect 4786 24894 4788 24946
rect 4732 24882 4788 24894
rect 6972 24722 7028 24734
rect 6972 24670 6974 24722
rect 7026 24670 7028 24722
rect 5964 24612 6020 24622
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4060 23998 4062 24050
rect 4114 23998 4116 24050
rect 4060 23986 4116 23998
rect 5628 23828 5684 23838
rect 3612 23538 3668 23548
rect 5516 23826 5684 23828
rect 5516 23774 5630 23826
rect 5682 23774 5684 23826
rect 5516 23772 5684 23774
rect 3500 23380 3556 23390
rect 3388 18564 3444 18574
rect 3388 15426 3444 18508
rect 3500 17556 3556 23324
rect 5516 23378 5572 23772
rect 5628 23762 5684 23772
rect 5964 23826 6020 24556
rect 6860 24164 6916 24174
rect 5964 23774 5966 23826
rect 6018 23774 6020 23826
rect 5516 23326 5518 23378
rect 5570 23326 5572 23378
rect 5516 23314 5572 23326
rect 5516 23156 5572 23166
rect 5964 23156 6020 23774
rect 6636 23826 6692 23838
rect 6636 23774 6638 23826
rect 6690 23774 6692 23826
rect 6636 23716 6692 23774
rect 6636 23650 6692 23660
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4060 22484 4116 22494
rect 4060 22390 4116 22428
rect 5516 22372 5572 23100
rect 5404 22370 5572 22372
rect 5404 22318 5518 22370
rect 5570 22318 5572 22370
rect 5404 22316 5572 22318
rect 3836 21924 3892 21934
rect 3836 20914 3892 21868
rect 4732 21588 4788 21598
rect 3836 20862 3838 20914
rect 3890 20862 3892 20914
rect 3836 20850 3892 20862
rect 4060 21586 4788 21588
rect 4060 21534 4734 21586
rect 4786 21534 4788 21586
rect 4060 21532 4788 21534
rect 3836 20580 3892 20590
rect 3836 19346 3892 20524
rect 3836 19294 3838 19346
rect 3890 19294 3892 19346
rect 3836 19282 3892 19294
rect 3948 19348 4004 19358
rect 3948 17778 4004 19292
rect 3948 17726 3950 17778
rect 4002 17726 4004 17778
rect 3948 17714 4004 17726
rect 3500 17490 3556 17500
rect 4060 16210 4116 21532
rect 4732 21522 4788 21532
rect 5404 21586 5460 22316
rect 5516 22306 5572 22316
rect 5852 23100 6244 23156
rect 5404 21534 5406 21586
rect 5458 21534 5460 21586
rect 5404 21476 5460 21534
rect 5852 21586 5908 23100
rect 6188 23044 6244 23100
rect 6524 23044 6580 23054
rect 6188 23042 6580 23044
rect 6188 22990 6526 23042
rect 6578 22990 6580 23042
rect 6188 22988 6580 22990
rect 6524 22978 6580 22988
rect 6076 22932 6132 22942
rect 6076 22838 6132 22876
rect 6748 22708 6804 22718
rect 6076 22372 6132 22382
rect 5852 21534 5854 21586
rect 5906 21534 5908 21586
rect 5852 21522 5908 21534
rect 5964 22370 6132 22372
rect 5964 22318 6078 22370
rect 6130 22318 6132 22370
rect 5964 22316 6132 22318
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5404 20804 5460 21420
rect 5516 20804 5572 20814
rect 5404 20802 5572 20804
rect 5404 20750 5518 20802
rect 5570 20750 5572 20802
rect 5404 20748 5572 20750
rect 5516 20188 5572 20748
rect 5404 20132 5572 20188
rect 4956 20020 5012 20030
rect 4060 16158 4062 16210
rect 4114 16158 4116 16210
rect 4060 16146 4116 16158
rect 4172 20018 5012 20020
rect 4172 19966 4958 20018
rect 5010 19966 5012 20018
rect 4172 19964 5012 19966
rect 4172 15988 4228 19964
rect 4956 19954 5012 19964
rect 5404 20018 5460 20132
rect 5404 19966 5406 20018
rect 5458 19966 5460 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4732 18452 4788 18462
rect 5292 18452 5348 18462
rect 5404 18452 5460 19966
rect 5964 19348 6020 22316
rect 6076 22306 6132 22316
rect 6076 22148 6132 22158
rect 6076 21698 6132 22092
rect 6076 21646 6078 21698
rect 6130 21646 6132 21698
rect 6076 21634 6132 21646
rect 6636 21476 6692 21486
rect 6636 21382 6692 21420
rect 6188 20802 6244 20814
rect 6188 20750 6190 20802
rect 6242 20750 6244 20802
rect 5964 19282 6020 19292
rect 6076 19684 6132 19694
rect 5964 19124 6020 19134
rect 5964 18674 6020 19068
rect 6076 19122 6132 19628
rect 6076 19070 6078 19122
rect 6130 19070 6132 19122
rect 6076 19058 6132 19070
rect 5964 18622 5966 18674
rect 6018 18622 6020 18674
rect 5964 18610 6020 18622
rect 4732 18450 4900 18452
rect 4732 18398 4734 18450
rect 4786 18398 4900 18450
rect 4732 18396 4900 18398
rect 4732 18386 4788 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 16884 4676 16894
rect 3388 15374 3390 15426
rect 3442 15374 3444 15426
rect 3388 15362 3444 15374
rect 3724 15932 4228 15988
rect 4284 16882 4676 16884
rect 4284 16830 4622 16882
rect 4674 16830 4676 16882
rect 4284 16828 4676 16830
rect 2940 15092 3220 15148
rect 2380 13972 2436 15092
rect 2716 14308 2772 14318
rect 2716 14214 2772 14252
rect 2380 13906 2436 13916
rect 2604 13746 2660 13758
rect 2604 13694 2606 13746
rect 2658 13694 2660 13746
rect 2380 12852 2436 12862
rect 2380 12758 2436 12796
rect 2604 12628 2660 13694
rect 2604 12562 2660 12572
rect 2268 12350 2270 12402
rect 2322 12350 2324 12402
rect 2268 12338 2324 12350
rect 2044 11890 2100 11900
rect 2380 11284 2436 11294
rect 2380 11190 2436 11228
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 10546 1876 10558
rect 2268 10612 2324 10622
rect 2940 10612 2996 15092
rect 3164 14308 3220 14318
rect 3164 13636 3220 14252
rect 3164 13570 3220 13580
rect 3724 13074 3780 15932
rect 3724 13022 3726 13074
rect 3778 13022 3780 13074
rect 3724 13010 3780 13022
rect 3836 14642 3892 14654
rect 3836 14590 3838 14642
rect 3890 14590 3892 14642
rect 3500 12628 3556 12638
rect 3500 11506 3556 12572
rect 3836 12180 3892 14590
rect 4284 13188 4340 16828
rect 4620 16818 4676 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16324 4900 18396
rect 5292 18450 5460 18452
rect 5292 18398 5294 18450
rect 5346 18398 5460 18450
rect 5292 18396 5460 18398
rect 5292 18386 5348 18396
rect 5404 18228 5460 18238
rect 5404 18134 5460 18172
rect 5068 17442 5124 17454
rect 5068 17390 5070 17442
rect 5122 17390 5124 17442
rect 4844 16258 4900 16268
rect 4956 16884 5012 16894
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4956 14418 5012 16828
rect 4956 14366 4958 14418
rect 5010 14366 5012 14418
rect 4956 14354 5012 14366
rect 5068 16884 5124 17390
rect 5852 17442 5908 17454
rect 5852 17390 5854 17442
rect 5906 17390 5908 17442
rect 5404 16884 5460 16894
rect 5068 16882 5460 16884
rect 5068 16830 5070 16882
rect 5122 16830 5406 16882
rect 5458 16830 5460 16882
rect 5068 16828 5460 16830
rect 5068 15316 5124 16828
rect 5404 16818 5460 16828
rect 5740 15876 5796 15886
rect 5852 15876 5908 17390
rect 6076 16882 6132 16894
rect 6076 16830 6078 16882
rect 6130 16830 6132 16882
rect 6076 16100 6132 16830
rect 6188 16212 6244 20750
rect 6748 19684 6804 22652
rect 6748 19618 6804 19628
rect 6860 19346 6916 24108
rect 6972 20580 7028 24670
rect 7644 24724 7700 24734
rect 7644 24630 7700 24668
rect 7980 24724 8036 26236
rect 8540 25732 8596 25742
rect 8540 25506 8596 25676
rect 8540 25454 8542 25506
rect 8594 25454 8596 25506
rect 8540 25442 8596 25454
rect 8652 25284 8708 27804
rect 8876 26908 8932 28364
rect 9884 27746 9940 28364
rect 10444 28420 10500 30828
rect 10892 30772 10948 33182
rect 11004 30994 11060 31006
rect 11004 30942 11006 30994
rect 11058 30942 11060 30994
rect 11004 30884 11060 30942
rect 11340 30884 11396 33966
rect 11452 33348 11508 34974
rect 12684 34802 12740 34814
rect 12684 34750 12686 34802
rect 12738 34750 12740 34802
rect 12348 34018 12404 34030
rect 12348 33966 12350 34018
rect 12402 33966 12404 34018
rect 12348 33570 12404 33966
rect 12348 33518 12350 33570
rect 12402 33518 12404 33570
rect 12348 33506 12404 33518
rect 12572 34018 12628 34030
rect 12572 33966 12574 34018
rect 12626 33966 12628 34018
rect 11900 33458 11956 33470
rect 11900 33406 11902 33458
rect 11954 33406 11956 33458
rect 11900 33348 11956 33406
rect 11900 33292 12516 33348
rect 11452 33282 11508 33292
rect 12348 33124 12404 33134
rect 12236 33122 12404 33124
rect 12236 33070 12350 33122
rect 12402 33070 12404 33122
rect 12236 33068 12404 33070
rect 12124 30996 12180 31006
rect 11452 30884 11508 30894
rect 11340 30828 11452 30884
rect 11004 30818 11060 30828
rect 11452 30790 11508 30828
rect 11676 30882 11732 30894
rect 11676 30830 11678 30882
rect 11730 30830 11732 30882
rect 10892 30706 10948 30716
rect 11676 29652 11732 30830
rect 11676 29586 11732 29596
rect 11788 30772 11844 30782
rect 11788 28866 11844 30716
rect 11788 28814 11790 28866
rect 11842 28814 11844 28866
rect 11788 28802 11844 28814
rect 10444 28354 10500 28364
rect 11228 28644 11284 28654
rect 11228 28418 11284 28588
rect 12012 28644 12068 28654
rect 12012 28550 12068 28588
rect 11228 28366 11230 28418
rect 11282 28366 11284 28418
rect 11228 28354 11284 28366
rect 12124 28532 12180 30940
rect 12236 30884 12292 33068
rect 12348 33058 12404 33068
rect 12460 32562 12516 33292
rect 12460 32510 12462 32562
rect 12514 32510 12516 32562
rect 12460 32498 12516 32510
rect 12236 30818 12292 30828
rect 12348 31554 12404 31566
rect 12348 31502 12350 31554
rect 12402 31502 12404 31554
rect 12348 30212 12404 31502
rect 12572 30994 12628 33966
rect 12572 30942 12574 30994
rect 12626 30942 12628 30994
rect 12572 30930 12628 30942
rect 12348 30146 12404 30156
rect 12460 30100 12516 30110
rect 12460 29986 12516 30044
rect 12460 29934 12462 29986
rect 12514 29934 12516 29986
rect 12460 29922 12516 29934
rect 12684 29988 12740 34750
rect 12796 31892 12852 37324
rect 13804 37380 13860 37390
rect 13804 37286 13860 37324
rect 15148 37154 15204 37166
rect 15148 37102 15150 37154
rect 15202 37102 15204 37154
rect 14812 36596 14868 36606
rect 13916 36594 14868 36596
rect 13916 36542 14814 36594
rect 14866 36542 14868 36594
rect 13916 36540 14868 36542
rect 13244 34356 13300 34366
rect 12908 33570 12964 33582
rect 12908 33518 12910 33570
rect 12962 33518 12964 33570
rect 12908 33122 12964 33518
rect 12908 33070 12910 33122
rect 12962 33070 12964 33122
rect 12908 32564 12964 33070
rect 13244 32786 13300 34300
rect 13580 34242 13636 34254
rect 13580 34190 13582 34242
rect 13634 34190 13636 34242
rect 13244 32734 13246 32786
rect 13298 32734 13300 32786
rect 13244 32722 13300 32734
rect 13356 33348 13412 33358
rect 13468 33348 13524 33358
rect 13356 33346 13468 33348
rect 13356 33294 13358 33346
rect 13410 33294 13468 33346
rect 13356 33292 13468 33294
rect 13132 32564 13188 32574
rect 13356 32564 13412 33292
rect 13468 33282 13524 33292
rect 12908 32562 13412 32564
rect 12908 32510 13134 32562
rect 13186 32510 13412 32562
rect 12908 32508 13412 32510
rect 13020 31892 13076 31902
rect 12796 31890 13076 31892
rect 12796 31838 13022 31890
rect 13074 31838 13076 31890
rect 12796 31836 13076 31838
rect 13020 31826 13076 31836
rect 13132 31780 13188 32508
rect 13356 31780 13412 31790
rect 13132 31778 13412 31780
rect 13132 31726 13358 31778
rect 13410 31726 13412 31778
rect 13132 31724 13412 31726
rect 13356 30996 13412 31724
rect 13356 30930 13412 30940
rect 13580 30772 13636 34190
rect 13916 31778 13972 36540
rect 14812 36530 14868 36540
rect 14700 35588 14756 35598
rect 14476 35586 14756 35588
rect 14476 35534 14702 35586
rect 14754 35534 14756 35586
rect 14476 35532 14756 35534
rect 14028 35252 14084 35262
rect 14028 33346 14084 35196
rect 14364 34020 14420 34030
rect 14028 33294 14030 33346
rect 14082 33294 14084 33346
rect 14028 33282 14084 33294
rect 14140 34018 14420 34020
rect 14140 33966 14366 34018
rect 14418 33966 14420 34018
rect 14140 33964 14420 33966
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 13916 31714 13972 31726
rect 14028 32674 14084 32686
rect 14028 32622 14030 32674
rect 14082 32622 14084 32674
rect 13020 30716 13636 30772
rect 13020 30210 13076 30716
rect 14028 30660 14084 32622
rect 14028 30594 14084 30604
rect 13020 30158 13022 30210
rect 13074 30158 13076 30210
rect 13020 30146 13076 30158
rect 13692 30210 13748 30222
rect 13692 30158 13694 30210
rect 13746 30158 13748 30210
rect 13468 30100 13524 30110
rect 13468 30006 13524 30044
rect 12684 29932 13188 29988
rect 12348 29652 12404 29662
rect 12348 29558 12404 29596
rect 13132 29650 13188 29932
rect 13132 29598 13134 29650
rect 13186 29598 13188 29650
rect 13132 29586 13188 29598
rect 13356 29426 13412 29438
rect 13356 29374 13358 29426
rect 13410 29374 13412 29426
rect 10108 27860 10164 27870
rect 10108 27766 10164 27804
rect 9884 27694 9886 27746
rect 9938 27694 9940 27746
rect 9772 27188 9828 27198
rect 8876 26852 9156 26908
rect 9100 26514 9156 26852
rect 9100 26462 9102 26514
rect 9154 26462 9156 26514
rect 9100 26450 9156 26462
rect 9660 26516 9716 26554
rect 9660 26450 9716 26460
rect 9660 26292 9716 26302
rect 9548 26180 9604 26190
rect 9548 26086 9604 26124
rect 7980 24658 8036 24668
rect 8428 25228 8708 25284
rect 8988 25732 9044 25742
rect 8988 25282 9044 25676
rect 9548 25508 9604 25518
rect 9660 25508 9716 26236
rect 9548 25506 9716 25508
rect 9548 25454 9550 25506
rect 9602 25454 9716 25506
rect 9548 25452 9716 25454
rect 9548 25442 9604 25452
rect 8988 25230 8990 25282
rect 9042 25230 9044 25282
rect 7868 24050 7924 24062
rect 7868 23998 7870 24050
rect 7922 23998 7924 24050
rect 7868 23940 7924 23998
rect 8428 24052 8484 25228
rect 8428 24050 8596 24052
rect 8428 23998 8430 24050
rect 8482 23998 8596 24050
rect 8428 23996 8596 23998
rect 8428 23986 8484 23996
rect 7868 23874 7924 23884
rect 8428 22148 8484 22158
rect 8428 22054 8484 22092
rect 6972 20514 7028 20524
rect 7756 22036 7812 22046
rect 6860 19294 6862 19346
rect 6914 19294 6916 19346
rect 6860 19282 6916 19294
rect 7644 20020 7700 20030
rect 7644 19346 7700 19964
rect 7644 19294 7646 19346
rect 7698 19294 7700 19346
rect 7644 19282 7700 19294
rect 6636 17666 6692 17678
rect 6636 17614 6638 17666
rect 6690 17614 6692 17666
rect 6636 17444 6692 17614
rect 6636 17378 6692 17388
rect 6972 16660 7028 16670
rect 6636 16212 6692 16222
rect 6188 16210 6692 16212
rect 6188 16158 6638 16210
rect 6690 16158 6692 16210
rect 6188 16156 6692 16158
rect 6636 16146 6692 16156
rect 6076 16044 6468 16100
rect 6300 15876 6356 15886
rect 5740 15874 6300 15876
rect 5740 15822 5742 15874
rect 5794 15822 6300 15874
rect 5740 15820 6300 15822
rect 4844 13972 4900 13982
rect 4844 13878 4900 13916
rect 5068 13524 5124 15260
rect 5628 15314 5684 15326
rect 5628 15262 5630 15314
rect 5682 15262 5684 15314
rect 5628 15092 5684 15262
rect 5740 15316 5796 15820
rect 6300 15782 6356 15820
rect 5740 15250 5796 15260
rect 5628 15036 6020 15092
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4396 13188 4452 13198
rect 4284 13132 4396 13188
rect 4396 13122 4452 13132
rect 5068 12404 5124 13468
rect 5516 14306 5572 14318
rect 5516 14254 5518 14306
rect 5570 14254 5572 14306
rect 5516 12628 5572 14254
rect 5852 13636 5908 13646
rect 5852 13542 5908 13580
rect 5628 13522 5684 13534
rect 5628 13470 5630 13522
rect 5682 13470 5684 13522
rect 5628 13076 5684 13470
rect 5628 13010 5684 13020
rect 5740 12740 5796 12750
rect 5516 12562 5572 12572
rect 5628 12738 5908 12740
rect 5628 12686 5742 12738
rect 5794 12686 5908 12738
rect 5628 12684 5908 12686
rect 5628 12404 5684 12684
rect 5740 12674 5796 12684
rect 5068 12402 5684 12404
rect 5068 12350 5630 12402
rect 5682 12350 5684 12402
rect 5068 12348 5684 12350
rect 4620 12180 4676 12190
rect 3836 12178 4676 12180
rect 3836 12126 4622 12178
rect 4674 12126 4676 12178
rect 3836 12124 4676 12126
rect 4620 12114 4676 12124
rect 5068 12178 5124 12348
rect 5628 12338 5684 12348
rect 5068 12126 5070 12178
rect 5122 12126 5124 12178
rect 5068 12114 5124 12126
rect 4284 11956 4340 11966
rect 4284 11620 4340 11900
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4284 11564 4564 11620
rect 3500 11454 3502 11506
rect 3554 11454 3556 11506
rect 3500 11442 3556 11454
rect 4508 10834 4564 11564
rect 4508 10782 4510 10834
rect 4562 10782 4564 10834
rect 4508 10770 4564 10782
rect 2268 10610 2996 10612
rect 2268 10558 2270 10610
rect 2322 10558 2996 10610
rect 2268 10556 2996 10558
rect 2268 10546 2324 10556
rect 5292 10386 5348 10398
rect 5292 10334 5294 10386
rect 5346 10334 5348 10386
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 5292 9716 5348 10334
rect 5852 9938 5908 12684
rect 5964 10498 6020 15036
rect 6188 14306 6244 14318
rect 6188 14254 6190 14306
rect 6242 14254 6244 14306
rect 6188 13858 6244 14254
rect 6188 13806 6190 13858
rect 6242 13806 6244 13858
rect 6188 13794 6244 13806
rect 6412 11506 6468 16044
rect 6524 14756 6580 14766
rect 6524 12850 6580 14700
rect 6972 13858 7028 16604
rect 7756 15986 7812 21980
rect 8540 21586 8596 23996
rect 8876 23716 8932 23726
rect 8988 23716 9044 25230
rect 9324 24724 9380 24734
rect 9660 24724 9716 25452
rect 9380 24722 9716 24724
rect 9380 24670 9662 24722
rect 9714 24670 9716 24722
rect 9380 24668 9716 24670
rect 9324 23938 9380 24668
rect 9660 24658 9716 24668
rect 9324 23886 9326 23938
rect 9378 23886 9380 23938
rect 9324 23874 9380 23886
rect 9660 23940 9716 23950
rect 9772 23940 9828 27132
rect 9884 26908 9940 27694
rect 11788 27746 11844 27758
rect 11788 27694 11790 27746
rect 11842 27694 11844 27746
rect 11676 26964 11732 27002
rect 9884 26852 10276 26908
rect 11676 26898 11732 26908
rect 9884 25508 9940 25518
rect 9884 25414 9940 25452
rect 10108 24722 10164 24734
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 10108 24164 10164 24670
rect 10108 24098 10164 24108
rect 9660 23938 9828 23940
rect 9660 23886 9662 23938
rect 9714 23886 9828 23938
rect 9660 23884 9828 23886
rect 9660 23874 9716 23884
rect 8876 23714 9044 23716
rect 8876 23662 8878 23714
rect 8930 23662 9044 23714
rect 8876 23660 9044 23662
rect 8876 23154 8932 23660
rect 8876 23102 8878 23154
rect 8930 23102 8932 23154
rect 8876 23044 8932 23102
rect 8876 22978 8932 22988
rect 9660 23044 9716 23054
rect 9716 22988 9828 23044
rect 9660 22950 9716 22988
rect 9548 22370 9604 22382
rect 9548 22318 9550 22370
rect 9602 22318 9604 22370
rect 9212 22148 9268 22158
rect 9212 22054 9268 22092
rect 8540 21534 8542 21586
rect 8594 21534 8596 21586
rect 8316 21476 8372 21486
rect 8316 20356 8372 21420
rect 8316 20300 8484 20356
rect 7868 19908 7924 19918
rect 7868 19906 8148 19908
rect 7868 19854 7870 19906
rect 7922 19854 8148 19906
rect 7868 19852 8148 19854
rect 7868 19842 7924 19852
rect 8092 19346 8148 19852
rect 8092 19294 8094 19346
rect 8146 19294 8148 19346
rect 7756 15934 7758 15986
rect 7810 15934 7812 15986
rect 7756 15922 7812 15934
rect 7980 18564 8036 18574
rect 7980 15428 8036 18508
rect 8092 17668 8148 19294
rect 8428 19236 8484 20300
rect 8540 20020 8596 21534
rect 9548 21588 9604 22318
rect 9548 21522 9604 21532
rect 9660 21474 9716 21486
rect 9660 21422 9662 21474
rect 9714 21422 9716 21474
rect 9660 21140 9716 21422
rect 8652 21084 9716 21140
rect 8652 20578 8708 21084
rect 9324 20692 9380 20702
rect 9324 20598 9380 20636
rect 8652 20526 8654 20578
rect 8706 20526 8708 20578
rect 8652 20514 8708 20526
rect 9212 20578 9268 20590
rect 9212 20526 9214 20578
rect 9266 20526 9268 20578
rect 8540 19926 8596 19964
rect 8540 19236 8596 19246
rect 8428 19234 8596 19236
rect 8428 19182 8542 19234
rect 8594 19182 8596 19234
rect 8428 19180 8596 19182
rect 8092 17602 8148 17612
rect 8204 18900 8260 18910
rect 8204 15538 8260 18844
rect 8428 18450 8484 18462
rect 8428 18398 8430 18450
rect 8482 18398 8484 18450
rect 8428 18228 8484 18398
rect 8540 18452 8596 19180
rect 8988 19234 9044 19246
rect 8988 19182 8990 19234
rect 9042 19182 9044 19234
rect 8876 18452 8932 18462
rect 8540 18450 8932 18452
rect 8540 18398 8878 18450
rect 8930 18398 8932 18450
rect 8540 18396 8932 18398
rect 8876 18386 8932 18396
rect 8428 18172 8932 18228
rect 8652 18004 8708 18014
rect 8316 17948 8652 18004
rect 8316 17778 8372 17948
rect 8316 17726 8318 17778
rect 8370 17726 8372 17778
rect 8316 17714 8372 17726
rect 8204 15486 8206 15538
rect 8258 15486 8260 15538
rect 8204 15474 8260 15486
rect 8316 16994 8372 17006
rect 8316 16942 8318 16994
rect 8370 16942 8372 16994
rect 8316 15540 8372 16942
rect 8540 16100 8596 16110
rect 8540 16006 8596 16044
rect 8316 15474 8372 15484
rect 7980 15372 8148 15428
rect 7980 15204 8036 15214
rect 6972 13806 6974 13858
rect 7026 13806 7028 13858
rect 6972 13794 7028 13806
rect 7868 15092 7924 15102
rect 7756 13412 7812 13422
rect 6524 12798 6526 12850
rect 6578 12798 6580 12850
rect 6524 12786 6580 12798
rect 6972 13188 7028 13198
rect 6412 11454 6414 11506
rect 6466 11454 6468 11506
rect 6412 11442 6468 11454
rect 6748 12628 6804 12638
rect 6748 10722 6804 12572
rect 6972 12066 7028 13132
rect 6972 12014 6974 12066
rect 7026 12014 7028 12066
rect 6972 12002 7028 12014
rect 7756 11282 7812 13356
rect 7868 13074 7924 15036
rect 7980 13634 8036 15148
rect 7980 13582 7982 13634
rect 8034 13582 8036 13634
rect 7980 13570 8036 13582
rect 7868 13022 7870 13074
rect 7922 13022 7924 13074
rect 7868 13010 7924 13022
rect 8092 12290 8148 15372
rect 8428 14868 8484 14878
rect 8652 14868 8708 17948
rect 8876 16436 8932 18172
rect 8988 17108 9044 19182
rect 9212 18676 9268 20526
rect 9212 18610 9268 18620
rect 9436 19794 9492 19806
rect 9436 19742 9438 19794
rect 9490 19742 9492 19794
rect 9436 18564 9492 19742
rect 9436 18498 9492 18508
rect 9436 18226 9492 18238
rect 9436 18174 9438 18226
rect 9490 18174 9492 18226
rect 8988 17042 9044 17052
rect 9212 17668 9268 17678
rect 9100 16660 9156 16670
rect 9100 16566 9156 16604
rect 8876 16380 9044 16436
rect 8876 16098 8932 16110
rect 8876 16046 8878 16098
rect 8930 16046 8932 16098
rect 8876 15204 8932 16046
rect 8876 15138 8932 15148
rect 8484 14812 8708 14868
rect 8764 15090 8820 15102
rect 8764 15038 8766 15090
rect 8818 15038 8820 15090
rect 8428 13636 8484 14812
rect 8428 13542 8484 13580
rect 8652 14530 8708 14542
rect 8652 14478 8654 14530
rect 8706 14478 8708 14530
rect 8652 12516 8708 14478
rect 8764 13412 8820 15038
rect 8988 15092 9044 16380
rect 8988 15026 9044 15036
rect 9212 16100 9268 17612
rect 9436 16884 9492 18174
rect 9436 16818 9492 16828
rect 9660 17666 9716 17678
rect 9660 17614 9662 17666
rect 9714 17614 9716 17666
rect 9212 15540 9268 16044
rect 9212 14532 9268 15484
rect 8876 14530 9268 14532
rect 8876 14478 9214 14530
rect 9266 14478 9268 14530
rect 8876 14476 9268 14478
rect 8876 13970 8932 14476
rect 9212 14466 9268 14476
rect 9436 16658 9492 16670
rect 9436 16606 9438 16658
rect 9490 16606 9492 16658
rect 8876 13918 8878 13970
rect 8930 13918 8932 13970
rect 8876 13906 8932 13918
rect 8764 13346 8820 13356
rect 9436 13412 9492 16606
rect 9548 15428 9604 15438
rect 9548 15334 9604 15372
rect 9660 14868 9716 17614
rect 9436 13346 9492 13356
rect 9548 14812 9716 14868
rect 9772 17444 9828 22988
rect 10220 23042 10276 26852
rect 11116 26852 11172 26862
rect 11116 26850 11284 26852
rect 11116 26798 11118 26850
rect 11170 26798 11284 26850
rect 11116 26796 11284 26798
rect 11116 26786 11172 26796
rect 11228 26402 11284 26796
rect 11228 26350 11230 26402
rect 11282 26350 11284 26402
rect 11228 26338 11284 26350
rect 11788 26292 11844 27694
rect 12124 27186 12180 28476
rect 12236 28756 12292 28766
rect 12236 28642 12292 28700
rect 12236 28590 12238 28642
rect 12290 28590 12292 28642
rect 12236 28420 12292 28590
rect 12236 28354 12292 28364
rect 12908 28642 12964 28654
rect 12908 28590 12910 28642
rect 12962 28590 12964 28642
rect 12908 27860 12964 28590
rect 12908 27794 12964 27804
rect 13356 28644 13412 29374
rect 13692 28756 13748 30158
rect 13916 29428 13972 29438
rect 14140 29428 14196 33964
rect 14364 33954 14420 33964
rect 14252 30212 14308 30222
rect 14252 30118 14308 30156
rect 13916 29426 14196 29428
rect 13916 29374 13918 29426
rect 13970 29374 14196 29426
rect 13916 29372 14196 29374
rect 13916 29362 13972 29372
rect 14476 29204 14532 35532
rect 14700 35522 14756 35532
rect 15148 35252 15204 37102
rect 15148 35186 15204 35196
rect 15820 36370 15876 36382
rect 15820 36318 15822 36370
rect 15874 36318 15876 36370
rect 14700 35028 14756 35038
rect 14700 34934 14756 34972
rect 15820 34356 15876 36318
rect 16044 35810 16100 35822
rect 16044 35758 16046 35810
rect 16098 35758 16100 35810
rect 15820 34290 15876 34300
rect 15932 34802 15988 34814
rect 15932 34750 15934 34802
rect 15986 34750 15988 34802
rect 15708 34242 15764 34254
rect 15708 34190 15710 34242
rect 15762 34190 15764 34242
rect 15596 33796 15652 33806
rect 15484 31668 15540 31678
rect 14924 31106 14980 31118
rect 14924 31054 14926 31106
rect 14978 31054 14980 31106
rect 14924 30322 14980 31054
rect 14924 30270 14926 30322
rect 14978 30270 14980 30322
rect 14924 30258 14980 30270
rect 13692 28690 13748 28700
rect 13916 29148 14532 29204
rect 14588 30100 14644 30110
rect 13356 27858 13412 28588
rect 13580 28642 13636 28654
rect 13580 28590 13582 28642
rect 13634 28590 13636 28642
rect 13580 28532 13636 28590
rect 13580 28466 13636 28476
rect 13356 27806 13358 27858
rect 13410 27806 13412 27858
rect 13356 27794 13412 27806
rect 13468 27860 13524 27870
rect 12124 27134 12126 27186
rect 12178 27134 12180 27186
rect 12124 27122 12180 27134
rect 13468 27076 13524 27804
rect 13916 27858 13972 29148
rect 14028 28756 14084 28766
rect 14028 28662 14084 28700
rect 14476 28756 14532 28766
rect 14588 28756 14644 30044
rect 15260 30100 15316 30110
rect 15260 30006 15316 30044
rect 14532 28700 14644 28756
rect 14476 28662 14532 28700
rect 13916 27806 13918 27858
rect 13970 27806 13972 27858
rect 13916 27794 13972 27806
rect 14924 28642 14980 28654
rect 14924 28590 14926 28642
rect 14978 28590 14980 28642
rect 14924 28532 14980 28590
rect 15148 28644 15204 28654
rect 15148 28550 15204 28588
rect 14924 27186 14980 28476
rect 14924 27134 14926 27186
rect 14978 27134 14980 27186
rect 14924 27122 14980 27134
rect 13468 26982 13524 27020
rect 12572 26962 12628 26974
rect 12572 26910 12574 26962
rect 12626 26910 12628 26962
rect 12572 26908 12628 26910
rect 12460 26852 12628 26908
rect 12908 26962 12964 26974
rect 12908 26910 12910 26962
rect 12962 26910 12964 26962
rect 11788 26198 11844 26236
rect 12348 26290 12404 26302
rect 12348 26238 12350 26290
rect 12402 26238 12404 26290
rect 10220 22990 10222 23042
rect 10274 22990 10276 23042
rect 10220 22978 10276 22990
rect 11564 26178 11620 26190
rect 11564 26126 11566 26178
rect 11618 26126 11620 26178
rect 11564 25508 11620 26126
rect 12348 25620 12404 26238
rect 12348 25554 12404 25564
rect 9884 22370 9940 22382
rect 9884 22318 9886 22370
rect 9938 22318 9940 22370
rect 9884 21924 9940 22318
rect 9884 21858 9940 21868
rect 11564 22148 11620 25452
rect 12236 25284 12292 25294
rect 12236 23714 12292 25228
rect 12460 25282 12516 26852
rect 12908 25508 12964 26910
rect 14924 26514 14980 26526
rect 14924 26462 14926 26514
rect 14978 26462 14980 26514
rect 13020 26404 13076 26414
rect 13020 25730 13076 26348
rect 13020 25678 13022 25730
rect 13074 25678 13076 25730
rect 13020 25666 13076 25678
rect 13244 26292 13300 26302
rect 12908 25442 12964 25452
rect 12460 25230 12462 25282
rect 12514 25230 12516 25282
rect 12460 25218 12516 25230
rect 12572 25396 12628 25406
rect 12572 24946 12628 25340
rect 12572 24894 12574 24946
rect 12626 24894 12628 24946
rect 12572 24882 12628 24894
rect 13244 24722 13300 26236
rect 13692 25508 13748 25518
rect 13692 25414 13748 25452
rect 14364 25508 14420 25518
rect 14364 25414 14420 25452
rect 13468 25396 13524 25406
rect 13468 25302 13524 25340
rect 14140 25394 14196 25406
rect 14140 25342 14142 25394
rect 14194 25342 14196 25394
rect 14140 25284 14196 25342
rect 14140 25218 14196 25228
rect 13244 24670 13246 24722
rect 13298 24670 13300 24722
rect 13244 24658 13300 24670
rect 13916 24722 13972 24734
rect 13916 24670 13918 24722
rect 13970 24670 13972 24722
rect 13132 24498 13188 24510
rect 13132 24446 13134 24498
rect 13186 24446 13188 24498
rect 13132 23828 13188 24446
rect 13132 23762 13188 23772
rect 12236 23662 12238 23714
rect 12290 23662 12292 23714
rect 12236 23650 12292 23662
rect 12796 23714 12852 23726
rect 12796 23662 12798 23714
rect 12850 23662 12852 23714
rect 12572 23154 12628 23166
rect 12572 23102 12574 23154
rect 12626 23102 12628 23154
rect 12572 23044 12628 23102
rect 11228 21700 11284 21710
rect 11564 21700 11620 22092
rect 11228 21698 11620 21700
rect 11228 21646 11230 21698
rect 11282 21646 11566 21698
rect 11618 21646 11620 21698
rect 11228 21644 11620 21646
rect 11228 21634 11284 21644
rect 11564 21634 11620 21644
rect 11676 22932 11732 22942
rect 9884 21586 9940 21598
rect 9884 21534 9886 21586
rect 9938 21534 9940 21586
rect 9884 21476 9940 21534
rect 9884 18004 9940 21420
rect 10556 21476 10612 21486
rect 10892 21476 10948 21486
rect 10556 21382 10612 21420
rect 10668 21474 10948 21476
rect 10668 21422 10894 21474
rect 10946 21422 10948 21474
rect 10668 21420 10948 21422
rect 10668 21140 10724 21420
rect 10892 21410 10948 21420
rect 10108 21084 10724 21140
rect 10108 20690 10164 21084
rect 10108 20638 10110 20690
rect 10162 20638 10164 20690
rect 10108 20626 10164 20638
rect 11676 20188 11732 22876
rect 12572 22372 12628 22988
rect 12796 22708 12852 23662
rect 13916 23492 13972 24670
rect 14924 24500 14980 26462
rect 15484 26292 15540 31612
rect 15596 30210 15652 33740
rect 15708 31218 15764 34190
rect 15708 31166 15710 31218
rect 15762 31166 15764 31218
rect 15708 31154 15764 31166
rect 15820 31780 15876 31790
rect 15596 30158 15598 30210
rect 15650 30158 15652 30210
rect 15596 30146 15652 30158
rect 15820 28642 15876 31724
rect 15932 29988 15988 34750
rect 16044 33684 16100 35758
rect 16492 35586 16548 35598
rect 16492 35534 16494 35586
rect 16546 35534 16548 35586
rect 16044 33618 16100 33628
rect 16380 35252 16436 35262
rect 16380 32562 16436 35196
rect 16492 33122 16548 35534
rect 16828 35586 16884 35598
rect 16828 35534 16830 35586
rect 16882 35534 16884 35586
rect 16604 34692 16660 34702
rect 16828 34692 16884 35534
rect 16660 34636 16884 34692
rect 16604 34598 16660 34636
rect 16492 33070 16494 33122
rect 16546 33070 16548 33122
rect 16492 33058 16548 33070
rect 16828 33684 16884 33694
rect 16380 32510 16382 32562
rect 16434 32510 16436 32562
rect 16380 32498 16436 32510
rect 16492 32340 16548 32350
rect 16492 31554 16548 32284
rect 16828 31668 16884 33628
rect 17052 33570 17108 37884
rect 17500 37380 17556 37390
rect 17052 33518 17054 33570
rect 17106 33518 17108 33570
rect 17052 33506 17108 33518
rect 17164 37378 17556 37380
rect 17164 37326 17502 37378
rect 17554 37326 17556 37378
rect 17164 37324 17556 37326
rect 16940 32562 16996 32574
rect 16940 32510 16942 32562
rect 16994 32510 16996 32562
rect 16940 31780 16996 32510
rect 17052 32004 17108 32014
rect 17164 32004 17220 37324
rect 17500 37314 17556 37324
rect 17836 35252 17892 38110
rect 18844 37940 18900 37950
rect 18844 37846 18900 37884
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 17836 35186 17892 35196
rect 18620 37154 18676 37166
rect 18620 37102 18622 37154
rect 18674 37102 18676 37154
rect 17612 35026 17668 35038
rect 17612 34974 17614 35026
rect 17666 34974 17668 35026
rect 17500 34018 17556 34030
rect 17500 33966 17502 34018
rect 17554 33966 17556 34018
rect 17052 32002 17220 32004
rect 17052 31950 17054 32002
rect 17106 31950 17220 32002
rect 17052 31948 17220 31950
rect 17276 33572 17332 33582
rect 17052 31938 17108 31948
rect 17164 31780 17220 31790
rect 16940 31778 17220 31780
rect 16940 31726 17166 31778
rect 17218 31726 17220 31778
rect 16940 31724 17220 31726
rect 16828 31612 16996 31668
rect 16492 31502 16494 31554
rect 16546 31502 16548 31554
rect 16492 31490 16548 31502
rect 16156 30882 16212 30894
rect 16492 30884 16548 30894
rect 16156 30830 16158 30882
rect 16210 30830 16212 30882
rect 16156 30100 16212 30830
rect 16156 30034 16212 30044
rect 16380 30882 16548 30884
rect 16380 30830 16494 30882
rect 16546 30830 16548 30882
rect 16380 30828 16548 30830
rect 16380 30098 16436 30828
rect 16492 30818 16548 30828
rect 16828 30882 16884 30894
rect 16828 30830 16830 30882
rect 16882 30830 16884 30882
rect 16380 30046 16382 30098
rect 16434 30046 16436 30098
rect 16380 30034 16436 30046
rect 16828 30100 16884 30830
rect 16828 30034 16884 30044
rect 15932 29922 15988 29932
rect 15820 28590 15822 28642
rect 15874 28590 15876 28642
rect 15820 28578 15876 28590
rect 16268 29764 16324 29774
rect 16268 27298 16324 29708
rect 16380 29652 16436 29662
rect 16380 29558 16436 29596
rect 16940 29650 16996 31612
rect 16940 29598 16942 29650
rect 16994 29598 16996 29650
rect 16940 29586 16996 29598
rect 17164 30212 17220 31724
rect 17276 31218 17332 33516
rect 17500 33348 17556 33966
rect 17388 33234 17444 33246
rect 17388 33182 17390 33234
rect 17442 33182 17444 33234
rect 17388 32340 17444 33182
rect 17500 32786 17556 33292
rect 17500 32734 17502 32786
rect 17554 32734 17556 32786
rect 17500 32722 17556 32734
rect 17388 32274 17444 32284
rect 17612 31780 17668 34974
rect 18508 34802 18564 34814
rect 18508 34750 18510 34802
rect 18562 34750 18564 34802
rect 17948 34692 18004 34702
rect 17948 34018 18004 34636
rect 17948 33966 17950 34018
rect 18002 33966 18004 34018
rect 17612 31714 17668 31724
rect 17724 33236 17780 33246
rect 17948 33236 18004 33966
rect 18396 34020 18452 34030
rect 18396 33926 18452 33964
rect 17724 33234 18004 33236
rect 17724 33182 17726 33234
rect 17778 33182 18004 33234
rect 17724 33180 18004 33182
rect 18396 33234 18452 33246
rect 18396 33182 18398 33234
rect 18450 33182 18452 33234
rect 17276 31166 17278 31218
rect 17330 31166 17332 31218
rect 17276 31154 17332 31166
rect 16940 29428 16996 29438
rect 16268 27246 16270 27298
rect 16322 27246 16324 27298
rect 16268 27234 16324 27246
rect 16380 28082 16436 28094
rect 16380 28030 16382 28082
rect 16434 28030 16436 28082
rect 16380 26908 16436 28030
rect 16940 28082 16996 29372
rect 17164 28644 17220 30156
rect 17388 30660 17444 30670
rect 17388 29538 17444 30604
rect 17388 29486 17390 29538
rect 17442 29486 17444 29538
rect 17388 29474 17444 29486
rect 17612 30100 17668 30110
rect 17724 30100 17780 33180
rect 18172 32674 18228 32686
rect 18172 32622 18174 32674
rect 18226 32622 18228 32674
rect 18060 32116 18116 32126
rect 17836 31892 17892 31902
rect 17836 31778 17892 31836
rect 17836 31726 17838 31778
rect 17890 31726 17892 31778
rect 17836 31714 17892 31726
rect 18060 31218 18116 32060
rect 18060 31166 18062 31218
rect 18114 31166 18116 31218
rect 18060 31154 18116 31166
rect 17668 30044 17780 30100
rect 17164 28578 17220 28588
rect 17612 29426 17668 30044
rect 18172 29764 18228 32622
rect 18396 30772 18452 33182
rect 18396 30706 18452 30716
rect 18508 30436 18564 34750
rect 18172 29698 18228 29708
rect 18284 30380 18564 30436
rect 17612 29374 17614 29426
rect 17666 29374 17668 29426
rect 16940 28030 16942 28082
rect 16994 28030 16996 28082
rect 16940 28018 16996 28030
rect 17500 28084 17556 28094
rect 17612 28084 17668 29374
rect 18284 29428 18340 30380
rect 18620 30210 18676 37102
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 18732 36594 18788 36606
rect 18732 36542 18734 36594
rect 18786 36542 18788 36594
rect 18732 31892 18788 36542
rect 22428 36594 22484 36606
rect 22428 36542 22430 36594
rect 22482 36542 22484 36594
rect 19740 36372 19796 36382
rect 19628 36370 19796 36372
rect 19628 36318 19742 36370
rect 19794 36318 19796 36370
rect 19628 36316 19796 36318
rect 19516 35810 19572 35822
rect 19516 35758 19518 35810
rect 19570 35758 19572 35810
rect 19516 33796 19572 35758
rect 19516 33730 19572 33740
rect 19628 33572 19684 36316
rect 19740 36306 19796 36316
rect 21196 36372 21252 36382
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20636 35588 20692 35598
rect 20188 35586 20692 35588
rect 20188 35534 20638 35586
rect 20690 35534 20692 35586
rect 20188 35532 20692 35534
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19740 34244 19796 34254
rect 19740 34150 19796 34188
rect 19628 33506 19684 33516
rect 19516 33458 19572 33470
rect 19516 33406 19518 33458
rect 19570 33406 19572 33458
rect 19180 32452 19236 32462
rect 18732 31826 18788 31836
rect 18844 32450 19236 32452
rect 18844 32398 19182 32450
rect 19234 32398 19236 32450
rect 18844 32396 19236 32398
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18620 30146 18676 30158
rect 18732 30772 18788 30782
rect 18284 29362 18340 29372
rect 18396 29426 18452 29438
rect 18396 29374 18398 29426
rect 18450 29374 18452 29426
rect 18284 28532 18340 28542
rect 17500 28082 17668 28084
rect 17500 28030 17502 28082
rect 17554 28030 17668 28082
rect 17500 28028 17668 28030
rect 18060 28418 18116 28430
rect 18060 28366 18062 28418
rect 18114 28366 18116 28418
rect 17500 28018 17556 28028
rect 17388 27076 17444 27086
rect 17388 26908 17444 27020
rect 16380 26852 16548 26908
rect 16492 26402 16548 26852
rect 17052 26850 17108 26862
rect 17388 26852 17556 26908
rect 17052 26798 17054 26850
rect 17106 26798 17108 26850
rect 17052 26516 17108 26798
rect 17052 26450 17108 26460
rect 17500 26514 17556 26796
rect 17500 26462 17502 26514
rect 17554 26462 17556 26514
rect 17500 26450 17556 26462
rect 18060 26514 18116 28366
rect 18284 27858 18340 28476
rect 18396 27972 18452 29374
rect 18732 28868 18788 30716
rect 18844 29426 18900 32396
rect 19180 32386 19236 32396
rect 19068 30212 19124 30222
rect 18844 29374 18846 29426
rect 18898 29374 18900 29426
rect 18844 29362 18900 29374
rect 18956 30156 19068 30212
rect 18844 28868 18900 28878
rect 18732 28866 18900 28868
rect 18732 28814 18846 28866
rect 18898 28814 18900 28866
rect 18732 28812 18900 28814
rect 18844 28802 18900 28812
rect 18396 27906 18452 27916
rect 18284 27806 18286 27858
rect 18338 27806 18340 27858
rect 18284 26852 18340 27806
rect 18284 26786 18340 26796
rect 18060 26462 18062 26514
rect 18114 26462 18116 26514
rect 18060 26450 18116 26462
rect 18844 26516 18900 26526
rect 16492 26350 16494 26402
rect 16546 26350 16548 26402
rect 16492 26338 16548 26350
rect 18844 26402 18900 26460
rect 18844 26350 18846 26402
rect 18898 26350 18900 26402
rect 18844 26338 18900 26350
rect 15484 26226 15540 26236
rect 15820 26178 15876 26190
rect 15820 26126 15822 26178
rect 15874 26126 15876 26178
rect 15484 26068 15540 26078
rect 15484 26066 15764 26068
rect 15484 26014 15486 26066
rect 15538 26014 15764 26066
rect 15484 26012 15764 26014
rect 15484 26002 15540 26012
rect 15372 25394 15428 25406
rect 15372 25342 15374 25394
rect 15426 25342 15428 25394
rect 15372 24948 15428 25342
rect 15372 24882 15428 24892
rect 14924 24434 14980 24444
rect 14924 24052 14980 24062
rect 15148 24052 15204 24062
rect 14924 24050 15148 24052
rect 14924 23998 14926 24050
rect 14978 23998 15148 24050
rect 14924 23996 15148 23998
rect 14924 23986 14980 23996
rect 15148 23986 15204 23996
rect 14028 23940 14084 23950
rect 14028 23826 14084 23884
rect 14028 23774 14030 23826
rect 14082 23774 14084 23826
rect 14028 23762 14084 23774
rect 13916 23426 13972 23436
rect 15260 23492 15316 23502
rect 13916 23266 13972 23278
rect 13916 23214 13918 23266
rect 13970 23214 13972 23266
rect 13132 22932 13188 22942
rect 13132 22838 13188 22876
rect 12796 22642 12852 22652
rect 12572 22306 12628 22316
rect 12684 22484 12740 22494
rect 12236 22148 12292 22158
rect 11900 22146 12292 22148
rect 11900 22094 12238 22146
rect 12290 22094 12292 22146
rect 11900 22092 12292 22094
rect 11900 21698 11956 22092
rect 12236 22082 12292 22092
rect 11900 21646 11902 21698
rect 11954 21646 11956 21698
rect 11900 21634 11956 21646
rect 12124 21588 12180 21598
rect 12124 21494 12180 21532
rect 12684 21586 12740 22428
rect 13804 22372 13860 22382
rect 13804 22278 13860 22316
rect 13020 22260 13076 22270
rect 13020 22166 13076 22204
rect 12684 21534 12686 21586
rect 12738 21534 12740 21586
rect 12684 21522 12740 21534
rect 13356 21812 13412 21822
rect 10220 20130 10276 20142
rect 10220 20078 10222 20130
rect 10274 20078 10276 20130
rect 10220 19908 10276 20078
rect 11564 20132 11732 20188
rect 12460 20802 12516 20814
rect 12460 20750 12462 20802
rect 12514 20750 12516 20802
rect 12460 20188 12516 20750
rect 13020 20804 13076 20814
rect 13356 20804 13412 21756
rect 13916 21700 13972 23214
rect 15036 22260 15092 22270
rect 14476 22148 14532 22158
rect 14476 22054 14532 22092
rect 15036 21810 15092 22204
rect 15036 21758 15038 21810
rect 15090 21758 15092 21810
rect 15036 21746 15092 21758
rect 13916 21634 13972 21644
rect 13020 20802 13412 20804
rect 13020 20750 13022 20802
rect 13074 20750 13358 20802
rect 13410 20750 13412 20802
rect 13020 20748 13412 20750
rect 13020 20738 13076 20748
rect 13356 20738 13412 20748
rect 14028 20802 14084 20814
rect 14028 20750 14030 20802
rect 14082 20750 14084 20802
rect 14028 20188 14084 20750
rect 12460 20132 12852 20188
rect 14028 20132 14308 20188
rect 10668 20020 10724 20030
rect 10220 19842 10276 19852
rect 10556 19964 10668 20020
rect 9884 17938 9940 17948
rect 10220 18562 10276 18574
rect 10220 18510 10222 18562
rect 10274 18510 10276 18562
rect 10220 17668 10276 18510
rect 10220 17602 10276 17612
rect 8652 12450 8708 12460
rect 9324 13076 9380 13086
rect 8092 12238 8094 12290
rect 8146 12238 8148 12290
rect 8092 12226 8148 12238
rect 7756 11230 7758 11282
rect 7810 11230 7812 11282
rect 7756 11218 7812 11230
rect 9324 11282 9380 13020
rect 9548 12068 9604 14812
rect 9772 14756 9828 17388
rect 10108 17108 10164 17118
rect 9996 15540 10052 15550
rect 9884 15204 9940 15214
rect 9884 14868 9940 15148
rect 9884 14802 9940 14812
rect 9660 14700 9828 14756
rect 9660 14642 9716 14700
rect 9996 14644 10052 15484
rect 9660 14590 9662 14642
rect 9714 14590 9716 14642
rect 9660 14578 9716 14590
rect 9772 14642 10052 14644
rect 9772 14590 9998 14642
rect 10050 14590 10052 14642
rect 9772 14588 10052 14590
rect 9660 13972 9716 13982
rect 9772 13972 9828 14588
rect 9996 14578 10052 14588
rect 9660 13970 9828 13972
rect 9660 13918 9662 13970
rect 9714 13918 9828 13970
rect 9660 13916 9828 13918
rect 9660 13906 9716 13916
rect 10108 13076 10164 17052
rect 10220 16996 10276 17006
rect 10220 16902 10276 16940
rect 10444 16324 10500 16334
rect 10332 15540 10388 15550
rect 10332 15446 10388 15484
rect 10444 14642 10500 16268
rect 10444 14590 10446 14642
rect 10498 14590 10500 14642
rect 10444 14578 10500 14590
rect 10556 14420 10612 19964
rect 10668 19954 10724 19964
rect 11452 19124 11508 19134
rect 11452 19010 11508 19068
rect 11452 18958 11454 19010
rect 11506 18958 11508 19010
rect 11452 18946 11508 18958
rect 11228 18676 11284 18686
rect 10444 14364 10612 14420
rect 10668 16884 10724 16894
rect 10220 13076 10276 13086
rect 10108 13074 10276 13076
rect 10108 13022 10222 13074
rect 10274 13022 10276 13074
rect 10108 13020 10276 13022
rect 10220 13010 10276 13020
rect 9660 12068 9716 12078
rect 9548 12012 9660 12068
rect 9660 12002 9716 12012
rect 10444 11506 10500 14364
rect 10444 11454 10446 11506
rect 10498 11454 10500 11506
rect 10444 11442 10500 11454
rect 10556 12516 10612 12526
rect 9324 11230 9326 11282
rect 9378 11230 9380 11282
rect 9324 11218 9380 11230
rect 6748 10670 6750 10722
rect 6802 10670 6804 10722
rect 6748 10658 6804 10670
rect 5964 10446 5966 10498
rect 6018 10446 6020 10498
rect 5964 10434 6020 10446
rect 10556 10498 10612 12460
rect 10556 10446 10558 10498
rect 10610 10446 10612 10498
rect 10556 10434 10612 10446
rect 5852 9886 5854 9938
rect 5906 9886 5908 9938
rect 5852 9874 5908 9886
rect 10556 9940 10612 9950
rect 10668 9940 10724 16828
rect 10780 15204 10836 15214
rect 10780 15110 10836 15148
rect 11228 12850 11284 18620
rect 11452 17556 11508 17566
rect 11452 15874 11508 17500
rect 11452 15822 11454 15874
rect 11506 15822 11508 15874
rect 11452 15810 11508 15822
rect 11564 14420 11620 20132
rect 12460 20020 12516 20030
rect 12460 19926 12516 19964
rect 12236 19124 12292 19134
rect 12236 19030 12292 19068
rect 12572 19124 12628 19134
rect 12572 19030 12628 19068
rect 12012 19010 12068 19022
rect 12012 18958 12014 19010
rect 12066 18958 12068 19010
rect 12012 17220 12068 18958
rect 12124 18564 12180 18574
rect 12124 17442 12180 18508
rect 12124 17390 12126 17442
rect 12178 17390 12180 17442
rect 12124 17378 12180 17390
rect 12572 18450 12628 18462
rect 12572 18398 12574 18450
rect 12626 18398 12628 18450
rect 11900 17164 12068 17220
rect 11900 15426 11956 17164
rect 12460 16884 12516 16894
rect 12460 16790 12516 16828
rect 11900 15374 11902 15426
rect 11954 15374 11956 15426
rect 11900 15362 11956 15374
rect 12012 15874 12068 15886
rect 12012 15822 12014 15874
rect 12066 15822 12068 15874
rect 11676 14420 11732 14430
rect 11564 14418 11732 14420
rect 11564 14366 11678 14418
rect 11730 14366 11732 14418
rect 11564 14364 11732 14366
rect 11676 14354 11732 14364
rect 11228 12798 11230 12850
rect 11282 12798 11284 12850
rect 11228 12786 11284 12798
rect 11788 13412 11844 13422
rect 11788 10722 11844 13356
rect 12012 12292 12068 15822
rect 12348 15876 12404 15886
rect 12348 15204 12404 15820
rect 12348 15138 12404 15148
rect 12572 13634 12628 18398
rect 12684 17442 12740 17454
rect 12684 17390 12686 17442
rect 12738 17390 12740 17442
rect 12684 15652 12740 17390
rect 12684 15586 12740 15596
rect 12796 15202 12852 20132
rect 13020 20020 13076 20030
rect 13244 20020 13300 20030
rect 13020 20018 13300 20020
rect 13020 19966 13022 20018
rect 13074 19966 13246 20018
rect 13298 19966 13300 20018
rect 13020 19964 13300 19966
rect 13020 18452 13076 19964
rect 13244 19954 13300 19964
rect 13916 20018 13972 20030
rect 13916 19966 13918 20018
rect 13970 19966 13972 20018
rect 13692 19234 13748 19246
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13468 19122 13524 19134
rect 13468 19070 13470 19122
rect 13522 19070 13524 19122
rect 13468 18564 13524 19070
rect 13468 18498 13524 18508
rect 13692 19124 13748 19182
rect 13244 18452 13300 18462
rect 13020 18450 13300 18452
rect 13020 18398 13022 18450
rect 13074 18398 13246 18450
rect 13298 18398 13300 18450
rect 13020 18396 13300 18398
rect 13020 17444 13076 18396
rect 13244 18386 13300 18396
rect 13020 16884 13076 17388
rect 13468 17668 13524 17678
rect 13468 16994 13524 17612
rect 13692 17668 13748 19068
rect 13916 18676 13972 19966
rect 14140 19124 14196 19134
rect 14140 19030 14196 19068
rect 13916 18620 14196 18676
rect 13916 18452 13972 18462
rect 13916 18450 14084 18452
rect 13916 18398 13918 18450
rect 13970 18398 14084 18450
rect 13916 18396 14084 18398
rect 13916 18386 13972 18396
rect 13804 17668 13860 17678
rect 13692 17666 13860 17668
rect 13692 17614 13806 17666
rect 13858 17614 13860 17666
rect 13692 17612 13860 17614
rect 13580 17556 13636 17566
rect 13580 17462 13636 17500
rect 13468 16942 13470 16994
rect 13522 16942 13524 16994
rect 13468 16930 13524 16942
rect 13020 16882 13412 16884
rect 13020 16830 13022 16882
rect 13074 16830 13412 16882
rect 13020 16828 13412 16830
rect 12908 15876 12964 15886
rect 12908 15782 12964 15820
rect 13020 15540 13076 16828
rect 13356 16660 13412 16828
rect 13692 16882 13748 17612
rect 13804 17602 13860 17612
rect 13692 16830 13694 16882
rect 13746 16830 13748 16882
rect 13692 16772 13748 16830
rect 13356 16604 13636 16660
rect 13580 16210 13636 16604
rect 13580 16158 13582 16210
rect 13634 16158 13636 16210
rect 13580 16146 13636 16158
rect 13692 15876 13748 16716
rect 14028 16212 14084 18396
rect 14140 16884 14196 18620
rect 14140 16818 14196 16828
rect 14028 16146 14084 16156
rect 13692 15810 13748 15820
rect 14028 15876 14084 15886
rect 14028 15782 14084 15820
rect 13020 15474 13076 15484
rect 13580 15652 13636 15662
rect 12796 15150 12798 15202
rect 12850 15150 12852 15202
rect 12796 15138 12852 15150
rect 13580 13858 13636 15596
rect 13580 13806 13582 13858
rect 13634 13806 13636 13858
rect 13580 13794 13636 13806
rect 12572 13582 12574 13634
rect 12626 13582 12628 13634
rect 12572 13570 12628 13582
rect 14252 13076 14308 20132
rect 14812 19460 14868 19470
rect 14700 19404 14812 19460
rect 14364 19236 14420 19246
rect 14364 19142 14420 19180
rect 14364 17444 14420 17454
rect 14364 17350 14420 17388
rect 14700 16994 14756 19404
rect 14812 19394 14868 19404
rect 14924 19236 14980 19246
rect 14924 19142 14980 19180
rect 15148 19010 15204 19022
rect 15148 18958 15150 19010
rect 15202 18958 15204 19010
rect 14924 17668 14980 17678
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 14812 17442 14868 17454
rect 14812 17390 14814 17442
rect 14866 17390 14868 17442
rect 14812 16772 14868 17390
rect 14812 16706 14868 16716
rect 14588 16100 14644 16110
rect 14588 15202 14644 16044
rect 14924 16098 14980 17612
rect 15148 17108 15204 18958
rect 15260 17778 15316 23436
rect 15708 23380 15764 26012
rect 15820 25508 15876 26126
rect 15820 25442 15876 25452
rect 16044 26178 16100 26190
rect 16044 26126 16046 26178
rect 16098 26126 16100 26178
rect 16044 24948 16100 26126
rect 16828 26180 16884 26190
rect 16828 26086 16884 26124
rect 17948 26180 18004 26190
rect 17948 26086 18004 26124
rect 18620 26180 18676 26190
rect 16380 25618 16436 25630
rect 16380 25566 16382 25618
rect 16434 25566 16436 25618
rect 16156 24948 16212 24958
rect 16044 24946 16212 24948
rect 16044 24894 16158 24946
rect 16210 24894 16212 24946
rect 16044 24892 16212 24894
rect 16156 24882 16212 24892
rect 16380 24388 16436 25566
rect 17500 24724 17556 24734
rect 17500 24630 17556 24668
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 16940 24500 16996 24510
rect 17500 24500 17556 24510
rect 16940 24498 17332 24500
rect 16940 24446 16942 24498
rect 16994 24446 17332 24498
rect 16940 24444 17332 24446
rect 16940 24434 16996 24444
rect 16380 24322 16436 24332
rect 16268 23716 16324 23726
rect 16268 23622 16324 23660
rect 17052 23716 17108 23726
rect 17052 23622 17108 23660
rect 15708 23324 16548 23380
rect 16156 23156 16212 23166
rect 15932 23154 16212 23156
rect 15932 23102 16158 23154
rect 16210 23102 16212 23154
rect 15932 23100 16212 23102
rect 15820 21362 15876 21374
rect 15820 21310 15822 21362
rect 15874 21310 15876 21362
rect 15820 19460 15876 21310
rect 15820 19394 15876 19404
rect 15932 19236 15988 23100
rect 16156 23090 16212 23100
rect 16380 22260 16436 22270
rect 16380 22166 16436 22204
rect 16380 21700 16436 21710
rect 16380 21606 16436 21644
rect 16380 20578 16436 20590
rect 16380 20526 16382 20578
rect 16434 20526 16436 20578
rect 16156 20132 16212 20142
rect 16156 20130 16324 20132
rect 16156 20078 16158 20130
rect 16210 20078 16324 20130
rect 16156 20076 16324 20078
rect 16156 20066 16212 20076
rect 15820 19180 15988 19236
rect 15260 17726 15262 17778
rect 15314 17726 15316 17778
rect 15260 17714 15316 17726
rect 15708 18340 15764 18350
rect 15148 17052 15652 17108
rect 15148 16884 15204 16894
rect 14924 16046 14926 16098
rect 14978 16046 14980 16098
rect 14924 16034 14980 16046
rect 15036 16324 15092 16334
rect 14588 15150 14590 15202
rect 14642 15150 14644 15202
rect 14588 15138 14644 15150
rect 15036 14418 15092 16268
rect 15148 15148 15204 16828
rect 15484 16212 15540 16222
rect 15260 16100 15316 16110
rect 15260 16006 15316 16044
rect 15148 15092 15428 15148
rect 15036 14366 15038 14418
rect 15090 14366 15092 14418
rect 15036 14354 15092 14366
rect 15372 13634 15428 15092
rect 15372 13582 15374 13634
rect 15426 13582 15428 13634
rect 15372 13570 15428 13582
rect 14364 13076 14420 13086
rect 14252 13020 14364 13076
rect 14364 13010 14420 13020
rect 15484 13074 15540 16156
rect 15596 13860 15652 17052
rect 15708 15426 15764 18284
rect 15820 16770 15876 19180
rect 15932 19012 15988 19022
rect 15932 18918 15988 18956
rect 16268 18452 16324 20076
rect 16380 19348 16436 20526
rect 16380 19282 16436 19292
rect 16268 18386 16324 18396
rect 16380 18674 16436 18686
rect 16380 18622 16382 18674
rect 16434 18622 16436 18674
rect 16380 17108 16436 18622
rect 16492 17554 16548 23324
rect 16828 23154 16884 23166
rect 16828 23102 16830 23154
rect 16882 23102 16884 23154
rect 16716 23044 16772 23054
rect 16716 22482 16772 22988
rect 16716 22430 16718 22482
rect 16770 22430 16772 22482
rect 16716 22148 16772 22430
rect 16828 22372 16884 23102
rect 17164 22372 17220 22382
rect 16828 22370 17220 22372
rect 16828 22318 17166 22370
rect 17218 22318 17220 22370
rect 16828 22316 17220 22318
rect 16716 21698 16772 22092
rect 17164 21924 17220 22316
rect 17164 21858 17220 21868
rect 16716 21646 16718 21698
rect 16770 21646 16772 21698
rect 16716 21634 16772 21646
rect 17052 20578 17108 20590
rect 17052 20526 17054 20578
rect 17106 20526 17108 20578
rect 16940 19796 16996 19806
rect 16828 19794 16996 19796
rect 16828 19742 16942 19794
rect 16994 19742 16996 19794
rect 16828 19740 16996 19742
rect 16716 18340 16772 18350
rect 16828 18340 16884 19740
rect 16940 19730 16996 19740
rect 16772 18284 16884 18340
rect 16716 18274 16772 18284
rect 16940 18228 16996 18238
rect 16492 17502 16494 17554
rect 16546 17502 16548 17554
rect 16492 17490 16548 17502
rect 16828 18226 16996 18228
rect 16828 18174 16942 18226
rect 16994 18174 16996 18226
rect 16828 18172 16996 18174
rect 16380 17042 16436 17052
rect 15820 16718 15822 16770
rect 15874 16718 15876 16770
rect 15820 16706 15876 16718
rect 15708 15374 15710 15426
rect 15762 15374 15764 15426
rect 15708 15362 15764 15374
rect 16268 16436 16324 16446
rect 16268 14642 16324 16380
rect 16828 16324 16884 18172
rect 16940 18162 16996 18172
rect 16940 17668 16996 17678
rect 16940 17574 16996 17612
rect 16828 16258 16884 16268
rect 17052 15148 17108 20526
rect 17164 20578 17220 20590
rect 17164 20526 17166 20578
rect 17218 20526 17220 20578
rect 17164 15540 17220 20526
rect 17164 15474 17220 15484
rect 17276 15428 17332 24444
rect 17500 23378 17556 24444
rect 17836 24276 17892 24670
rect 17836 24210 17892 24220
rect 17500 23326 17502 23378
rect 17554 23326 17556 23378
rect 17500 23314 17556 23326
rect 17388 23044 17444 23054
rect 17388 22950 17444 22988
rect 18060 23044 18116 23054
rect 17836 22370 17892 22382
rect 17836 22318 17838 22370
rect 17890 22318 17892 22370
rect 17724 22036 17780 22046
rect 17724 20020 17780 21980
rect 17836 20356 17892 22318
rect 17948 21586 18004 21598
rect 17948 21534 17950 21586
rect 18002 21534 18004 21586
rect 17948 20804 18004 21534
rect 17948 20738 18004 20748
rect 17948 20580 18004 20590
rect 18060 20580 18116 22988
rect 18172 23042 18228 23054
rect 18172 22990 18174 23042
rect 18226 22990 18228 23042
rect 18172 22036 18228 22990
rect 18172 21970 18228 21980
rect 18508 21924 18564 21934
rect 18508 21474 18564 21868
rect 18508 21422 18510 21474
rect 18562 21422 18564 21474
rect 18508 21410 18564 21422
rect 17948 20578 18116 20580
rect 17948 20526 17950 20578
rect 18002 20526 18116 20578
rect 17948 20524 18116 20526
rect 17948 20514 18004 20524
rect 17836 20300 18564 20356
rect 17836 20020 17892 20030
rect 17724 19964 17836 20020
rect 17836 19926 17892 19964
rect 18284 19234 18340 19246
rect 18284 19182 18286 19234
rect 18338 19182 18340 19234
rect 17836 18452 17892 18462
rect 18172 18452 18228 18462
rect 17836 18358 17892 18396
rect 18060 18396 18172 18452
rect 17500 17666 17556 17678
rect 17500 17614 17502 17666
rect 17554 17614 17556 17666
rect 17500 16436 17556 17614
rect 17724 17108 17780 17118
rect 17724 16994 17780 17052
rect 17724 16942 17726 16994
rect 17778 16942 17780 16994
rect 17724 16930 17780 16942
rect 18060 16996 18116 18396
rect 18172 18358 18228 18396
rect 18284 17220 18340 19182
rect 18508 17220 18564 20300
rect 18620 19906 18676 26124
rect 18956 25618 19012 30156
rect 19068 30118 19124 30156
rect 19068 29652 19124 29662
rect 19068 28754 19124 29596
rect 19068 28702 19070 28754
rect 19122 28702 19124 28754
rect 19068 28690 19124 28702
rect 19292 28644 19348 28654
rect 19180 28642 19348 28644
rect 19180 28590 19294 28642
rect 19346 28590 19348 28642
rect 19180 28588 19348 28590
rect 19068 27972 19124 27982
rect 19068 27746 19124 27916
rect 19068 27694 19070 27746
rect 19122 27694 19124 27746
rect 19068 27682 19124 27694
rect 19180 26908 19236 28588
rect 19292 28578 19348 28588
rect 19404 27076 19460 27086
rect 19516 27076 19572 33406
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 30996 20244 35532
rect 20636 35522 20692 35532
rect 20636 35028 20692 35038
rect 20524 34972 20636 35028
rect 20300 31556 20356 31566
rect 20300 31554 20468 31556
rect 20300 31502 20302 31554
rect 20354 31502 20468 31554
rect 20300 31500 20468 31502
rect 20300 31490 20356 31500
rect 20300 30996 20356 31006
rect 20188 30994 20356 30996
rect 20188 30942 20302 30994
rect 20354 30942 20356 30994
rect 20188 30940 20356 30942
rect 20300 30930 20356 30940
rect 20412 30210 20468 31500
rect 20412 30158 20414 30210
rect 20466 30158 20468 30210
rect 20412 30146 20468 30158
rect 20524 29988 20580 34972
rect 20636 34962 20692 34972
rect 20636 32562 20692 32574
rect 20636 32510 20638 32562
rect 20690 32510 20692 32562
rect 20636 30996 20692 32510
rect 20860 32004 20916 32014
rect 20860 31890 20916 31948
rect 20860 31838 20862 31890
rect 20914 31838 20916 31890
rect 20860 31826 20916 31838
rect 21196 31890 21252 36316
rect 22316 35028 22372 35038
rect 22316 34934 22372 34972
rect 21308 34580 21364 34590
rect 21308 32562 21364 34524
rect 22428 34580 22484 36542
rect 23548 36372 23604 36382
rect 23548 36278 23604 36316
rect 22652 35812 22708 35822
rect 22652 35810 22820 35812
rect 22652 35758 22654 35810
rect 22706 35758 22820 35810
rect 22652 35756 22820 35758
rect 22652 35746 22708 35756
rect 22428 34514 22484 34524
rect 21532 34244 21588 34254
rect 21308 32510 21310 32562
rect 21362 32510 21364 32562
rect 21308 32498 21364 32510
rect 21420 34242 21588 34244
rect 21420 34190 21534 34242
rect 21586 34190 21588 34242
rect 21420 34188 21588 34190
rect 21196 31838 21198 31890
rect 21250 31838 21252 31890
rect 21196 31826 21252 31838
rect 20748 30996 20804 31006
rect 21084 30996 21140 31006
rect 20636 30994 21140 30996
rect 20636 30942 20750 30994
rect 20802 30942 21086 30994
rect 21138 30942 21140 30994
rect 20636 30940 21140 30942
rect 20636 30212 20692 30940
rect 20748 30930 20804 30940
rect 21084 30930 21140 30940
rect 21420 30324 21476 34188
rect 21532 34178 21588 34188
rect 22652 34020 22708 34030
rect 21868 34018 22708 34020
rect 21868 33966 22654 34018
rect 22706 33966 22708 34018
rect 21868 33964 22708 33966
rect 21644 33234 21700 33246
rect 21644 33182 21646 33234
rect 21698 33182 21700 33234
rect 21532 33122 21588 33134
rect 21532 33070 21534 33122
rect 21586 33070 21588 33122
rect 21532 32116 21588 33070
rect 21532 32050 21588 32060
rect 21644 33124 21700 33182
rect 20636 30146 20692 30156
rect 21308 30268 21476 30324
rect 20748 30100 20804 30110
rect 20748 30006 20804 30044
rect 20188 29932 20580 29988
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19404 27074 19572 27076
rect 19404 27022 19406 27074
rect 19458 27022 19572 27074
rect 19404 27020 19572 27022
rect 19740 27972 19796 27982
rect 19740 27074 19796 27916
rect 19740 27022 19742 27074
rect 19794 27022 19796 27074
rect 19404 27010 19460 27020
rect 19740 26964 19796 27022
rect 19068 26852 19236 26908
rect 19628 26852 19796 26908
rect 19068 26290 19124 26852
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 26180 19124 26238
rect 19628 26290 19684 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26226 19684 26238
rect 20188 26290 20244 29932
rect 21196 29540 21252 29550
rect 20300 29538 21252 29540
rect 20300 29486 21198 29538
rect 21250 29486 21252 29538
rect 20300 29484 21252 29486
rect 20300 27186 20356 29484
rect 21196 29474 21252 29484
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 20300 27122 20356 27134
rect 20524 28868 20580 28878
rect 20524 27186 20580 28812
rect 20748 28644 20804 28654
rect 20524 27134 20526 27186
rect 20578 27134 20580 27186
rect 20524 27122 20580 27134
rect 20636 28588 20748 28644
rect 20188 26238 20190 26290
rect 20242 26238 20244 26290
rect 20188 26226 20244 26238
rect 19068 26114 19124 26124
rect 18956 25566 18958 25618
rect 19010 25566 19012 25618
rect 18956 25554 19012 25566
rect 20300 25506 20356 25518
rect 20300 25454 20302 25506
rect 20354 25454 20356 25506
rect 20300 25284 20356 25454
rect 20636 25284 20692 28588
rect 20748 28550 20804 28588
rect 21308 28420 21364 30268
rect 21532 30212 21588 30222
rect 21644 30212 21700 33068
rect 21756 33012 21812 33022
rect 21756 30994 21812 32956
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 21756 30930 21812 30942
rect 21532 30210 21700 30212
rect 21532 30158 21534 30210
rect 21586 30158 21700 30210
rect 21532 30156 21700 30158
rect 21532 30146 21588 30156
rect 21644 30100 21700 30156
rect 21644 28868 21700 30044
rect 20748 28364 21364 28420
rect 21532 28756 21588 28766
rect 20748 28082 20804 28364
rect 20748 28030 20750 28082
rect 20802 28030 20804 28082
rect 20748 28018 20804 28030
rect 21532 28082 21588 28700
rect 21644 28754 21700 28812
rect 21644 28702 21646 28754
rect 21698 28702 21700 28754
rect 21644 28690 21700 28702
rect 21756 30098 21812 30110
rect 21756 30046 21758 30098
rect 21810 30046 21812 30098
rect 21532 28030 21534 28082
rect 21586 28030 21588 28082
rect 21532 28018 21588 28030
rect 21196 27074 21252 27086
rect 21196 27022 21198 27074
rect 21250 27022 21252 27074
rect 21196 26964 21252 27022
rect 20748 25284 20804 25294
rect 20636 25228 20748 25284
rect 20300 25218 20356 25228
rect 20748 25190 20804 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20412 24946 20468 24958
rect 20412 24894 20414 24946
rect 20466 24894 20468 24946
rect 19964 24724 20020 24734
rect 19292 23940 19348 23950
rect 18620 19854 18622 19906
rect 18674 19854 18676 19906
rect 18620 18562 18676 19854
rect 18620 18510 18622 18562
rect 18674 18510 18676 18562
rect 18620 18452 18676 18510
rect 18620 18386 18676 18396
rect 18732 23938 19348 23940
rect 18732 23886 19294 23938
rect 19346 23886 19348 23938
rect 18732 23884 19348 23886
rect 18508 17164 18676 17220
rect 18284 17154 18340 17164
rect 18060 16902 18116 16940
rect 18620 16772 18676 17164
rect 17500 16370 17556 16380
rect 18508 16716 18676 16772
rect 17836 15988 17892 15998
rect 17836 15874 17892 15932
rect 17836 15822 17838 15874
rect 17890 15822 17892 15874
rect 17836 15810 17892 15822
rect 18396 15874 18452 15886
rect 18396 15822 18398 15874
rect 18450 15822 18452 15874
rect 17500 15428 17556 15438
rect 17276 15426 17556 15428
rect 17276 15374 17502 15426
rect 17554 15374 17556 15426
rect 17276 15372 17556 15374
rect 17500 15362 17556 15372
rect 17052 15092 18004 15148
rect 16268 14590 16270 14642
rect 16322 14590 16324 14642
rect 16268 14578 16324 14590
rect 16828 13972 16884 13982
rect 16716 13916 16828 13972
rect 16380 13860 16436 13870
rect 15596 13858 16436 13860
rect 15596 13806 16382 13858
rect 16434 13806 16436 13858
rect 15596 13804 16436 13806
rect 16380 13794 16436 13804
rect 15484 13022 15486 13074
rect 15538 13022 15540 13074
rect 15484 13010 15540 13022
rect 16716 12850 16772 13916
rect 16828 13906 16884 13916
rect 16716 12798 16718 12850
rect 16770 12798 16772 12850
rect 16716 12786 16772 12798
rect 13020 12292 13076 12302
rect 12012 12290 13076 12292
rect 12012 12238 13022 12290
rect 13074 12238 13076 12290
rect 12012 12236 13076 12238
rect 13020 12226 13076 12236
rect 17948 12290 18004 15092
rect 18396 13972 18452 15822
rect 18508 15148 18564 16716
rect 18620 15988 18676 15998
rect 18620 15894 18676 15932
rect 18732 15202 18788 23884
rect 19292 23874 19348 23884
rect 19964 23938 20020 24668
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 19964 23874 20020 23886
rect 20188 24388 20244 24398
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19404 23268 19460 23278
rect 19404 23174 19460 23212
rect 19628 23154 19684 23166
rect 19628 23102 19630 23154
rect 19682 23102 19684 23154
rect 19068 23044 19124 23054
rect 19068 22950 19124 22988
rect 19404 22260 19460 22270
rect 19292 22204 19404 22260
rect 19180 19346 19236 19358
rect 19180 19294 19182 19346
rect 19234 19294 19236 19346
rect 18844 19236 18900 19246
rect 18844 19234 19124 19236
rect 18844 19182 18846 19234
rect 18898 19182 19124 19234
rect 18844 19180 19124 19182
rect 18844 19170 18900 19180
rect 18844 18676 18900 18686
rect 18844 16994 18900 18620
rect 19068 18452 19124 19180
rect 19180 19012 19236 19294
rect 19180 18946 19236 18956
rect 19292 18900 19348 22204
rect 19404 22194 19460 22204
rect 19628 21924 19684 23102
rect 20188 23154 20244 24332
rect 20412 24050 20468 24894
rect 20972 24948 21028 24958
rect 20972 24854 21028 24892
rect 21196 24724 21252 26908
rect 21756 26908 21812 30046
rect 21868 27074 21924 33964
rect 22652 33954 22708 33964
rect 22764 32004 22820 35756
rect 23660 35588 23716 35598
rect 23660 35586 24276 35588
rect 23660 35534 23662 35586
rect 23714 35534 24276 35586
rect 23660 35532 24276 35534
rect 23660 35522 23716 35532
rect 23548 34802 23604 34814
rect 23548 34750 23550 34802
rect 23602 34750 23604 34802
rect 22764 31938 22820 31948
rect 22988 33234 23044 33246
rect 22988 33182 22990 33234
rect 23042 33182 23044 33234
rect 21980 31668 22036 31678
rect 22988 31668 23044 33182
rect 21980 31666 23044 31668
rect 21980 31614 21982 31666
rect 22034 31614 23044 31666
rect 21980 31612 23044 31614
rect 23212 33236 23268 33246
rect 21980 31602 22036 31612
rect 22204 31444 22260 31454
rect 22092 31388 22204 31444
rect 21980 29988 22036 29998
rect 21980 29894 22036 29932
rect 21980 29652 22036 29662
rect 22092 29652 22148 31388
rect 22204 31378 22260 31388
rect 22764 29988 22820 29998
rect 22764 29894 22820 29932
rect 21980 29650 22148 29652
rect 21980 29598 21982 29650
rect 22034 29598 22148 29650
rect 21980 29596 22148 29598
rect 21980 29586 22036 29596
rect 22652 29538 22708 29550
rect 22652 29486 22654 29538
rect 22706 29486 22708 29538
rect 22652 27300 22708 29486
rect 22652 27234 22708 27244
rect 21868 27022 21870 27074
rect 21922 27022 21924 27074
rect 21868 27010 21924 27022
rect 21756 26852 22484 26908
rect 22428 26514 22484 26852
rect 22428 26462 22430 26514
rect 22482 26462 22484 26514
rect 22428 26450 22484 26462
rect 23212 26514 23268 33180
rect 23324 33234 23380 33246
rect 23324 33182 23326 33234
rect 23378 33182 23380 33234
rect 23324 33124 23380 33182
rect 23324 33058 23380 33068
rect 23548 32900 23604 34750
rect 23436 32844 23604 32900
rect 23436 32452 23492 32844
rect 23772 32786 23828 32798
rect 23772 32734 23774 32786
rect 23826 32734 23828 32786
rect 23436 32396 23604 32452
rect 23548 31444 23604 32396
rect 23548 31378 23604 31388
rect 23772 30884 23828 32734
rect 24220 31778 24276 35532
rect 34636 35476 34692 35486
rect 25116 35026 25172 35038
rect 32620 35028 32676 35038
rect 25116 34974 25118 35026
rect 25170 34974 25172 35026
rect 24332 34804 24388 34814
rect 24332 32786 24388 34748
rect 24668 33460 24724 33470
rect 24332 32734 24334 32786
rect 24386 32734 24388 32786
rect 24332 32722 24388 32734
rect 24444 33458 24724 33460
rect 24444 33406 24670 33458
rect 24722 33406 24724 33458
rect 24444 33404 24724 33406
rect 24220 31726 24222 31778
rect 24274 31726 24276 31778
rect 24220 31714 24276 31726
rect 24220 31218 24276 31230
rect 24220 31166 24222 31218
rect 24274 31166 24276 31218
rect 24220 31108 24276 31166
rect 24220 31042 24276 31052
rect 23772 30818 23828 30828
rect 24444 30660 24500 33404
rect 24668 33394 24724 33404
rect 24892 33124 24948 33134
rect 24780 31780 24836 31790
rect 24780 31686 24836 31724
rect 24780 31220 24836 31230
rect 24892 31220 24948 33068
rect 25116 33012 25172 34974
rect 32060 35026 32676 35028
rect 32060 34974 32622 35026
rect 32674 34974 32676 35026
rect 32060 34972 32676 34974
rect 26124 34804 26180 34814
rect 31500 34804 31556 34814
rect 26124 34710 26180 34748
rect 30380 34802 31556 34804
rect 30380 34750 31502 34802
rect 31554 34750 31556 34802
rect 30380 34748 31556 34750
rect 27244 34242 27300 34254
rect 27244 34190 27246 34242
rect 27298 34190 27300 34242
rect 26236 34018 26292 34030
rect 26236 33966 26238 34018
rect 26290 33966 26292 34018
rect 25788 33348 25844 33358
rect 25676 33236 25732 33246
rect 25676 33142 25732 33180
rect 25116 32946 25172 32956
rect 24780 31218 24948 31220
rect 24780 31166 24782 31218
rect 24834 31166 24948 31218
rect 24780 31164 24948 31166
rect 25116 31892 25172 31902
rect 24780 31154 24836 31164
rect 23884 30604 24500 30660
rect 23660 29314 23716 29326
rect 23660 29262 23662 29314
rect 23714 29262 23716 29314
rect 23660 27860 23716 29262
rect 23772 28642 23828 28654
rect 23772 28590 23774 28642
rect 23826 28590 23828 28642
rect 23772 28532 23828 28590
rect 23772 28466 23828 28476
rect 23660 27794 23716 27804
rect 23884 27858 23940 30604
rect 25116 30210 25172 31836
rect 25228 31780 25284 31790
rect 25228 31686 25284 31724
rect 25676 31780 25732 31790
rect 25788 31780 25844 33292
rect 26236 31892 26292 33966
rect 27244 33124 27300 34190
rect 28924 34244 28980 34254
rect 27244 33058 27300 33068
rect 28252 33234 28308 33246
rect 28252 33182 28254 33234
rect 28306 33182 28308 33234
rect 26236 31826 26292 31836
rect 26572 32562 26628 32574
rect 26572 32510 26574 32562
rect 26626 32510 26628 32562
rect 25676 31778 25844 31780
rect 25676 31726 25678 31778
rect 25730 31726 25844 31778
rect 25676 31724 25844 31726
rect 26012 31780 26068 31790
rect 25676 31714 25732 31724
rect 25228 31108 25284 31118
rect 25228 31014 25284 31052
rect 26012 30994 26068 31724
rect 26572 31780 26628 32510
rect 26572 31714 26628 31724
rect 27244 32562 27300 32574
rect 27244 32510 27246 32562
rect 27298 32510 27300 32562
rect 26012 30942 26014 30994
rect 26066 30942 26068 30994
rect 25116 30158 25118 30210
rect 25170 30158 25172 30210
rect 25116 30146 25172 30158
rect 25228 30884 25284 30894
rect 24892 30100 24948 30110
rect 24444 28868 24500 28878
rect 24220 28756 24276 28766
rect 24220 28662 24276 28700
rect 24444 28642 24500 28812
rect 24444 28590 24446 28642
rect 24498 28590 24500 28642
rect 24444 28578 24500 28590
rect 23884 27806 23886 27858
rect 23938 27806 23940 27858
rect 23884 27794 23940 27806
rect 24444 27858 24500 27870
rect 24444 27806 24446 27858
rect 24498 27806 24500 27858
rect 24108 27748 24164 27758
rect 24108 26962 24164 27692
rect 24444 27188 24500 27806
rect 24892 27298 24948 30044
rect 25228 29538 25284 30828
rect 25228 29486 25230 29538
rect 25282 29486 25284 29538
rect 25228 29474 25284 29486
rect 25564 30882 25620 30894
rect 25564 30830 25566 30882
rect 25618 30830 25620 30882
rect 25452 29428 25508 29438
rect 25564 29428 25620 30830
rect 25676 30212 25732 30222
rect 25676 30118 25732 30156
rect 26012 30212 26068 30942
rect 26684 30996 26740 31006
rect 26684 30902 26740 30940
rect 27244 30884 27300 32510
rect 28252 32564 28308 33182
rect 28700 33236 28756 33246
rect 28140 32452 28196 32462
rect 28140 31554 28196 32396
rect 28140 31502 28142 31554
rect 28194 31502 28196 31554
rect 28140 31490 28196 31502
rect 27244 30818 27300 30828
rect 26908 30324 26964 30334
rect 26012 30146 26068 30156
rect 26796 30322 26964 30324
rect 26796 30270 26910 30322
rect 26962 30270 26964 30322
rect 26796 30268 26964 30270
rect 26012 29988 26068 29998
rect 26012 29650 26068 29932
rect 26012 29598 26014 29650
rect 26066 29598 26068 29650
rect 26012 29586 26068 29598
rect 25900 29428 25956 29438
rect 25452 29426 25956 29428
rect 25452 29374 25454 29426
rect 25506 29374 25902 29426
rect 25954 29374 25956 29426
rect 25452 29372 25956 29374
rect 25452 28868 25508 29372
rect 25900 29362 25956 29372
rect 25004 28642 25060 28654
rect 25004 28590 25006 28642
rect 25058 28590 25060 28642
rect 25004 28532 25060 28590
rect 25004 27636 25060 28476
rect 25452 27858 25508 28812
rect 26572 28644 26628 28654
rect 26572 28550 26628 28588
rect 25452 27806 25454 27858
rect 25506 27806 25508 27858
rect 25452 27794 25508 27806
rect 25228 27748 25284 27758
rect 25228 27654 25284 27692
rect 25004 27570 25060 27580
rect 24892 27246 24894 27298
rect 24946 27246 24948 27298
rect 24892 27234 24948 27246
rect 25004 27300 25060 27310
rect 25004 27206 25060 27244
rect 24444 27122 24500 27132
rect 25116 27188 25172 27198
rect 24108 26910 24110 26962
rect 24162 26910 24164 26962
rect 24108 26898 24164 26910
rect 25004 26964 25060 26974
rect 23212 26462 23214 26514
rect 23266 26462 23268 26514
rect 23212 26450 23268 26462
rect 22204 26292 22260 26302
rect 22092 25394 22148 25406
rect 22092 25342 22094 25394
rect 22146 25342 22148 25394
rect 22092 24948 22148 25342
rect 22092 24882 22148 24892
rect 21196 24630 21252 24668
rect 21644 24722 21700 24734
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 20412 23998 20414 24050
rect 20466 23998 20468 24050
rect 20412 23986 20468 23998
rect 21644 24052 21700 24670
rect 21644 23986 21700 23996
rect 22204 24052 22260 26236
rect 23100 26292 23156 26302
rect 23100 25618 23156 26236
rect 23100 25566 23102 25618
rect 23154 25566 23156 25618
rect 23100 25554 23156 25566
rect 23884 26290 23940 26302
rect 23884 26238 23886 26290
rect 23938 26238 23940 26290
rect 23660 25172 23716 25182
rect 22204 23958 22260 23996
rect 23324 24052 23380 24062
rect 23212 23940 23268 23950
rect 20748 23828 20804 23838
rect 20748 23268 20804 23772
rect 21308 23826 21364 23838
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23716 21364 23774
rect 21308 23650 21364 23660
rect 21644 23828 21700 23838
rect 20748 23202 20804 23212
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 20188 23090 20244 23102
rect 21196 23044 21252 23054
rect 20300 22146 20356 22158
rect 20860 22148 20916 22158
rect 20300 22094 20302 22146
rect 20354 22094 20356 22146
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21858 19684 21868
rect 20188 20802 20244 20814
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19852 19348 19908 19358
rect 19404 19236 19460 19246
rect 19404 19234 19796 19236
rect 19404 19182 19406 19234
rect 19458 19182 19796 19234
rect 19404 19180 19796 19182
rect 19404 19170 19460 19180
rect 19740 19122 19796 19180
rect 19740 19070 19742 19122
rect 19794 19070 19796 19122
rect 19740 19012 19796 19070
rect 19628 18956 19796 19012
rect 19852 19010 19908 19292
rect 19852 18958 19854 19010
rect 19906 18958 19908 19010
rect 19292 18844 19572 18900
rect 19180 18452 19236 18462
rect 19068 18450 19236 18452
rect 19068 18398 19182 18450
rect 19234 18398 19236 18450
rect 19068 18396 19236 18398
rect 18956 18340 19012 18350
rect 18956 18246 19012 18284
rect 19180 17668 19236 18396
rect 19180 17602 19236 17612
rect 19068 17220 19124 17230
rect 18844 16942 18846 16994
rect 18898 16942 18900 16994
rect 18844 16930 18900 16942
rect 18956 16996 19012 17006
rect 18956 16210 19012 16940
rect 18956 16158 18958 16210
rect 19010 16158 19012 16210
rect 18956 16146 19012 16158
rect 18732 15150 18734 15202
rect 18786 15150 18788 15202
rect 18508 15092 18676 15148
rect 18732 15138 18788 15150
rect 18620 14642 18676 15092
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 18396 13906 18452 13916
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 12226 18004 12238
rect 12012 12068 12068 12078
rect 12012 11974 12068 12012
rect 19068 12066 19124 17164
rect 19516 16772 19572 18844
rect 19628 18452 19684 18956
rect 19852 18946 19908 18958
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18386 19684 18396
rect 19740 18450 19796 18462
rect 19740 18398 19742 18450
rect 19794 18398 19796 18450
rect 19740 17444 19796 18398
rect 19852 18340 19908 18350
rect 19852 17554 19908 18284
rect 20188 18004 20244 20750
rect 20300 20580 20356 22094
rect 20748 22146 20916 22148
rect 20748 22094 20862 22146
rect 20914 22094 20916 22146
rect 20748 22092 20916 22094
rect 20412 21364 20468 21374
rect 20412 21362 20580 21364
rect 20412 21310 20414 21362
rect 20466 21310 20580 21362
rect 20412 21308 20580 21310
rect 20412 21298 20468 21308
rect 20300 20514 20356 20524
rect 20412 20804 20468 20814
rect 20412 20130 20468 20748
rect 20412 20078 20414 20130
rect 20466 20078 20468 20130
rect 20412 20066 20468 20078
rect 20300 19572 20356 19582
rect 20300 18676 20356 19516
rect 20524 19348 20580 21308
rect 20748 19572 20804 22092
rect 20860 22082 20916 22092
rect 21196 21810 21252 22988
rect 21420 22372 21476 22382
rect 21420 22278 21476 22316
rect 21196 21758 21198 21810
rect 21250 21758 21252 21810
rect 21196 21746 21252 21758
rect 21532 20916 21588 20926
rect 20860 20804 20916 20814
rect 21532 20804 21588 20860
rect 20860 20802 21588 20804
rect 20860 20750 20862 20802
rect 20914 20750 21588 20802
rect 20860 20748 21588 20750
rect 20860 20738 20916 20748
rect 20748 19506 20804 19516
rect 20860 20020 20916 20030
rect 20972 20020 21028 20748
rect 21420 20580 21476 20590
rect 21084 20020 21140 20030
rect 20972 20018 21140 20020
rect 20972 19966 21086 20018
rect 21138 19966 21140 20018
rect 20972 19964 21140 19966
rect 20860 19906 20916 19964
rect 20860 19854 20862 19906
rect 20914 19854 20916 19906
rect 20524 19292 20804 19348
rect 20300 18610 20356 18620
rect 20524 19012 20580 19022
rect 20188 17948 20356 18004
rect 19852 17502 19854 17554
rect 19906 17502 19908 17554
rect 19852 17490 19908 17502
rect 20188 17668 20244 17678
rect 19628 17388 19796 17444
rect 19628 16996 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16940 19796 16996
rect 19628 16772 19684 16782
rect 19516 16770 19684 16772
rect 19516 16718 19630 16770
rect 19682 16718 19684 16770
rect 19516 16716 19684 16718
rect 19628 16706 19684 16716
rect 19740 15988 19796 16940
rect 19628 15932 19796 15988
rect 19628 13634 19684 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15540 19796 15550
rect 19740 14418 19796 15484
rect 20188 15314 20244 17612
rect 20188 15262 20190 15314
rect 20242 15262 20244 15314
rect 20188 15250 20244 15262
rect 20300 15204 20356 17948
rect 20300 15138 20356 15148
rect 19740 14366 19742 14418
rect 19794 14366 19796 14418
rect 19740 14354 19796 14366
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13582 19630 13634
rect 19682 13582 19684 13634
rect 19628 13570 19684 13582
rect 19292 13076 19348 13086
rect 19292 12982 19348 13020
rect 20524 12850 20580 18956
rect 20748 18004 20804 19292
rect 20860 18452 20916 19854
rect 20860 18386 20916 18396
rect 20748 17948 21028 18004
rect 20636 17442 20692 17454
rect 20636 17390 20638 17442
rect 20690 17390 20692 17442
rect 20636 13858 20692 17390
rect 20636 13806 20638 13858
rect 20690 13806 20692 13858
rect 20636 13794 20692 13806
rect 20860 15314 20916 15326
rect 20860 15262 20862 15314
rect 20914 15262 20916 15314
rect 20860 13636 20916 15262
rect 20972 13860 21028 17948
rect 21084 17668 21140 19964
rect 21420 19346 21476 20524
rect 21644 20244 21700 23772
rect 22428 23828 22484 23838
rect 22428 23734 22484 23772
rect 22540 23714 22596 23726
rect 22540 23662 22542 23714
rect 22594 23662 22596 23714
rect 22540 23378 22596 23662
rect 22540 23326 22542 23378
rect 22594 23326 22596 23378
rect 22540 23314 22596 23326
rect 23212 23380 23268 23884
rect 23324 23938 23380 23996
rect 23324 23886 23326 23938
rect 23378 23886 23380 23938
rect 23324 23874 23380 23886
rect 23660 23604 23716 25116
rect 23324 23380 23380 23390
rect 23212 23378 23380 23380
rect 23212 23326 23326 23378
rect 23378 23326 23380 23378
rect 23212 23324 23380 23326
rect 23324 23314 23380 23324
rect 23548 23044 23604 23054
rect 23548 22950 23604 22988
rect 21868 22370 21924 22382
rect 21868 22318 21870 22370
rect 21922 22318 21924 22370
rect 21868 22260 21924 22318
rect 21868 22194 21924 22204
rect 23436 21588 23492 21598
rect 23436 21494 23492 21532
rect 23660 20804 23716 23548
rect 23884 23828 23940 26238
rect 23996 26178 24052 26190
rect 23996 26126 23998 26178
rect 24050 26126 24052 26178
rect 23996 24946 24052 26126
rect 24556 25508 24612 25518
rect 24556 25414 24612 25452
rect 25004 25506 25060 26908
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 25004 25442 25060 25454
rect 25116 26290 25172 27132
rect 26796 26964 26852 30268
rect 26908 30258 26964 30268
rect 28140 30212 28196 30222
rect 27916 30100 27972 30110
rect 27916 30006 27972 30044
rect 27580 29540 27636 29550
rect 27580 29446 27636 29484
rect 27916 29426 27972 29438
rect 27916 29374 27918 29426
rect 27970 29374 27972 29426
rect 27020 29314 27076 29326
rect 27020 29262 27022 29314
rect 27074 29262 27076 29314
rect 27020 28644 27076 29262
rect 27356 29314 27412 29326
rect 27356 29262 27358 29314
rect 27410 29262 27412 29314
rect 27020 28578 27076 28588
rect 27132 28756 27188 28766
rect 27132 27858 27188 28700
rect 27356 28084 27412 29262
rect 27356 28018 27412 28028
rect 27132 27806 27134 27858
rect 27186 27806 27188 27858
rect 27132 27794 27188 27806
rect 27468 27860 27524 27870
rect 27468 27766 27524 27804
rect 26796 26898 26852 26908
rect 27580 27188 27636 27198
rect 25788 26850 25844 26862
rect 25788 26798 25790 26850
rect 25842 26798 25844 26850
rect 25116 26238 25118 26290
rect 25170 26238 25172 26290
rect 25116 25508 25172 26238
rect 25676 26292 25732 26302
rect 25676 26198 25732 26236
rect 25116 25442 25172 25452
rect 25676 25508 25732 25518
rect 23996 24894 23998 24946
rect 24050 24894 24052 24946
rect 23996 24882 24052 24894
rect 24780 24948 24836 24958
rect 24780 24854 24836 24892
rect 25676 24722 25732 25452
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 25676 24658 25732 24670
rect 23884 23268 23940 23772
rect 24332 23604 24388 23614
rect 24332 23378 24388 23548
rect 24332 23326 24334 23378
rect 24386 23326 24388 23378
rect 24332 23314 24388 23326
rect 23884 23174 23940 23212
rect 24556 23268 24612 23278
rect 24444 22372 24500 22382
rect 24332 22146 24388 22158
rect 24332 22094 24334 22146
rect 24386 22094 24388 22146
rect 24332 21698 24388 22094
rect 24332 21646 24334 21698
rect 24386 21646 24388 21698
rect 24332 21634 24388 21646
rect 23884 21586 23940 21598
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 20916 23940 21534
rect 23884 20850 23940 20860
rect 23660 20710 23716 20748
rect 24444 20802 24500 22316
rect 24556 21586 24612 23212
rect 25788 23042 25844 26798
rect 26012 25396 26068 25406
rect 26012 23268 26068 25340
rect 27244 25282 27300 25294
rect 27244 25230 27246 25282
rect 27298 25230 27300 25282
rect 26348 24722 26404 24734
rect 26348 24670 26350 24722
rect 26402 24670 26404 24722
rect 26348 24052 26404 24670
rect 26348 23986 26404 23996
rect 26572 24164 26628 24174
rect 26572 23378 26628 24108
rect 27244 24164 27300 25230
rect 27244 24098 27300 24108
rect 26572 23326 26574 23378
rect 26626 23326 26628 23378
rect 26572 23314 26628 23326
rect 26796 23826 26852 23838
rect 26796 23774 26798 23826
rect 26850 23774 26852 23826
rect 26796 23604 26852 23774
rect 26012 23174 26068 23212
rect 26684 23156 26740 23166
rect 26684 23062 26740 23100
rect 25788 22990 25790 23042
rect 25842 22990 25844 23042
rect 25788 22978 25844 22990
rect 25004 22372 25060 22382
rect 25060 22316 25172 22372
rect 25004 22278 25060 22316
rect 24892 22148 24948 22158
rect 24892 22054 24948 22092
rect 25116 21700 25172 22316
rect 25676 22370 25732 22382
rect 25676 22318 25678 22370
rect 25730 22318 25732 22370
rect 25340 21700 25396 21710
rect 25116 21644 25340 21700
rect 24556 21534 24558 21586
rect 24610 21534 24612 21586
rect 24556 21522 24612 21534
rect 25340 21586 25396 21644
rect 25340 21534 25342 21586
rect 25394 21534 25396 21586
rect 25340 21522 25396 21534
rect 25676 21252 25732 22318
rect 25676 21186 25732 21196
rect 25788 21700 25844 21710
rect 24444 20750 24446 20802
rect 24498 20750 24500 20802
rect 24444 20738 24500 20750
rect 25116 20802 25172 20814
rect 25116 20750 25118 20802
rect 25170 20750 25172 20802
rect 21644 20188 21924 20244
rect 21756 20020 21812 20030
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21532 20018 21812 20020
rect 21532 19966 21758 20018
rect 21810 19966 21812 20018
rect 21532 19964 21812 19966
rect 21084 16882 21140 17612
rect 21532 17556 21588 19964
rect 21756 19954 21812 19964
rect 21868 19796 21924 20188
rect 23996 20130 24052 20142
rect 23996 20078 23998 20130
rect 24050 20078 24052 20130
rect 21756 19740 21924 19796
rect 23100 19908 23156 19918
rect 21756 19346 21812 19740
rect 21756 19294 21758 19346
rect 21810 19294 21812 19346
rect 21756 19282 21812 19294
rect 23100 19122 23156 19852
rect 23100 19070 23102 19122
rect 23154 19070 23156 19122
rect 23100 19058 23156 19070
rect 22316 19012 22372 19022
rect 22316 18918 22372 18956
rect 22092 18564 22148 18574
rect 21644 18562 22148 18564
rect 21644 18510 22094 18562
rect 22146 18510 22148 18562
rect 21644 18508 22148 18510
rect 21644 17778 21700 18508
rect 22092 18498 22148 18508
rect 23996 18562 24052 20078
rect 24780 19796 24836 19806
rect 23996 18510 23998 18562
rect 24050 18510 24052 18562
rect 23996 18498 24052 18510
rect 24668 19794 24836 19796
rect 24668 19742 24782 19794
rect 24834 19742 24836 19794
rect 24668 19740 24836 19742
rect 22540 18452 22596 18462
rect 21644 17726 21646 17778
rect 21698 17726 21700 17778
rect 21644 17714 21700 17726
rect 21868 17780 21924 17790
rect 21868 17686 21924 17724
rect 22540 17780 22596 18396
rect 23660 18452 23716 18462
rect 23660 18358 23716 18396
rect 24332 18452 24388 18462
rect 23324 18340 23380 18350
rect 23212 18338 23380 18340
rect 23212 18286 23326 18338
rect 23378 18286 23380 18338
rect 23212 18284 23380 18286
rect 22540 17686 22596 17724
rect 22876 18226 22932 18238
rect 22876 18174 22878 18226
rect 22930 18174 22932 18226
rect 22764 17668 22820 17678
rect 22764 17574 22820 17612
rect 21532 17490 21588 17500
rect 22204 17554 22260 17566
rect 22204 17502 22206 17554
rect 22258 17502 22260 17554
rect 21084 16830 21086 16882
rect 21138 16830 21140 16882
rect 21084 16818 21140 16830
rect 21756 16882 21812 16894
rect 21756 16830 21758 16882
rect 21810 16830 21812 16882
rect 21756 15988 21812 16830
rect 21756 15922 21812 15932
rect 21980 15988 22036 15998
rect 22204 15988 22260 17502
rect 21980 15986 22260 15988
rect 21980 15934 21982 15986
rect 22034 15934 22260 15986
rect 21980 15932 22260 15934
rect 22428 17556 22484 17566
rect 21980 15922 22036 15932
rect 21196 15874 21252 15886
rect 21196 15822 21198 15874
rect 21250 15822 21252 15874
rect 21196 15148 21252 15822
rect 21196 15092 21588 15148
rect 21308 13860 21364 13870
rect 20972 13858 21364 13860
rect 20972 13806 21310 13858
rect 21362 13806 21364 13858
rect 20972 13804 21364 13806
rect 21308 13794 21364 13804
rect 20860 13570 20916 13580
rect 20524 12798 20526 12850
rect 20578 12798 20580 12850
rect 20524 12786 20580 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19068 12014 19070 12066
rect 19122 12014 19124 12066
rect 19068 12002 19124 12014
rect 21532 11282 21588 15092
rect 22428 13634 22484 17500
rect 22876 16660 22932 18174
rect 22876 16594 22932 16604
rect 22428 13582 22430 13634
rect 22482 13582 22484 13634
rect 22428 13570 22484 13582
rect 22652 15988 22708 15998
rect 22652 11506 22708 15932
rect 23212 15538 23268 18284
rect 23324 18274 23380 18284
rect 23436 17666 23492 17678
rect 23436 17614 23438 17666
rect 23490 17614 23492 17666
rect 23436 15876 23492 17614
rect 24108 17106 24164 17118
rect 24108 17054 24110 17106
rect 24162 17054 24164 17106
rect 23436 15810 23492 15820
rect 23660 16660 23716 16670
rect 23212 15486 23214 15538
rect 23266 15486 23268 15538
rect 23212 15474 23268 15486
rect 23660 15148 23716 16604
rect 23996 16100 24052 16110
rect 22876 15092 22932 15102
rect 23660 15092 23828 15148
rect 22876 12850 22932 15036
rect 22876 12798 22878 12850
rect 22930 12798 22932 12850
rect 22876 12786 22932 12798
rect 22988 13636 23044 13646
rect 22988 12066 23044 13580
rect 23772 12292 23828 15092
rect 23884 15092 23940 15102
rect 23884 14998 23940 15036
rect 23884 14644 23940 14654
rect 23884 13074 23940 14588
rect 23996 14530 24052 16044
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 23996 14466 24052 14478
rect 24108 13860 24164 17054
rect 24220 16098 24276 16110
rect 24220 16046 24222 16098
rect 24274 16046 24276 16098
rect 24220 14644 24276 16046
rect 24332 15426 24388 18396
rect 24668 15876 24724 19740
rect 24780 19730 24836 19740
rect 25116 19572 25172 20750
rect 25452 20020 25508 20030
rect 25340 20018 25508 20020
rect 25340 19966 25454 20018
rect 25506 19966 25508 20018
rect 25340 19964 25508 19966
rect 25228 19908 25284 19918
rect 25228 19814 25284 19852
rect 25116 19506 25172 19516
rect 25340 18452 25396 19964
rect 25452 19954 25508 19964
rect 25452 19236 25508 19246
rect 25788 19236 25844 21644
rect 26012 21586 26068 21598
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 26012 19908 26068 21534
rect 26796 20916 26852 23548
rect 26908 23154 26964 23166
rect 26908 23102 26910 23154
rect 26962 23102 26964 23154
rect 26908 21700 26964 23102
rect 27580 23154 27636 27132
rect 27916 27076 27972 29374
rect 28140 28756 28196 30156
rect 28252 29540 28308 32508
rect 28364 33122 28420 33134
rect 28364 33070 28366 33122
rect 28418 33070 28420 33122
rect 28364 31220 28420 33070
rect 28700 31890 28756 33180
rect 28700 31838 28702 31890
rect 28754 31838 28756 31890
rect 28700 31826 28756 31838
rect 28924 31444 28980 34188
rect 30268 34242 30324 34254
rect 30268 34190 30270 34242
rect 30322 34190 30324 34242
rect 29036 34018 29092 34030
rect 29036 33966 29038 34018
rect 29090 33966 29092 34018
rect 29036 33348 29092 33966
rect 29036 33282 29092 33292
rect 30156 33458 30212 33470
rect 30156 33406 30158 33458
rect 30210 33406 30212 33458
rect 29036 33124 29092 33134
rect 29036 31890 29092 33068
rect 29820 33012 29876 33022
rect 29708 32786 29764 32798
rect 29708 32734 29710 32786
rect 29762 32734 29764 32786
rect 29708 32676 29764 32734
rect 29708 32610 29764 32620
rect 29036 31838 29038 31890
rect 29090 31838 29092 31890
rect 29036 31826 29092 31838
rect 29820 31666 29876 32956
rect 29820 31614 29822 31666
rect 29874 31614 29876 31666
rect 29820 31602 29876 31614
rect 30044 31780 30100 31790
rect 28924 31388 29092 31444
rect 28924 31220 28980 31230
rect 28364 31218 28980 31220
rect 28364 31166 28926 31218
rect 28978 31166 28980 31218
rect 28364 31164 28980 31166
rect 28924 31154 28980 31164
rect 28252 29474 28308 29484
rect 28476 30660 28532 30670
rect 28476 29426 28532 30604
rect 28476 29374 28478 29426
rect 28530 29374 28532 29426
rect 28476 29362 28532 29374
rect 29036 28866 29092 31388
rect 29820 31332 29876 31342
rect 29708 31108 29764 31118
rect 29708 31014 29764 31052
rect 29260 30212 29316 30222
rect 29260 30118 29316 30156
rect 29708 30212 29764 30222
rect 29820 30212 29876 31276
rect 30044 31220 30100 31724
rect 30044 31126 30100 31164
rect 30156 30660 30212 33406
rect 30268 33124 30324 34190
rect 30268 33058 30324 33068
rect 30268 32788 30324 32798
rect 30380 32788 30436 34748
rect 31500 34738 31556 34748
rect 30828 34020 30884 34030
rect 30268 32786 30436 32788
rect 30268 32734 30270 32786
rect 30322 32734 30436 32786
rect 30268 32732 30436 32734
rect 30716 34018 30884 34020
rect 30716 33966 30830 34018
rect 30882 33966 30884 34018
rect 30716 33964 30884 33966
rect 30268 32722 30324 32732
rect 30492 32676 30548 32686
rect 30492 32582 30548 32620
rect 30716 32564 30772 33964
rect 30828 33954 30884 33964
rect 31052 34018 31108 34030
rect 31052 33966 31054 34018
rect 31106 33966 31108 34018
rect 31052 33012 31108 33966
rect 31164 33236 31220 33246
rect 31164 33142 31220 33180
rect 31052 32946 31108 32956
rect 30716 32470 30772 32508
rect 31388 32564 31444 32574
rect 31388 32470 31444 32508
rect 31836 32564 31892 32574
rect 31892 32508 32004 32564
rect 31836 32470 31892 32508
rect 31164 32452 31220 32462
rect 31164 32358 31220 32396
rect 31948 31332 32004 32508
rect 32060 31778 32116 34972
rect 32620 34962 32676 34972
rect 33404 34244 33460 34254
rect 32732 34242 33460 34244
rect 32732 34190 33406 34242
rect 33458 34190 33460 34242
rect 32732 34188 33460 34190
rect 32060 31726 32062 31778
rect 32114 31726 32116 31778
rect 32060 31714 32116 31726
rect 32172 32450 32228 32462
rect 32172 32398 32174 32450
rect 32226 32398 32228 32450
rect 31948 31276 32116 31332
rect 31500 31220 31556 31230
rect 30940 30884 30996 30922
rect 30940 30818 30996 30828
rect 30156 30594 30212 30604
rect 30940 30660 30996 30670
rect 29708 30210 29876 30212
rect 29708 30158 29710 30210
rect 29762 30158 29876 30210
rect 29708 30156 29876 30158
rect 29708 30146 29764 30156
rect 30604 29764 30660 29774
rect 29036 28814 29038 28866
rect 29090 28814 29092 28866
rect 29036 28802 29092 28814
rect 29820 29316 29876 29326
rect 28140 28662 28196 28700
rect 29820 28530 29876 29260
rect 29820 28478 29822 28530
rect 29874 28478 29876 28530
rect 29820 28466 29876 28478
rect 29820 28084 29876 28094
rect 29820 27990 29876 28028
rect 30604 28082 30660 29708
rect 30940 29650 30996 30604
rect 30940 29598 30942 29650
rect 30994 29598 30996 29650
rect 30940 29586 30996 29598
rect 31500 29650 31556 31164
rect 31948 31108 32004 31118
rect 31948 31014 32004 31052
rect 31500 29598 31502 29650
rect 31554 29598 31556 29650
rect 31500 29586 31556 29598
rect 31612 29652 31668 29662
rect 30604 28030 30606 28082
rect 30658 28030 30660 28082
rect 30604 28018 30660 28030
rect 31500 28084 31556 28094
rect 31612 28084 31668 29596
rect 32060 29652 32116 31276
rect 32172 29986 32228 32398
rect 32508 31778 32564 31790
rect 32508 31726 32510 31778
rect 32562 31726 32564 31778
rect 32396 31444 32452 31454
rect 32396 30660 32452 31388
rect 32396 30594 32452 30604
rect 32396 30324 32452 30334
rect 32172 29934 32174 29986
rect 32226 29934 32228 29986
rect 32172 29922 32228 29934
rect 32284 30268 32396 30324
rect 32060 29538 32116 29596
rect 32060 29486 32062 29538
rect 32114 29486 32116 29538
rect 32060 29474 32116 29486
rect 31724 29316 31780 29326
rect 31724 29222 31780 29260
rect 32172 28644 32228 28654
rect 32284 28644 32340 30268
rect 32396 30258 32452 30268
rect 32172 28642 32340 28644
rect 32172 28590 32174 28642
rect 32226 28590 32340 28642
rect 32172 28588 32340 28590
rect 32508 30212 32564 31726
rect 32508 28644 32564 30156
rect 32732 30210 32788 34188
rect 33404 34178 33460 34188
rect 34524 34020 34580 34030
rect 33628 34018 34580 34020
rect 33628 33966 34526 34018
rect 34578 33966 34580 34018
rect 33628 33964 34580 33966
rect 33180 33458 33236 33470
rect 33180 33406 33182 33458
rect 33234 33406 33236 33458
rect 32956 32676 33012 32686
rect 32732 30158 32734 30210
rect 32786 30158 32788 30210
rect 32732 30146 32788 30158
rect 32844 30772 32900 30782
rect 32844 30210 32900 30716
rect 32844 30158 32846 30210
rect 32898 30158 32900 30210
rect 32844 30146 32900 30158
rect 32844 28644 32900 28654
rect 32508 28642 32900 28644
rect 32508 28590 32510 28642
rect 32562 28590 32846 28642
rect 32898 28590 32900 28642
rect 32508 28588 32900 28590
rect 32172 28578 32228 28588
rect 32508 28578 32564 28588
rect 32844 28578 32900 28588
rect 31500 28082 31668 28084
rect 31500 28030 31502 28082
rect 31554 28030 31668 28082
rect 31500 28028 31668 28030
rect 31500 28018 31556 28028
rect 30268 27860 30324 27870
rect 27916 27010 27972 27020
rect 28140 27074 28196 27086
rect 28140 27022 28142 27074
rect 28194 27022 28196 27074
rect 28140 25620 28196 27022
rect 28700 27076 28756 27086
rect 28700 26982 28756 27020
rect 30156 27076 30212 27086
rect 30268 27076 30324 27804
rect 31836 27860 31892 27870
rect 31836 27766 31892 27804
rect 31836 27636 31892 27646
rect 30156 27074 30324 27076
rect 30156 27022 30158 27074
rect 30210 27022 30324 27074
rect 30156 27020 30324 27022
rect 30156 27010 30212 27020
rect 29372 26964 29428 26974
rect 28140 25554 28196 25564
rect 28252 26514 28308 26526
rect 28252 26462 28254 26514
rect 28306 26462 28308 26514
rect 28252 25618 28308 26462
rect 29036 26290 29092 26302
rect 29036 26238 29038 26290
rect 29090 26238 29092 26290
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 28812 26066 28868 26078
rect 28812 26014 28814 26066
rect 28866 26014 28868 26066
rect 28588 25396 28644 25406
rect 28588 25302 28644 25340
rect 28028 25282 28084 25294
rect 28028 25230 28030 25282
rect 28082 25230 28084 25282
rect 28028 24500 28084 25230
rect 28028 24434 28084 24444
rect 28588 24834 28644 24846
rect 28588 24782 28590 24834
rect 28642 24782 28644 24834
rect 28588 23268 28644 24782
rect 28812 23828 28868 26014
rect 28812 23762 28868 23772
rect 29036 23940 29092 26238
rect 29372 24946 29428 26908
rect 30156 25620 30212 25630
rect 29596 25396 29652 25406
rect 29596 25302 29652 25340
rect 29372 24894 29374 24946
rect 29426 24894 29428 24946
rect 29372 24882 29428 24894
rect 30044 24276 30100 24286
rect 29260 23940 29316 23950
rect 29036 23938 29316 23940
rect 29036 23886 29262 23938
rect 29314 23886 29316 23938
rect 29036 23884 29316 23886
rect 28588 23202 28644 23212
rect 29036 23716 29092 23884
rect 29260 23874 29316 23884
rect 27580 23102 27582 23154
rect 27634 23102 27636 23154
rect 27580 23090 27636 23102
rect 29036 23044 29092 23660
rect 30044 23378 30100 24220
rect 30156 24050 30212 25564
rect 30268 25396 30324 27020
rect 31388 27076 31444 27086
rect 31388 26178 31444 27020
rect 31836 27076 31892 27580
rect 31836 26982 31892 27020
rect 32956 26514 33012 32620
rect 33068 32450 33124 32462
rect 33068 32398 33070 32450
rect 33122 32398 33124 32450
rect 33068 31444 33124 32398
rect 33068 31378 33124 31388
rect 33180 31332 33236 33406
rect 33292 32564 33348 32574
rect 33292 31892 33348 32508
rect 33292 31826 33348 31836
rect 33180 31266 33236 31276
rect 33068 30994 33124 31006
rect 33068 30942 33070 30994
rect 33122 30942 33124 30994
rect 33068 29428 33124 30942
rect 33628 30994 33684 33964
rect 34524 33954 34580 33964
rect 34076 33234 34132 33246
rect 34076 33182 34078 33234
rect 34130 33182 34132 33234
rect 33852 32676 33908 32686
rect 33852 32582 33908 32620
rect 33628 30942 33630 30994
rect 33682 30942 33684 30994
rect 33628 30930 33684 30942
rect 33964 31890 34020 31902
rect 33964 31838 33966 31890
rect 34018 31838 34020 31890
rect 33516 30884 33572 30894
rect 33404 30828 33516 30884
rect 33180 29652 33236 29662
rect 33180 29538 33236 29596
rect 33180 29486 33182 29538
rect 33234 29486 33236 29538
rect 33180 29474 33236 29486
rect 33068 29362 33124 29372
rect 33404 28642 33460 30828
rect 33516 30818 33572 30828
rect 33964 30324 34020 31838
rect 34076 31220 34132 33182
rect 34636 31780 34692 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35644 32676 35700 32686
rect 35196 32452 35252 32462
rect 35196 32450 35588 32452
rect 35196 32398 35198 32450
rect 35250 32398 35588 32450
rect 35196 32396 35588 32398
rect 35196 32386 35252 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34636 31714 34692 31724
rect 34076 31154 34132 31164
rect 34972 31666 35028 31678
rect 34972 31614 34974 31666
rect 35026 31614 35028 31666
rect 33964 30258 34020 30268
rect 33516 29986 33572 29998
rect 33516 29934 33518 29986
rect 33570 29934 33572 29986
rect 33516 29538 33572 29934
rect 33516 29486 33518 29538
rect 33570 29486 33572 29538
rect 33516 29474 33572 29486
rect 34300 29876 34356 29886
rect 33852 29428 33908 29438
rect 33404 28590 33406 28642
rect 33458 28590 33460 28642
rect 33404 28578 33460 28590
rect 33516 28756 33572 28766
rect 32956 26462 32958 26514
rect 33010 26462 33012 26514
rect 32956 26450 33012 26462
rect 31388 26126 31390 26178
rect 31442 26126 31444 26178
rect 31052 25508 31108 25518
rect 30940 25506 31108 25508
rect 30940 25454 31054 25506
rect 31106 25454 31108 25506
rect 30940 25452 31108 25454
rect 31388 25508 31444 26126
rect 32172 26292 32228 26302
rect 31612 25508 31668 25518
rect 31388 25506 31668 25508
rect 31388 25454 31614 25506
rect 31666 25454 31668 25506
rect 31388 25452 31668 25454
rect 30380 25396 30436 25406
rect 30268 25394 30436 25396
rect 30268 25342 30382 25394
rect 30434 25342 30436 25394
rect 30268 25340 30436 25342
rect 30380 24612 30436 25340
rect 30380 24546 30436 24556
rect 30828 25394 30884 25406
rect 30828 25342 30830 25394
rect 30882 25342 30884 25394
rect 30828 24276 30884 25342
rect 30828 24210 30884 24220
rect 30156 23998 30158 24050
rect 30210 23998 30212 24050
rect 30156 23986 30212 23998
rect 30044 23326 30046 23378
rect 30098 23326 30100 23378
rect 30044 23314 30100 23326
rect 30604 23604 30660 23614
rect 30604 23378 30660 23548
rect 30604 23326 30606 23378
rect 30658 23326 30660 23378
rect 30604 23314 30660 23326
rect 30940 23156 30996 25452
rect 31052 25442 31108 25452
rect 31612 25442 31668 25452
rect 32172 24722 32228 26236
rect 32284 25508 32340 25518
rect 32284 25414 32340 25452
rect 32956 25284 33012 25294
rect 32956 24724 33012 25228
rect 32172 24670 32174 24722
rect 32226 24670 32228 24722
rect 32172 24658 32228 24670
rect 32844 24722 33012 24724
rect 32844 24670 32958 24722
rect 33010 24670 33012 24722
rect 32844 24668 33012 24670
rect 33516 24724 33572 28700
rect 33852 27858 33908 29372
rect 33852 27806 33854 27858
rect 33906 27806 33908 27858
rect 33852 27794 33908 27806
rect 33964 27972 34020 27982
rect 33740 26404 33796 26414
rect 33740 26310 33796 26348
rect 33964 26292 34020 27916
rect 34300 27858 34356 29820
rect 34972 29764 35028 31614
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34972 29698 35028 29708
rect 35308 30212 35364 30222
rect 35308 29428 35364 30156
rect 35532 29876 35588 32396
rect 35532 29810 35588 29820
rect 35644 29652 35700 32620
rect 35756 31892 35812 31902
rect 35756 31798 35812 31836
rect 35868 31554 35924 31566
rect 35868 31502 35870 31554
rect 35922 31502 35924 31554
rect 35868 31218 35924 31502
rect 35868 31166 35870 31218
rect 35922 31166 35924 31218
rect 35868 31154 35924 31166
rect 35980 30996 36036 31006
rect 35308 29334 35364 29372
rect 35532 29596 35700 29652
rect 35756 30436 35812 30446
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34300 27806 34302 27858
rect 34354 27806 34356 27858
rect 34300 27794 34356 27806
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34524 27188 34580 27198
rect 35532 27188 35588 29596
rect 35756 29426 35812 30380
rect 35980 30210 36036 30940
rect 35980 30158 35982 30210
rect 36034 30158 36036 30210
rect 35980 30146 36036 30158
rect 35756 29374 35758 29426
rect 35810 29374 35812 29426
rect 35756 29362 35812 29374
rect 35980 28420 36036 28430
rect 35980 28326 36036 28364
rect 36316 28196 36372 38892
rect 38108 37378 38164 37390
rect 38108 37326 38110 37378
rect 38162 37326 38164 37378
rect 37436 36370 37492 36382
rect 37436 36318 37438 36370
rect 37490 36318 37492 36370
rect 37212 35028 37268 35038
rect 36652 33572 36708 33582
rect 36652 31218 36708 33516
rect 36652 31166 36654 31218
rect 36706 31166 36708 31218
rect 36652 31154 36708 31166
rect 36764 33460 36820 33470
rect 36540 31108 36596 31118
rect 36428 31052 36540 31108
rect 36428 28868 36484 31052
rect 36540 31042 36596 31052
rect 36540 30212 36596 30222
rect 36540 30118 36596 30156
rect 36540 28868 36596 28878
rect 36428 28866 36596 28868
rect 36428 28814 36542 28866
rect 36594 28814 36596 28866
rect 36428 28812 36596 28814
rect 36540 28802 36596 28812
rect 36428 28196 36484 28206
rect 36316 28140 36428 28196
rect 36428 28130 36484 28140
rect 36540 27972 36596 27982
rect 35756 27970 36596 27972
rect 35756 27918 36542 27970
rect 36594 27918 36596 27970
rect 35756 27916 36596 27918
rect 35532 27132 35700 27188
rect 34524 27094 34580 27132
rect 33964 26226 34020 26236
rect 34076 27076 34132 27086
rect 33628 24724 33684 24734
rect 33516 24722 33684 24724
rect 33516 24670 33630 24722
rect 33682 24670 33684 24722
rect 33516 24668 33684 24670
rect 31052 24612 31108 24622
rect 31052 23940 31108 24556
rect 31052 23874 31108 23884
rect 32060 23940 32116 23950
rect 31164 23828 31220 23838
rect 31164 23734 31220 23772
rect 32060 23266 32116 23884
rect 32060 23214 32062 23266
rect 32114 23214 32116 23266
rect 32060 23202 32116 23214
rect 31052 23156 31108 23166
rect 30940 23100 31052 23156
rect 28588 22988 29092 23044
rect 31052 23042 31108 23100
rect 32508 23156 32564 23166
rect 31052 22990 31054 23042
rect 31106 22990 31108 23042
rect 28028 22146 28084 22158
rect 28028 22094 28030 22146
rect 28082 22094 28084 22146
rect 26908 21634 26964 21644
rect 27356 21924 27412 21934
rect 26796 20850 26852 20860
rect 27132 21252 27188 21262
rect 26012 19842 26068 19852
rect 26908 20130 26964 20142
rect 26908 20078 26910 20130
rect 26962 20078 26964 20130
rect 25452 19234 25620 19236
rect 25452 19182 25454 19234
rect 25506 19182 25620 19234
rect 25452 19180 25620 19182
rect 25452 19170 25508 19180
rect 25340 17556 25396 18396
rect 25340 17490 25396 17500
rect 25564 17220 25620 19180
rect 25788 19142 25844 19180
rect 26124 19794 26180 19806
rect 26124 19742 26126 19794
rect 26178 19742 26180 19794
rect 25676 18450 25732 18462
rect 25676 18398 25678 18450
rect 25730 18398 25732 18450
rect 25676 18228 25732 18398
rect 25676 18162 25732 18172
rect 25900 17444 25956 17454
rect 25900 17442 26068 17444
rect 25900 17390 25902 17442
rect 25954 17390 26068 17442
rect 25900 17388 26068 17390
rect 25900 17378 25956 17388
rect 25564 17164 25844 17220
rect 24780 16660 24836 16670
rect 25116 16660 25172 16670
rect 24780 16566 24836 16604
rect 25004 16658 25172 16660
rect 25004 16606 25118 16658
rect 25170 16606 25172 16658
rect 25004 16604 25172 16606
rect 24892 16100 24948 16110
rect 24892 16006 24948 16044
rect 24668 15820 24948 15876
rect 24332 15374 24334 15426
rect 24386 15374 24388 15426
rect 24332 15148 24388 15374
rect 24668 15652 24724 15662
rect 24668 15426 24724 15596
rect 24668 15374 24670 15426
rect 24722 15374 24724 15426
rect 24668 15362 24724 15374
rect 24332 15092 24612 15148
rect 24220 14578 24276 14588
rect 24444 14530 24500 14542
rect 24444 14478 24446 14530
rect 24498 14478 24500 14530
rect 24332 13860 24388 13870
rect 24108 13858 24388 13860
rect 24108 13806 24334 13858
rect 24386 13806 24388 13858
rect 24108 13804 24388 13806
rect 24332 13794 24388 13804
rect 23884 13022 23886 13074
rect 23938 13022 23940 13074
rect 23884 13010 23940 13022
rect 23996 12292 24052 12302
rect 23772 12290 24052 12292
rect 23772 12238 23998 12290
rect 24050 12238 24052 12290
rect 23772 12236 24052 12238
rect 23996 12226 24052 12236
rect 22988 12014 22990 12066
rect 23042 12014 23044 12066
rect 22988 12002 23044 12014
rect 22652 11454 22654 11506
rect 22706 11454 22708 11506
rect 22652 11442 22708 11454
rect 21532 11230 21534 11282
rect 21586 11230 21588 11282
rect 21532 11218 21588 11230
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 11788 10670 11790 10722
rect 11842 10670 11844 10722
rect 11788 10658 11844 10670
rect 24444 10500 24500 14478
rect 24556 13746 24612 15092
rect 24892 15092 24948 15820
rect 24892 15026 24948 15036
rect 24556 13694 24558 13746
rect 24610 13694 24612 13746
rect 24556 13682 24612 13694
rect 25004 13412 25060 16604
rect 25116 16594 25172 16604
rect 25116 16100 25172 16138
rect 25116 16034 25172 16044
rect 25676 16098 25732 16110
rect 25676 16046 25678 16098
rect 25730 16046 25732 16098
rect 25004 13346 25060 13356
rect 25116 15876 25172 15886
rect 25116 11508 25172 15820
rect 25676 12068 25732 16046
rect 25788 13076 25844 17164
rect 25900 16994 25956 17006
rect 25900 16942 25902 16994
rect 25954 16942 25956 16994
rect 25900 15540 25956 16942
rect 26012 15652 26068 17388
rect 26012 15586 26068 15596
rect 25900 15474 25956 15484
rect 26124 13860 26180 19742
rect 26908 18452 26964 20078
rect 26908 18386 26964 18396
rect 26684 17554 26740 17566
rect 26684 17502 26686 17554
rect 26738 17502 26740 17554
rect 26460 17442 26516 17454
rect 26460 17390 26462 17442
rect 26514 17390 26516 17442
rect 26236 16660 26292 16670
rect 26292 16604 26404 16660
rect 26236 16594 26292 16604
rect 26236 15204 26292 15242
rect 26236 15138 26292 15148
rect 26124 13794 26180 13804
rect 26348 13188 26404 16604
rect 26460 15428 26516 17390
rect 26460 15362 26516 15372
rect 26684 14418 26740 17502
rect 27020 17556 27076 17566
rect 27020 17462 27076 17500
rect 26684 14366 26686 14418
rect 26738 14366 26740 14418
rect 26684 14354 26740 14366
rect 27132 13634 27188 21196
rect 27356 15426 27412 21868
rect 27804 20916 27860 20926
rect 27580 20578 27636 20590
rect 27580 20526 27582 20578
rect 27634 20526 27636 20578
rect 27580 19348 27636 20526
rect 27580 19282 27636 19292
rect 27804 19346 27860 20860
rect 28028 19796 28084 22094
rect 28476 21810 28532 21822
rect 28476 21758 28478 21810
rect 28530 21758 28532 21810
rect 28140 20578 28196 20590
rect 28140 20526 28142 20578
rect 28194 20526 28196 20578
rect 28140 20132 28196 20526
rect 28140 20066 28196 20076
rect 28476 20020 28532 21758
rect 28588 20916 28644 22988
rect 31052 22978 31108 22990
rect 32172 23044 32228 23054
rect 32172 22370 32228 22988
rect 32172 22318 32174 22370
rect 32226 22318 32228 22370
rect 32172 22306 32228 22318
rect 28588 20822 28644 20860
rect 28700 22146 28756 22158
rect 28700 22094 28702 22146
rect 28754 22094 28756 22146
rect 28476 19954 28532 19964
rect 28028 19730 28084 19740
rect 27804 19294 27806 19346
rect 27858 19294 27860 19346
rect 27804 19282 27860 19294
rect 28588 19236 28644 19246
rect 28588 18338 28644 19180
rect 28588 18286 28590 18338
rect 28642 18286 28644 18338
rect 28588 18274 28644 18286
rect 27356 15374 27358 15426
rect 27410 15374 27412 15426
rect 27356 15362 27412 15374
rect 27580 18226 27636 18238
rect 27580 18174 27582 18226
rect 27634 18174 27636 18226
rect 27580 17666 27636 18174
rect 28252 18228 28308 18238
rect 28252 17778 28308 18172
rect 28252 17726 28254 17778
rect 28306 17726 28308 17778
rect 28252 17714 28308 17726
rect 27580 17614 27582 17666
rect 27634 17614 27636 17666
rect 27580 17556 27636 17614
rect 27580 15428 27636 17500
rect 27804 17556 27860 17566
rect 27804 17554 27972 17556
rect 27804 17502 27806 17554
rect 27858 17502 27972 17554
rect 27804 17500 27972 17502
rect 27804 17490 27860 17500
rect 27916 15986 27972 17500
rect 28700 17220 28756 22094
rect 29036 22146 29092 22158
rect 29036 22094 29038 22146
rect 29090 22094 29092 22146
rect 29036 21924 29092 22094
rect 29036 21858 29092 21868
rect 29820 22146 29876 22158
rect 29820 22094 29822 22146
rect 29874 22094 29876 22146
rect 29820 21812 29876 22094
rect 29820 21746 29876 21756
rect 32172 21700 32228 21710
rect 32172 21606 32228 21644
rect 32508 21698 32564 23100
rect 32732 22372 32788 22382
rect 32844 22372 32900 24668
rect 32956 24658 33012 24668
rect 33628 24658 33684 24668
rect 33964 24500 34020 24510
rect 32956 24052 33012 24062
rect 32956 23958 33012 23996
rect 33964 23826 34020 24444
rect 33964 23774 33966 23826
rect 34018 23774 34020 23826
rect 33964 23762 34020 23774
rect 33068 23268 33124 23278
rect 33068 23174 33124 23212
rect 33292 23156 33348 23166
rect 32732 22370 32900 22372
rect 32732 22318 32734 22370
rect 32786 22318 32900 22370
rect 32732 22316 32900 22318
rect 33068 22372 33124 22382
rect 33180 22372 33236 22382
rect 33068 22370 33180 22372
rect 33068 22318 33070 22370
rect 33122 22318 33180 22370
rect 33068 22316 33180 22318
rect 32732 22306 32788 22316
rect 33068 22306 33124 22316
rect 32508 21646 32510 21698
rect 32562 21646 32564 21698
rect 32508 21634 32564 21646
rect 31276 21586 31332 21598
rect 31276 21534 31278 21586
rect 31330 21534 31332 21586
rect 29484 21476 29540 21486
rect 29148 21474 29540 21476
rect 29148 21422 29486 21474
rect 29538 21422 29540 21474
rect 29148 21420 29540 21422
rect 29036 21362 29092 21374
rect 29036 21310 29038 21362
rect 29090 21310 29092 21362
rect 29036 20804 29092 21310
rect 28924 20748 29092 20804
rect 28924 18676 28980 20748
rect 29148 20188 29204 21420
rect 29484 21410 29540 21420
rect 30268 20916 30324 20926
rect 29036 20132 29204 20188
rect 29260 20802 29316 20814
rect 29260 20750 29262 20802
rect 29314 20750 29316 20802
rect 29036 19012 29092 20132
rect 29148 20018 29204 20030
rect 29148 19966 29150 20018
rect 29202 19966 29204 20018
rect 29148 19460 29204 19966
rect 29148 19394 29204 19404
rect 29260 20020 29316 20750
rect 29708 20802 29764 20814
rect 29708 20750 29710 20802
rect 29762 20750 29764 20802
rect 29596 20020 29652 20030
rect 29260 20018 29652 20020
rect 29260 19966 29598 20018
rect 29650 19966 29652 20018
rect 29260 19964 29652 19966
rect 29260 19236 29316 19964
rect 29596 19954 29652 19964
rect 29260 19170 29316 19180
rect 29372 19234 29428 19246
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29372 19012 29428 19182
rect 29036 18956 29428 19012
rect 28924 18610 28980 18620
rect 29372 17668 29428 18956
rect 29708 18564 29764 20750
rect 30044 19460 30100 19470
rect 29820 19234 29876 19246
rect 29820 19182 29822 19234
rect 29874 19182 29876 19234
rect 29820 18788 29876 19182
rect 29820 18722 29876 18732
rect 29708 18498 29764 18508
rect 29372 17612 29652 17668
rect 28700 17164 29428 17220
rect 27916 15934 27918 15986
rect 27970 15934 27972 15986
rect 27916 15922 27972 15934
rect 28252 16882 28308 16894
rect 28252 16830 28254 16882
rect 28306 16830 28308 16882
rect 28140 15540 28196 15550
rect 28140 15446 28196 15484
rect 28028 15428 28084 15438
rect 27580 15426 28084 15428
rect 27580 15374 28030 15426
rect 28082 15374 28084 15426
rect 27580 15372 28084 15374
rect 28028 15362 28084 15372
rect 27916 15204 27972 15214
rect 27132 13582 27134 13634
rect 27186 13582 27188 13634
rect 27132 13570 27188 13582
rect 27244 15092 27300 15102
rect 26348 13132 26740 13188
rect 26236 13076 26292 13086
rect 25788 13074 26292 13076
rect 25788 13022 26238 13074
rect 26290 13022 26292 13074
rect 25788 13020 26292 13022
rect 26236 13010 26292 13020
rect 26572 12068 26628 12078
rect 25676 12066 26628 12068
rect 25676 12014 26574 12066
rect 26626 12014 26628 12066
rect 25676 12012 26628 12014
rect 26572 12002 26628 12012
rect 25228 11508 25284 11518
rect 25116 11506 25284 11508
rect 25116 11454 25230 11506
rect 25282 11454 25284 11506
rect 25116 11452 25284 11454
rect 25228 11442 25284 11452
rect 26572 11284 26628 11294
rect 26684 11284 26740 13132
rect 27244 12850 27300 15036
rect 27244 12798 27246 12850
rect 27298 12798 27300 12850
rect 27244 12786 27300 12798
rect 27468 14306 27524 14318
rect 27468 14254 27470 14306
rect 27522 14254 27524 14306
rect 27468 12292 27524 14254
rect 27468 12226 27524 12236
rect 27580 13412 27636 13422
rect 27580 12290 27636 13356
rect 27580 12238 27582 12290
rect 27634 12238 27636 12290
rect 27580 12226 27636 12238
rect 26572 11282 26740 11284
rect 26572 11230 26574 11282
rect 26626 11230 26740 11282
rect 26572 11228 26740 11230
rect 26572 11218 26628 11228
rect 27916 10722 27972 15148
rect 28028 13860 28084 13870
rect 28028 13766 28084 13804
rect 28252 12068 28308 16830
rect 28812 16884 28868 16894
rect 28924 16884 28980 16894
rect 28812 16882 28924 16884
rect 28812 16830 28814 16882
rect 28866 16830 28924 16882
rect 28812 16828 28924 16830
rect 28812 16818 28868 16828
rect 28924 16100 28980 16828
rect 29036 16100 29092 16110
rect 28980 16098 29092 16100
rect 28980 16046 29038 16098
rect 29090 16046 29092 16098
rect 28980 16044 29092 16046
rect 28700 15876 28756 15886
rect 28700 15874 28868 15876
rect 28700 15822 28702 15874
rect 28754 15822 28868 15874
rect 28700 15820 28868 15822
rect 28700 15810 28756 15820
rect 28252 12002 28308 12012
rect 28476 12740 28532 12750
rect 27916 10670 27918 10722
rect 27970 10670 27972 10722
rect 27916 10658 27972 10670
rect 24444 10434 24500 10444
rect 26572 10500 26628 10510
rect 26572 10406 26628 10444
rect 10556 9938 10724 9940
rect 10556 9886 10558 9938
rect 10610 9886 10724 9938
rect 10556 9884 10724 9886
rect 24108 10052 24164 10062
rect 10556 9874 10612 9884
rect 5292 9650 5348 9660
rect 9212 9716 9268 9726
rect 9212 9622 9268 9660
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2828 8258 2884 8270
rect 2828 8206 2830 8258
rect 2882 8206 2884 8258
rect 2044 8146 2100 8158
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 7476 2100 8094
rect 2828 8036 2884 8206
rect 2828 7970 2884 7980
rect 3388 8036 3444 8046
rect 3388 7942 3444 7980
rect 18396 8036 18452 8046
rect 2044 7410 2100 7420
rect 2940 7474 2996 7486
rect 2940 7422 2942 7474
rect 2994 7422 2996 7474
rect 1932 7362 1988 7374
rect 1932 7310 1934 7362
rect 1986 7310 1988 7362
rect 1932 6804 1988 7310
rect 2940 7364 2996 7422
rect 2940 7298 2996 7308
rect 3500 7364 3556 7374
rect 3500 7270 3556 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 1932 6738 1988 6748
rect 2940 6692 2996 6702
rect 2940 6598 2996 6636
rect 16604 6692 16660 6702
rect 2044 6578 2100 6590
rect 2044 6526 2046 6578
rect 2098 6526 2100 6578
rect 2044 6132 2100 6526
rect 2044 6066 2100 6076
rect 2156 6356 2212 6366
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5460 1988 5742
rect 2156 5572 2212 6300
rect 2940 5908 2996 5918
rect 2940 5814 2996 5852
rect 1932 5394 1988 5404
rect 2044 5516 2212 5572
rect 8876 5684 8932 5694
rect 4476 5516 4740 5526
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 4788 1764 5070
rect 2044 5010 2100 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2156 5012 2212 5022
rect 1708 4722 1764 4732
rect 2044 4564 2100 4574
rect 2156 4564 2212 4956
rect 2492 4788 2548 5070
rect 2492 4722 2548 4732
rect 2044 4562 2212 4564
rect 2044 4510 2046 4562
rect 2098 4510 2212 4562
rect 2044 4508 2212 4510
rect 8876 4562 8932 5628
rect 10556 5572 10612 5582
rect 10108 5348 10164 5358
rect 8876 4510 8878 4562
rect 8930 4510 8932 4562
rect 2044 4498 2100 4508
rect 8876 4498 8932 4510
rect 9436 4898 9492 4910
rect 9436 4846 9438 4898
rect 9490 4846 9492 4898
rect 1708 4338 1764 4350
rect 1708 4286 1710 4338
rect 1762 4286 1764 4338
rect 1708 4116 1764 4286
rect 9436 4340 9492 4846
rect 9996 4564 10052 4574
rect 10108 4564 10164 5292
rect 9996 4562 10164 4564
rect 9996 4510 9998 4562
rect 10050 4510 10164 4562
rect 9996 4508 10164 4510
rect 9996 4498 10052 4508
rect 10332 4452 10388 4462
rect 10108 4450 10388 4452
rect 10108 4398 10334 4450
rect 10386 4398 10388 4450
rect 10108 4396 10388 4398
rect 9660 4340 9716 4350
rect 9436 4338 9716 4340
rect 9436 4286 9662 4338
rect 9714 4286 9716 4338
rect 9436 4284 9716 4286
rect 1708 4050 1764 4060
rect 2044 4228 2100 4238
rect 1708 3444 1764 3454
rect 1708 3350 1764 3388
rect 2044 3442 2100 4172
rect 2492 4226 2548 4238
rect 2492 4174 2494 4226
rect 2546 4174 2548 4226
rect 2492 4116 2548 4174
rect 8092 4116 8148 4126
rect 2492 4050 2548 4060
rect 7756 4114 8148 4116
rect 7756 4062 8094 4114
rect 8146 4062 8148 4114
rect 7756 4060 8148 4062
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 7196 3780 7252 3790
rect 2044 3390 2046 3442
rect 2098 3390 2100 3442
rect 2044 3378 2100 3390
rect 2940 3444 2996 3454
rect 6860 3444 6916 3454
rect 2940 3350 2996 3388
rect 6748 3442 7140 3444
rect 6748 3390 6862 3442
rect 6914 3390 7140 3442
rect 6748 3388 7140 3390
rect 2380 3330 2436 3342
rect 2380 3278 2382 3330
rect 2434 3278 2436 3330
rect 2380 2772 2436 3278
rect 2380 2706 2436 2716
rect 6748 800 6804 3388
rect 6860 3378 6916 3388
rect 7084 3220 7140 3388
rect 7196 3442 7252 3724
rect 7196 3390 7198 3442
rect 7250 3390 7252 3442
rect 7196 3378 7252 3390
rect 7644 3442 7700 3454
rect 7644 3390 7646 3442
rect 7698 3390 7700 3442
rect 7644 3220 7700 3390
rect 7084 3164 7700 3220
rect 7756 2100 7812 4060
rect 8092 4050 8148 4060
rect 8764 3556 8820 3566
rect 8764 3462 8820 3500
rect 7980 3332 8036 3342
rect 7980 3330 8148 3332
rect 7980 3278 7982 3330
rect 8034 3278 8148 3330
rect 7980 3276 8148 3278
rect 7980 3266 8036 3276
rect 7420 2044 7812 2100
rect 7420 800 7476 2044
rect 8092 800 8148 3276
rect 9660 3108 9716 4284
rect 9436 3052 9716 3108
rect 9772 3330 9828 3342
rect 9772 3278 9774 3330
rect 9826 3278 9828 3330
rect 8876 980 8932 990
rect 8764 978 8932 980
rect 8764 926 8878 978
rect 8930 926 8932 978
rect 8764 924 8932 926
rect 8764 800 8820 924
rect 8876 914 8932 924
rect 9436 800 9492 3052
rect 9772 978 9828 3278
rect 9772 926 9774 978
rect 9826 926 9828 978
rect 9772 914 9828 926
rect 10108 800 10164 4396
rect 10332 4386 10388 4396
rect 10556 3554 10612 5516
rect 12572 5236 12628 5246
rect 12460 5180 12572 5236
rect 11788 5012 11844 5022
rect 12236 5012 12292 5022
rect 11452 4226 11508 4238
rect 11452 4174 11454 4226
rect 11506 4174 11508 4226
rect 11452 3892 11508 4174
rect 10556 3502 10558 3554
rect 10610 3502 10612 3554
rect 10556 3490 10612 3502
rect 10892 3836 11508 3892
rect 11564 4114 11620 4126
rect 11564 4062 11566 4114
rect 11618 4062 11620 4114
rect 10892 3444 10948 3836
rect 11004 3668 11060 3678
rect 11060 3612 11284 3668
rect 11004 3602 11060 3612
rect 10780 3442 10948 3444
rect 10780 3390 10894 3442
rect 10946 3390 10948 3442
rect 10780 3388 10948 3390
rect 10780 800 10836 3388
rect 10892 3378 10948 3388
rect 11228 3330 11284 3612
rect 11564 3444 11620 4062
rect 11228 3278 11230 3330
rect 11282 3278 11284 3330
rect 11228 3266 11284 3278
rect 11452 3442 11620 3444
rect 11452 3390 11566 3442
rect 11618 3390 11620 3442
rect 11452 3388 11620 3390
rect 11788 3444 11844 4956
rect 11900 5010 12292 5012
rect 11900 4958 12238 5010
rect 12290 4958 12292 5010
rect 11900 4956 12292 4958
rect 11900 3780 11956 4956
rect 12236 4946 12292 4956
rect 12012 4226 12068 4238
rect 12012 4174 12014 4226
rect 12066 4174 12068 4226
rect 12012 4114 12068 4174
rect 12348 4116 12404 4126
rect 12012 4062 12014 4114
rect 12066 4062 12068 4114
rect 12012 4050 12068 4062
rect 12124 4114 12404 4116
rect 12124 4062 12350 4114
rect 12402 4062 12404 4114
rect 12124 4060 12404 4062
rect 11900 3714 11956 3724
rect 11788 3388 11956 3444
rect 11452 800 11508 3388
rect 11564 3378 11620 3388
rect 11900 3330 11956 3388
rect 11900 3278 11902 3330
rect 11954 3278 11956 3330
rect 11900 3266 11956 3278
rect 12124 800 12180 4060
rect 12348 4050 12404 4060
rect 12236 3556 12292 3566
rect 12236 3462 12292 3500
rect 12460 3444 12516 5180
rect 12572 5170 12628 5180
rect 14700 5236 14756 5246
rect 13692 5124 13748 5134
rect 13692 5030 13748 5068
rect 14700 5122 14756 5180
rect 14700 5070 14702 5122
rect 14754 5070 14756 5122
rect 14700 5058 14756 5070
rect 14812 5124 14868 5134
rect 12572 4900 12628 4910
rect 13468 4900 13524 4910
rect 12572 4898 13076 4900
rect 12572 4846 12574 4898
rect 12626 4846 13076 4898
rect 12572 4844 13076 4846
rect 12572 4834 12628 4844
rect 13020 4338 13076 4844
rect 13468 4898 13860 4900
rect 13468 4846 13470 4898
rect 13522 4846 13860 4898
rect 13468 4844 13860 4846
rect 13468 4834 13524 4844
rect 13020 4286 13022 4338
rect 13074 4286 13076 4338
rect 13020 4274 13076 4286
rect 13580 4228 13636 4238
rect 13468 4226 13636 4228
rect 13468 4174 13582 4226
rect 13634 4174 13636 4226
rect 13468 4172 13636 4174
rect 13468 3556 13524 4172
rect 13580 4162 13636 4172
rect 12572 3444 12628 3454
rect 12460 3442 12628 3444
rect 12460 3390 12574 3442
rect 12626 3390 12628 3442
rect 12460 3388 12628 3390
rect 12572 3378 12628 3388
rect 13132 3332 13188 3342
rect 12796 3330 13188 3332
rect 12796 3278 13134 3330
rect 13186 3278 13188 3330
rect 12796 3276 13188 3278
rect 12796 800 12852 3276
rect 13132 3266 13188 3276
rect 13468 800 13524 3500
rect 13804 3554 13860 4844
rect 14700 4564 14756 4574
rect 14812 4564 14868 5068
rect 15596 5124 15652 5134
rect 15596 5030 15652 5068
rect 16380 5124 16436 5134
rect 14700 4562 14868 4564
rect 14700 4510 14702 4562
rect 14754 4510 14868 4562
rect 14700 4508 14868 4510
rect 15036 4898 15092 4910
rect 15036 4846 15038 4898
rect 15090 4846 15092 4898
rect 15036 4562 15092 4846
rect 15932 4900 15988 4910
rect 15932 4898 16324 4900
rect 15932 4846 15934 4898
rect 15986 4846 16324 4898
rect 15932 4844 16324 4846
rect 15932 4834 15988 4844
rect 15036 4510 15038 4562
rect 15090 4510 15092 4562
rect 14700 4498 14756 4508
rect 15036 4498 15092 4510
rect 14364 4338 14420 4350
rect 14364 4286 14366 4338
rect 14418 4286 14420 4338
rect 13804 3502 13806 3554
rect 13858 3502 13860 3554
rect 13804 3490 13860 3502
rect 14140 4228 14196 4238
rect 14364 4228 14420 4286
rect 15484 4228 15540 4238
rect 14140 4226 14420 4228
rect 14140 4174 14142 4226
rect 14194 4174 14420 4226
rect 14140 4172 14420 4174
rect 14812 4226 15540 4228
rect 14812 4174 15486 4226
rect 15538 4174 15540 4226
rect 14812 4172 15540 4174
rect 14140 800 14196 4172
rect 14812 800 14868 4172
rect 15484 4162 15540 4172
rect 16268 3554 16324 4844
rect 16268 3502 16270 3554
rect 16322 3502 16324 3554
rect 16268 3490 16324 3502
rect 16380 3388 16436 5068
rect 16604 5010 16660 6636
rect 18284 5796 18340 5806
rect 16940 5124 16996 5134
rect 17500 5124 17556 5134
rect 16940 5122 17332 5124
rect 16940 5070 16942 5122
rect 16994 5070 17332 5122
rect 16940 5068 17332 5070
rect 16940 5058 16996 5068
rect 16604 4958 16606 5010
rect 16658 4958 16660 5010
rect 16604 4946 16660 4958
rect 17276 5010 17332 5068
rect 17500 5030 17556 5068
rect 18060 5124 18116 5134
rect 18060 5030 18116 5068
rect 17276 4958 17278 5010
rect 17330 4958 17332 5010
rect 17276 4946 17332 4958
rect 17724 4564 17780 4574
rect 17724 4470 17780 4508
rect 17388 4338 17444 4350
rect 17388 4286 17390 4338
rect 17442 4286 17444 4338
rect 15596 3332 15652 3342
rect 15484 3330 15652 3332
rect 15484 3278 15598 3330
rect 15650 3278 15652 3330
rect 15484 3276 15652 3278
rect 15484 800 15540 3276
rect 15596 3266 15652 3276
rect 16156 3332 16436 3388
rect 16828 4228 16884 4238
rect 17388 4228 17444 4286
rect 16828 4226 17444 4228
rect 16828 4174 16830 4226
rect 16882 4174 17444 4226
rect 16828 4172 17444 4174
rect 18284 4228 18340 5740
rect 18396 5010 18452 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 22204 7364 22260 7374
rect 18620 6356 18676 6366
rect 18396 4958 18398 5010
rect 18450 4958 18452 5010
rect 18396 4946 18452 4958
rect 18508 5236 18564 5246
rect 16156 800 16212 3332
rect 16828 800 16884 4172
rect 18284 4162 18340 4172
rect 18396 4450 18452 4462
rect 18396 4398 18398 4450
rect 18450 4398 18452 4450
rect 18396 3388 18452 4398
rect 18508 3554 18564 5180
rect 18620 5122 18676 6300
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 22204 6130 22260 7308
rect 22204 6078 22206 6130
rect 22258 6078 22260 6130
rect 22204 6066 22260 6078
rect 23884 6132 23940 6142
rect 20748 6020 20804 6030
rect 20748 5926 20804 5964
rect 22988 6018 23044 6030
rect 22988 5966 22990 6018
rect 23042 5966 23044 6018
rect 20972 5906 21028 5918
rect 20972 5854 20974 5906
rect 21026 5854 21028 5906
rect 20412 5796 20468 5806
rect 20412 5702 20468 5740
rect 20972 5796 21028 5854
rect 20972 5730 21028 5740
rect 21644 5908 21700 5918
rect 19740 5124 19796 5134
rect 18620 5070 18622 5122
rect 18674 5070 18676 5122
rect 18620 5058 18676 5070
rect 19404 5122 19796 5124
rect 19404 5070 19742 5122
rect 19794 5070 19796 5122
rect 19404 5068 19796 5070
rect 19404 4562 19460 5068
rect 19740 5058 19796 5068
rect 20412 5010 20468 5022
rect 20412 4958 20414 5010
rect 20466 4958 20468 5010
rect 19404 4510 19406 4562
rect 19458 4510 19460 4562
rect 19404 4498 19460 4510
rect 19516 4898 19572 4910
rect 19516 4846 19518 4898
rect 19570 4846 19572 4898
rect 19516 4452 19572 4846
rect 20076 4900 20132 4910
rect 20076 4898 20244 4900
rect 20076 4846 20078 4898
rect 20130 4846 20244 4898
rect 20076 4844 20244 4846
rect 20076 4834 20132 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19740 4452 19796 4462
rect 19516 4450 19796 4452
rect 19516 4398 19742 4450
rect 19794 4398 19796 4450
rect 19516 4396 19796 4398
rect 18508 3502 18510 3554
rect 18562 3502 18564 3554
rect 18508 3490 18564 3502
rect 19068 4338 19124 4350
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 3666 19124 4286
rect 19068 3614 19070 3666
rect 19122 3614 19124 3666
rect 19068 3388 19124 3614
rect 17836 3332 17892 3342
rect 17500 3330 17892 3332
rect 17500 3278 17838 3330
rect 17890 3278 17892 3330
rect 17500 3276 17892 3278
rect 17500 800 17556 3276
rect 17836 3266 17892 3276
rect 18172 3332 18452 3388
rect 18844 3332 19124 3388
rect 18172 800 18228 3332
rect 18844 800 18900 3332
rect 19516 800 19572 4396
rect 19740 4386 19796 4396
rect 20076 4452 20132 4490
rect 20076 4386 20132 4396
rect 19740 3666 19796 3678
rect 19740 3614 19742 3666
rect 19794 3614 19796 3666
rect 19740 3388 19796 3614
rect 20188 3554 20244 4844
rect 20412 4452 20468 4958
rect 20748 4898 20804 4910
rect 20748 4846 20750 4898
rect 20802 4846 20804 4898
rect 20748 4564 20804 4846
rect 21084 4564 21140 4574
rect 20748 4562 21140 4564
rect 20748 4510 21086 4562
rect 21138 4510 21140 4562
rect 20748 4508 21140 4510
rect 21084 4498 21140 4508
rect 20412 4386 20468 4396
rect 21532 4228 21588 4238
rect 21308 4226 21588 4228
rect 21308 4174 21534 4226
rect 21586 4174 21588 4226
rect 21308 4172 21588 4174
rect 20188 3502 20190 3554
rect 20242 3502 20244 3554
rect 20188 3490 20244 3502
rect 21196 3554 21252 3566
rect 21196 3502 21198 3554
rect 21250 3502 21252 3554
rect 21196 3444 21252 3502
rect 19740 3332 20244 3388
rect 21196 3378 21252 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3332
rect 21308 1764 21364 4172
rect 21532 4162 21588 4172
rect 21420 3444 21476 3454
rect 21644 3444 21700 5852
rect 22428 5908 22484 5918
rect 22428 5814 22484 5852
rect 22204 5572 22260 5582
rect 21756 5012 21812 5022
rect 22204 5012 22260 5516
rect 22988 5236 23044 5966
rect 23660 6018 23716 6030
rect 23660 5966 23662 6018
rect 23714 5966 23716 6018
rect 23212 5906 23268 5918
rect 23212 5854 23214 5906
rect 23266 5854 23268 5906
rect 22988 5170 23044 5180
rect 23100 5348 23156 5358
rect 22764 5124 22820 5134
rect 22764 5030 22820 5068
rect 23100 5122 23156 5292
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 23100 5058 23156 5070
rect 22428 5012 22484 5022
rect 22204 5010 22484 5012
rect 22204 4958 22430 5010
rect 22482 4958 22484 5010
rect 22204 4956 22484 4958
rect 21756 4918 21812 4956
rect 22428 4946 22484 4956
rect 22652 5012 22708 5022
rect 22092 4898 22148 4910
rect 22092 4846 22094 4898
rect 22146 4846 22148 4898
rect 22092 4452 22148 4846
rect 22652 4562 22708 4956
rect 22652 4510 22654 4562
rect 22706 4510 22708 4562
rect 22652 4498 22708 4510
rect 23212 4564 23268 5854
rect 23660 5684 23716 5966
rect 23660 5618 23716 5628
rect 23436 5124 23492 5134
rect 23436 5010 23492 5068
rect 23884 5122 23940 6076
rect 23884 5070 23886 5122
rect 23938 5070 23940 5122
rect 23884 5058 23940 5070
rect 23996 5906 24052 5918
rect 23996 5854 23998 5906
rect 24050 5854 24052 5906
rect 23436 4958 23438 5010
rect 23490 4958 23492 5010
rect 23436 4946 23492 4958
rect 23212 4498 23268 4508
rect 22092 4396 22484 4452
rect 22316 4226 22372 4238
rect 22316 4174 22318 4226
rect 22370 4174 22372 4226
rect 21420 3442 21700 3444
rect 21420 3390 21422 3442
rect 21474 3390 21700 3442
rect 21420 3388 21700 3390
rect 22092 3444 22148 3454
rect 22316 3388 22372 4174
rect 22428 3554 22484 4396
rect 23324 4450 23380 4462
rect 23324 4398 23326 4450
rect 23378 4398 23380 4450
rect 22428 3502 22430 3554
rect 22482 3502 22484 3554
rect 22428 3490 22484 3502
rect 22876 4338 22932 4350
rect 22876 4286 22878 4338
rect 22930 4286 22932 4338
rect 22876 3668 22932 4286
rect 23212 3668 23268 3678
rect 22876 3666 23268 3668
rect 22876 3614 23214 3666
rect 23266 3614 23268 3666
rect 22876 3612 23268 3614
rect 21420 3378 21476 3388
rect 21756 3332 21812 3342
rect 22092 3332 22372 3388
rect 20860 1708 21364 1764
rect 21532 3330 21812 3332
rect 21532 3278 21758 3330
rect 21810 3278 21812 3330
rect 21532 3276 21812 3278
rect 20860 800 20916 1708
rect 21532 800 21588 3276
rect 21756 3266 21812 3276
rect 22204 800 22260 3332
rect 22876 800 22932 3612
rect 23212 3602 23268 3612
rect 23324 3556 23380 4398
rect 23548 4338 23604 4350
rect 23548 4286 23550 4338
rect 23602 4286 23604 4338
rect 23548 3668 23604 4286
rect 23548 3602 23604 3612
rect 23324 3490 23380 3500
rect 23660 3442 23716 3454
rect 23660 3390 23662 3442
rect 23714 3390 23716 3442
rect 23660 3388 23716 3390
rect 23996 3442 24052 5854
rect 24108 5010 24164 9996
rect 25228 8036 25284 8046
rect 24444 6132 24500 6142
rect 24444 6038 24500 6076
rect 25228 6132 25284 7980
rect 25228 6066 25284 6076
rect 26460 6018 26516 6030
rect 26460 5966 26462 6018
rect 26514 5966 26516 6018
rect 26236 5906 26292 5918
rect 26236 5854 26238 5906
rect 26290 5854 26292 5906
rect 24892 5236 24948 5246
rect 24780 5234 24948 5236
rect 24780 5182 24894 5234
rect 24946 5182 24948 5234
rect 24780 5180 24948 5182
rect 24444 5124 24500 5134
rect 24444 5030 24500 5068
rect 24108 4958 24110 5010
rect 24162 4958 24164 5010
rect 24108 4946 24164 4958
rect 24444 4450 24500 4462
rect 24444 4398 24446 4450
rect 24498 4398 24500 4450
rect 24220 4340 24276 4350
rect 24220 4246 24276 4284
rect 24444 3556 24500 4398
rect 24444 3490 24500 3500
rect 23996 3390 23998 3442
rect 24050 3390 24052 3442
rect 23548 3332 23940 3388
rect 23996 3378 24052 3390
rect 24668 3442 24724 3454
rect 24668 3390 24670 3442
rect 24722 3390 24724 3442
rect 24668 3388 24724 3390
rect 23548 800 23604 3332
rect 23884 3220 23940 3332
rect 24108 3332 24724 3388
rect 24108 3220 24164 3332
rect 23884 3164 24164 3220
rect 24780 1764 24836 5180
rect 24892 5170 24948 5180
rect 26124 5122 26180 5134
rect 26124 5070 26126 5122
rect 26178 5070 26180 5122
rect 26124 4004 26180 5070
rect 26236 4564 26292 5854
rect 26348 4898 26404 4910
rect 26348 4846 26350 4898
rect 26402 4846 26404 4898
rect 26348 4564 26404 4846
rect 26460 4788 26516 5966
rect 28252 5796 28308 5806
rect 27020 5684 27076 5694
rect 26460 4722 26516 4732
rect 26684 5010 26740 5022
rect 26684 4958 26686 5010
rect 26738 4958 26740 5010
rect 26460 4564 26516 4574
rect 26348 4562 26516 4564
rect 26348 4510 26462 4562
rect 26514 4510 26516 4562
rect 26348 4508 26516 4510
rect 26236 4498 26292 4508
rect 26460 4498 26516 4508
rect 26684 4340 26740 4958
rect 27020 5010 27076 5628
rect 28252 5122 28308 5740
rect 28252 5070 28254 5122
rect 28306 5070 28308 5122
rect 28252 5058 28308 5070
rect 27020 4958 27022 5010
rect 27074 4958 27076 5010
rect 27020 4946 27076 4958
rect 28476 5010 28532 12684
rect 28588 12628 28644 12638
rect 28588 10052 28644 12572
rect 28812 11396 28868 15820
rect 28924 15316 28980 16044
rect 29036 16034 29092 16044
rect 28924 15222 28980 15260
rect 29260 15314 29316 15326
rect 29260 15262 29262 15314
rect 29314 15262 29316 15314
rect 29260 11732 29316 15262
rect 29372 13860 29428 17164
rect 29484 16882 29540 16894
rect 29484 16830 29486 16882
rect 29538 16830 29540 16882
rect 29484 14196 29540 16830
rect 29596 16884 29652 17612
rect 29596 16818 29652 16828
rect 29708 16100 29764 16110
rect 29708 16098 29876 16100
rect 29708 16046 29710 16098
rect 29762 16046 29876 16098
rect 29708 16044 29876 16046
rect 29708 16034 29764 16044
rect 29708 15316 29764 15326
rect 29708 14530 29764 15260
rect 29708 14478 29710 14530
rect 29762 14478 29764 14530
rect 29708 14466 29764 14478
rect 29484 14140 29652 14196
rect 29484 13860 29540 13870
rect 29372 13858 29540 13860
rect 29372 13806 29486 13858
rect 29538 13806 29540 13858
rect 29372 13804 29540 13806
rect 29484 13794 29540 13804
rect 29372 12068 29428 12078
rect 29372 11974 29428 12012
rect 29260 11666 29316 11676
rect 29596 11508 29652 14140
rect 29820 13636 29876 16044
rect 29820 13570 29876 13580
rect 30044 13076 30100 19404
rect 30268 18450 30324 20860
rect 31276 20916 31332 21534
rect 33180 21586 33236 22316
rect 33180 21534 33182 21586
rect 33234 21534 33236 21586
rect 33180 21522 33236 21534
rect 31276 20850 31332 20860
rect 32172 20578 32228 20590
rect 32172 20526 32174 20578
rect 32226 20526 32228 20578
rect 32060 20132 32116 20142
rect 32060 20038 32116 20076
rect 31052 19908 31108 19918
rect 31052 19814 31108 19852
rect 31052 19348 31108 19358
rect 30268 18398 30270 18450
rect 30322 18398 30324 18450
rect 30268 18386 30324 18398
rect 30604 18564 30660 18574
rect 30268 17780 30324 17790
rect 30268 17686 30324 17724
rect 30492 17666 30548 17678
rect 30492 17614 30494 17666
rect 30546 17614 30548 17666
rect 30156 17442 30212 17454
rect 30156 17390 30158 17442
rect 30210 17390 30212 17442
rect 30156 15540 30212 17390
rect 30492 16884 30548 17614
rect 30492 16818 30548 16828
rect 30156 15474 30212 15484
rect 30380 14530 30436 14542
rect 30380 14478 30382 14530
rect 30434 14478 30436 14530
rect 30380 13188 30436 14478
rect 30604 13634 30660 18508
rect 31052 18562 31108 19292
rect 31948 19348 32004 19358
rect 31052 18510 31054 18562
rect 31106 18510 31108 18562
rect 31052 18498 31108 18510
rect 31276 18676 31332 18686
rect 31164 17666 31220 17678
rect 31164 17614 31166 17666
rect 31218 17614 31220 17666
rect 31164 14756 31220 17614
rect 31164 14690 31220 14700
rect 30604 13582 30606 13634
rect 30658 13582 30660 13634
rect 30604 13570 30660 13582
rect 30380 13122 30436 13132
rect 30268 13076 30324 13086
rect 30044 13074 30324 13076
rect 30044 13022 30270 13074
rect 30322 13022 30324 13074
rect 30044 13020 30324 13022
rect 30268 13010 30324 13020
rect 31276 12850 31332 18620
rect 31724 18452 31780 18462
rect 31724 18358 31780 18396
rect 31948 18450 32004 19292
rect 32172 18900 32228 20526
rect 32732 20578 32788 20590
rect 32732 20526 32734 20578
rect 32786 20526 32788 20578
rect 32508 19236 32564 19246
rect 32284 19012 32340 19022
rect 32284 18918 32340 18956
rect 32172 18834 32228 18844
rect 31948 18398 31950 18450
rect 32002 18398 32004 18450
rect 31388 18340 31444 18350
rect 31388 18246 31444 18284
rect 31948 18340 32004 18398
rect 31948 18274 32004 18284
rect 32508 18674 32564 19180
rect 32732 19124 32788 20526
rect 33068 20020 33124 20030
rect 33068 19926 33124 19964
rect 33292 20020 33348 23100
rect 33516 22372 33572 22382
rect 33404 22370 33572 22372
rect 33404 22318 33518 22370
rect 33570 22318 33572 22370
rect 33404 22316 33572 22318
rect 33404 20188 33460 22316
rect 33516 22306 33572 22316
rect 33628 21588 33684 21598
rect 33964 21588 34020 21598
rect 33628 21586 33908 21588
rect 33628 21534 33630 21586
rect 33682 21534 33908 21586
rect 33628 21532 33908 21534
rect 33628 21522 33684 21532
rect 33628 20578 33684 20590
rect 33628 20526 33630 20578
rect 33682 20526 33684 20578
rect 33404 20132 33572 20188
rect 33292 19348 33348 19964
rect 33516 19460 33572 20132
rect 33292 19282 33348 19292
rect 33404 19404 33572 19460
rect 33628 20132 33684 20526
rect 32732 19058 32788 19068
rect 32844 19012 32900 19022
rect 32844 19010 33348 19012
rect 32844 18958 32846 19010
rect 32898 18958 33348 19010
rect 32844 18956 33348 18958
rect 32844 18946 32900 18956
rect 32508 18622 32510 18674
rect 32562 18622 32564 18674
rect 32508 18228 32564 18622
rect 32508 18162 32564 18172
rect 33180 18450 33236 18462
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 31724 17332 31780 17342
rect 31612 15540 31668 15550
rect 31612 15446 31668 15484
rect 31276 12798 31278 12850
rect 31330 12798 31332 12850
rect 31276 12786 31332 12798
rect 30380 12292 30436 12302
rect 30380 12198 30436 12236
rect 29596 11442 29652 11452
rect 30492 11508 30548 11518
rect 30492 11414 30548 11452
rect 28812 11340 29428 11396
rect 29372 11282 29428 11340
rect 29372 11230 29374 11282
rect 29426 11230 29428 11282
rect 29372 11218 29428 11230
rect 28588 9986 28644 9996
rect 31724 8372 31780 17276
rect 31836 16994 31892 17006
rect 31836 16942 31838 16994
rect 31890 16942 31892 16994
rect 31836 15316 31892 16942
rect 33180 16884 33236 18398
rect 32620 16658 32676 16670
rect 32620 16606 32622 16658
rect 32674 16606 32676 16658
rect 32172 15874 32228 15886
rect 32172 15822 32174 15874
rect 32226 15822 32228 15874
rect 31836 15260 32004 15316
rect 31948 13860 32004 15260
rect 32172 14644 32228 15822
rect 32396 15092 32452 15102
rect 32396 14998 32452 15036
rect 32172 14578 32228 14588
rect 32396 14756 32452 14766
rect 32172 13860 32228 13870
rect 31948 13858 32228 13860
rect 31948 13806 32174 13858
rect 32226 13806 32228 13858
rect 31948 13804 32228 13806
rect 32172 13794 32228 13804
rect 32396 11620 32452 14700
rect 32508 13860 32564 13870
rect 32508 13766 32564 13804
rect 32620 13412 32676 16606
rect 33068 16100 33124 16110
rect 33180 16100 33236 16828
rect 33068 16098 33236 16100
rect 33068 16046 33070 16098
rect 33122 16046 33236 16098
rect 33068 16044 33236 16046
rect 33068 16034 33124 16044
rect 32732 15874 32788 15886
rect 32732 15822 32734 15874
rect 32786 15822 32788 15874
rect 32732 14980 32788 15822
rect 32732 14914 32788 14924
rect 32956 15090 33012 15102
rect 32956 15038 32958 15090
rect 33010 15038 33012 15090
rect 32844 14308 32900 14318
rect 32844 14214 32900 14252
rect 32620 13346 32676 13356
rect 32396 11554 32452 11564
rect 32732 13188 32788 13198
rect 32732 9938 32788 13132
rect 32956 10724 33012 15038
rect 33292 14756 33348 18956
rect 33404 14868 33460 19404
rect 33516 19236 33572 19246
rect 33628 19236 33684 20076
rect 33740 19908 33796 19918
rect 33740 19814 33796 19852
rect 33572 19180 33684 19236
rect 33516 19142 33572 19180
rect 33852 18564 33908 21532
rect 33964 20914 34020 21532
rect 33964 20862 33966 20914
rect 34018 20862 34020 20914
rect 33964 20850 34020 20862
rect 34076 20188 34132 27020
rect 35532 26964 35588 26974
rect 35532 26870 35588 26908
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35644 25844 35700 27132
rect 35196 25834 35460 25844
rect 35532 25788 35700 25844
rect 35308 25732 35364 25742
rect 35532 25732 35588 25788
rect 35308 25730 35588 25732
rect 35308 25678 35310 25730
rect 35362 25678 35588 25730
rect 35308 25676 35588 25678
rect 35308 25666 35364 25676
rect 34300 25508 34356 25518
rect 34300 20188 34356 25452
rect 34748 25282 34804 25294
rect 34748 25230 34750 25282
rect 34802 25230 34804 25282
rect 34748 23380 34804 25230
rect 35756 25282 35812 27916
rect 36540 27906 36596 27916
rect 36764 27748 36820 33404
rect 36540 27692 36820 27748
rect 36876 33236 36932 33246
rect 36428 26964 36484 26974
rect 36428 26870 36484 26908
rect 36092 26292 36148 26302
rect 36540 26292 36596 27692
rect 36764 26516 36820 26526
rect 36876 26516 36932 33180
rect 37100 31556 37156 31566
rect 36988 31554 37156 31556
rect 36988 31502 37102 31554
rect 37154 31502 37156 31554
rect 36988 31500 37156 31502
rect 36988 30882 37044 31500
rect 37100 31490 37156 31500
rect 36988 30830 36990 30882
rect 37042 30830 37044 30882
rect 36988 30212 37044 30830
rect 36988 30146 37044 30156
rect 36764 26514 36932 26516
rect 36764 26462 36766 26514
rect 36818 26462 36932 26514
rect 36764 26460 36932 26462
rect 36988 28644 37044 28654
rect 36988 27074 37044 28588
rect 36988 27022 36990 27074
rect 37042 27022 37044 27074
rect 36764 26450 36820 26460
rect 36092 26290 36596 26292
rect 36092 26238 36094 26290
rect 36146 26238 36596 26290
rect 36092 26236 36596 26238
rect 36652 26290 36708 26302
rect 36652 26238 36654 26290
rect 36706 26238 36708 26290
rect 36092 26226 36148 26236
rect 35756 25230 35758 25282
rect 35810 25230 35812 25282
rect 35756 25218 35812 25230
rect 35868 25394 35924 25406
rect 35868 25342 35870 25394
rect 35922 25342 35924 25394
rect 35868 25172 35924 25342
rect 36652 25284 36708 26238
rect 36652 25218 36708 25228
rect 35868 25106 35924 25116
rect 36876 25172 36932 25182
rect 35980 24946 36036 24958
rect 35980 24894 35982 24946
rect 36034 24894 36036 24946
rect 35532 24500 35588 24510
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34748 23314 34804 23324
rect 34972 24164 35028 24174
rect 34412 23154 34468 23166
rect 34412 23102 34414 23154
rect 34466 23102 34468 23154
rect 34412 22372 34468 23102
rect 34412 22306 34468 22316
rect 34860 23154 34916 23166
rect 34860 23102 34862 23154
rect 34914 23102 34916 23154
rect 34860 21924 34916 23102
rect 34972 23044 35028 24108
rect 35420 23940 35476 23950
rect 35532 23940 35588 24444
rect 35476 23884 35588 23940
rect 35420 23846 35476 23884
rect 34972 22978 35028 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34860 21858 34916 21868
rect 35756 22146 35812 22158
rect 35756 22094 35758 22146
rect 35810 22094 35812 22146
rect 34972 21700 35028 21710
rect 34972 20690 35028 21644
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34972 20638 34974 20690
rect 35026 20638 35028 20690
rect 34972 20626 35028 20638
rect 34076 20132 34244 20188
rect 34300 20132 34804 20188
rect 34076 20066 34132 20076
rect 33964 20020 34020 20030
rect 34188 20020 34244 20132
rect 34636 20020 34692 20030
rect 34188 20018 34692 20020
rect 34188 19966 34638 20018
rect 34690 19966 34692 20018
rect 34188 19964 34692 19966
rect 33964 19926 34020 19964
rect 34636 19954 34692 19964
rect 34636 19348 34692 19358
rect 33852 18498 33908 18508
rect 34076 19010 34132 19022
rect 34076 18958 34078 19010
rect 34130 18958 34132 19010
rect 33628 18450 33684 18462
rect 33628 18398 33630 18450
rect 33682 18398 33684 18450
rect 33628 17780 33684 18398
rect 34076 17780 34132 18958
rect 33628 17724 33908 17780
rect 33628 17556 33684 17566
rect 33628 17442 33684 17500
rect 33628 17390 33630 17442
rect 33682 17390 33684 17442
rect 33628 17378 33684 17390
rect 33628 16882 33684 16894
rect 33628 16830 33630 16882
rect 33682 16830 33684 16882
rect 33516 16098 33572 16110
rect 33516 16046 33518 16098
rect 33570 16046 33572 16098
rect 33516 15204 33572 16046
rect 33516 15138 33572 15148
rect 33404 14802 33460 14812
rect 33292 14690 33348 14700
rect 33068 14644 33124 14654
rect 33068 13858 33124 14588
rect 33404 14308 33460 14318
rect 33404 14306 33572 14308
rect 33404 14254 33406 14306
rect 33458 14254 33572 14306
rect 33404 14252 33572 14254
rect 33404 14242 33460 14252
rect 33068 13806 33070 13858
rect 33122 13806 33124 13858
rect 33068 13794 33124 13806
rect 33404 13860 33460 13870
rect 33404 13766 33460 13804
rect 33292 13636 33348 13646
rect 33292 13074 33348 13580
rect 33292 13022 33294 13074
rect 33346 13022 33348 13074
rect 33292 13010 33348 13022
rect 33404 11508 33460 11518
rect 33404 11414 33460 11452
rect 32956 10658 33012 10668
rect 32732 9886 32734 9938
rect 32786 9886 32788 9938
rect 32732 9874 32788 9886
rect 33404 9828 33460 9838
rect 31724 8306 31780 8316
rect 32844 8372 32900 8382
rect 30268 7924 30324 7934
rect 28812 5796 28868 5806
rect 28812 5702 28868 5740
rect 28476 4958 28478 5010
rect 28530 4958 28532 5010
rect 28476 4946 28532 4958
rect 29372 5122 29428 5134
rect 29372 5070 29374 5122
rect 29426 5070 29428 5122
rect 28588 4788 28644 4798
rect 28028 4564 28084 4574
rect 28028 4470 28084 4508
rect 26684 4284 27412 4340
rect 26236 4228 26292 4238
rect 26236 4134 26292 4172
rect 27132 4116 27188 4126
rect 26124 3948 26740 4004
rect 25564 3668 25620 3678
rect 25228 3666 25620 3668
rect 25228 3614 25566 3666
rect 25618 3614 25620 3666
rect 25228 3612 25620 3614
rect 25116 3556 25172 3566
rect 25116 3462 25172 3500
rect 25228 3388 25284 3612
rect 25564 3602 25620 3612
rect 25676 3556 25732 3566
rect 25676 3388 25732 3500
rect 26460 3556 26516 3566
rect 26460 3462 26516 3500
rect 24220 1708 24836 1764
rect 24892 3332 25284 3388
rect 25564 3332 25732 3388
rect 26236 3444 26292 3454
rect 24220 800 24276 1708
rect 24892 800 24948 3332
rect 25564 800 25620 3332
rect 26236 800 26292 3388
rect 26684 3442 26740 3948
rect 26908 3556 26964 3566
rect 26908 3462 26964 3500
rect 27132 3556 27188 4060
rect 26684 3390 26686 3442
rect 26738 3390 26740 3442
rect 26684 3378 26740 3390
rect 27132 3388 27188 3500
rect 26908 3332 27188 3388
rect 27244 4114 27300 4126
rect 27244 4062 27246 4114
rect 27298 4062 27300 4114
rect 27244 3444 27300 4062
rect 27244 3378 27300 3388
rect 27356 3442 27412 4284
rect 28252 4338 28308 4350
rect 28252 4286 28254 4338
rect 28306 4286 28308 4338
rect 27692 4228 27748 4238
rect 28252 4228 28308 4286
rect 27356 3390 27358 3442
rect 27410 3390 27412 3442
rect 27356 3378 27412 3390
rect 27580 4226 28308 4228
rect 27580 4174 27694 4226
rect 27746 4174 28308 4226
rect 27580 4172 28308 4174
rect 26908 800 26964 3332
rect 27580 800 27636 4172
rect 27692 4162 27748 4172
rect 27692 3556 27748 3566
rect 27692 3462 27748 3500
rect 28588 3554 28644 4732
rect 29148 4452 29204 4462
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 28924 4450 29204 4452
rect 28924 4398 29150 4450
rect 29202 4398 29204 4450
rect 28924 4396 29204 4398
rect 28252 3444 28308 3454
rect 28252 800 28308 3388
rect 28924 800 28980 4396
rect 29148 4386 29204 4396
rect 29372 4452 29428 5070
rect 30044 5124 30100 5134
rect 30044 5122 30212 5124
rect 30044 5070 30046 5122
rect 30098 5070 30212 5122
rect 30044 5068 30212 5070
rect 30044 5058 30100 5068
rect 29596 4900 29652 4910
rect 29596 4898 29876 4900
rect 29596 4846 29598 4898
rect 29650 4846 29876 4898
rect 29596 4844 29876 4846
rect 29596 4834 29652 4844
rect 29372 4386 29428 4396
rect 29820 4116 29876 4844
rect 30156 4676 30212 5068
rect 30268 5010 30324 7868
rect 31276 7028 31332 7038
rect 31276 5122 31332 6972
rect 32620 6132 32676 6142
rect 31276 5070 31278 5122
rect 31330 5070 31332 5122
rect 31276 5058 31332 5070
rect 31948 5122 32004 5134
rect 31948 5070 31950 5122
rect 32002 5070 32004 5122
rect 30268 4958 30270 5010
rect 30322 4958 30324 5010
rect 30268 4946 30324 4958
rect 30940 4898 30996 4910
rect 30940 4846 30942 4898
rect 30994 4846 30996 4898
rect 30156 4620 30548 4676
rect 30492 4562 30548 4620
rect 30492 4510 30494 4562
rect 30546 4510 30548 4562
rect 30492 4498 30548 4510
rect 30716 4338 30772 4350
rect 30716 4286 30718 4338
rect 30770 4286 30772 4338
rect 30268 4228 30324 4238
rect 30716 4228 30772 4286
rect 30268 4226 30772 4228
rect 30268 4174 30270 4226
rect 30322 4174 30772 4226
rect 30268 4172 30772 4174
rect 29820 4060 30100 4116
rect 29596 3668 29652 3678
rect 29260 3444 29316 3454
rect 29260 3350 29316 3388
rect 29596 800 29652 3612
rect 30044 3554 30100 4060
rect 30044 3502 30046 3554
rect 30098 3502 30100 3554
rect 30044 3490 30100 3502
rect 30268 800 30324 4172
rect 30940 4004 30996 4846
rect 31500 4900 31556 4910
rect 31500 4806 31556 4844
rect 31948 4564 32004 5070
rect 32620 5122 32676 6076
rect 32620 5070 32622 5122
rect 32674 5070 32676 5122
rect 32620 5058 32676 5070
rect 32844 5010 32900 8316
rect 33404 6130 33460 9772
rect 33516 9156 33572 14252
rect 33628 10500 33684 16830
rect 33740 15426 33796 15438
rect 33740 15374 33742 15426
rect 33794 15374 33796 15426
rect 33740 14644 33796 15374
rect 33740 14578 33796 14588
rect 33740 14308 33796 14318
rect 33740 13858 33796 14252
rect 33740 13806 33742 13858
rect 33794 13806 33796 13858
rect 33740 13794 33796 13806
rect 33852 12068 33908 17724
rect 33852 12002 33908 12012
rect 33964 14980 34020 14990
rect 33852 10836 33908 10846
rect 33740 10500 33796 10510
rect 33628 10444 33740 10500
rect 33740 10434 33796 10444
rect 33516 9090 33572 9100
rect 33628 9044 33684 9054
rect 33628 7028 33684 8988
rect 33628 6962 33684 6972
rect 33404 6078 33406 6130
rect 33458 6078 33460 6130
rect 33404 6066 33460 6078
rect 33852 6132 33908 10780
rect 33964 9714 34020 14924
rect 34076 13860 34132 17724
rect 34412 18900 34468 18910
rect 34412 17778 34468 18844
rect 34412 17726 34414 17778
rect 34466 17726 34468 17778
rect 34412 17714 34468 17726
rect 34636 17666 34692 19292
rect 34636 17614 34638 17666
rect 34690 17614 34692 17666
rect 34636 17602 34692 17614
rect 34188 17442 34244 17454
rect 34188 17390 34190 17442
rect 34242 17390 34244 17442
rect 34188 16772 34244 17390
rect 34188 16706 34244 16716
rect 34748 16660 34804 20132
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35644 18564 35700 18574
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35308 17780 35364 17790
rect 35308 17666 35364 17724
rect 35308 17614 35310 17666
rect 35362 17614 35364 17666
rect 35308 17602 35364 17614
rect 35084 17556 35140 17566
rect 35084 17462 35140 17500
rect 35644 16996 35700 18508
rect 35756 17778 35812 22094
rect 35868 21698 35924 21710
rect 35868 21646 35870 21698
rect 35922 21646 35924 21698
rect 35868 20132 35924 21646
rect 35980 20578 36036 24894
rect 36652 24498 36708 24510
rect 36652 24446 36654 24498
rect 36706 24446 36708 24498
rect 36204 24052 36260 24062
rect 36204 23958 36260 23996
rect 36652 22260 36708 24446
rect 36876 24052 36932 25116
rect 36988 24836 37044 27022
rect 37212 27076 37268 34972
rect 37324 34242 37380 34254
rect 37324 34190 37326 34242
rect 37378 34190 37380 34242
rect 37324 31108 37380 34190
rect 37436 31220 37492 36318
rect 38108 36260 38164 37326
rect 38108 36194 38164 36204
rect 37772 35588 37828 35598
rect 37436 31154 37492 31164
rect 37660 32450 37716 32462
rect 37660 32398 37662 32450
rect 37714 32398 37716 32450
rect 37324 31042 37380 31052
rect 37436 30884 37492 30894
rect 37324 30882 37492 30884
rect 37324 30830 37438 30882
rect 37490 30830 37492 30882
rect 37324 30828 37492 30830
rect 37324 30212 37380 30828
rect 37436 30818 37492 30828
rect 37324 28644 37380 30156
rect 37548 30324 37604 30334
rect 37324 28578 37380 28588
rect 37436 28868 37492 28878
rect 37324 28084 37380 28094
rect 37436 28084 37492 28812
rect 37548 28642 37604 30268
rect 37660 28756 37716 32398
rect 37772 30210 37828 35532
rect 38108 35026 38164 35038
rect 38108 34974 38110 35026
rect 38162 34974 38164 35026
rect 37996 33460 38052 33470
rect 37996 33366 38052 33404
rect 38108 30996 38164 34974
rect 38444 31948 38500 39676
rect 38556 39666 38612 39676
rect 43036 39732 43092 39742
rect 43036 39638 43092 39676
rect 42252 39506 42308 39518
rect 42252 39454 42254 39506
rect 42306 39454 42308 39506
rect 40236 38724 40292 38734
rect 39452 38164 39508 38174
rect 39228 37154 39284 37166
rect 39228 37102 39230 37154
rect 39282 37102 39284 37154
rect 38556 36596 38612 36606
rect 38556 36594 38724 36596
rect 38556 36542 38558 36594
rect 38610 36542 38724 36594
rect 38556 36540 38724 36542
rect 38556 36530 38612 36540
rect 38668 36484 38724 36540
rect 38668 36428 38836 36484
rect 38780 34132 38836 36428
rect 39116 35812 39172 35822
rect 38892 35588 38948 35598
rect 38892 35494 38948 35532
rect 38780 34066 38836 34076
rect 39004 34802 39060 34814
rect 39004 34750 39006 34802
rect 39058 34750 39060 34802
rect 38668 34018 38724 34030
rect 38668 33966 38670 34018
rect 38722 33966 38724 34018
rect 38444 31892 38612 31948
rect 38108 30930 38164 30940
rect 37884 30884 37940 30894
rect 37884 30790 37940 30828
rect 38556 30884 38612 31892
rect 38556 30818 38612 30828
rect 38668 30324 38724 33966
rect 39004 33572 39060 34750
rect 39004 33506 39060 33516
rect 39004 33236 39060 33246
rect 39004 33142 39060 33180
rect 39116 33012 39172 35756
rect 39004 32956 39172 33012
rect 38780 32676 38836 32686
rect 38780 32582 38836 32620
rect 38780 31554 38836 31566
rect 38780 31502 38782 31554
rect 38834 31502 38836 31554
rect 38780 31108 38836 31502
rect 38780 31042 38836 31052
rect 38892 31106 38948 31118
rect 38892 31054 38894 31106
rect 38946 31054 38948 31106
rect 38892 30772 38948 31054
rect 38892 30706 38948 30716
rect 39004 30548 39060 32956
rect 39228 32564 39284 37102
rect 39228 32498 39284 32508
rect 39116 31780 39172 31790
rect 39116 31686 39172 31724
rect 39452 31778 39508 38108
rect 39900 35812 39956 35822
rect 39900 35718 39956 35756
rect 40236 33572 40292 38668
rect 41916 38722 41972 38734
rect 41916 38670 41918 38722
rect 41970 38670 41972 38722
rect 41356 38164 41412 38174
rect 41356 38070 41412 38108
rect 41132 37940 41188 37950
rect 40908 36594 40964 36606
rect 40908 36542 40910 36594
rect 40962 36542 40964 36594
rect 40796 35028 40852 35038
rect 40796 34934 40852 34972
rect 40236 33506 40292 33516
rect 40348 34018 40404 34030
rect 40348 33966 40350 34018
rect 40402 33966 40404 34018
rect 40012 33124 40068 33134
rect 40348 33124 40404 33966
rect 40684 33346 40740 33358
rect 40684 33294 40686 33346
rect 40738 33294 40740 33346
rect 40460 33124 40516 33134
rect 40684 33124 40740 33294
rect 39900 33122 40740 33124
rect 39900 33070 40014 33122
rect 40066 33070 40462 33122
rect 40514 33070 40740 33122
rect 39900 33068 40740 33070
rect 39452 31726 39454 31778
rect 39506 31726 39508 31778
rect 39452 31714 39508 31726
rect 39676 32452 39732 32462
rect 39900 32452 39956 33068
rect 40012 33058 40068 33068
rect 40460 33058 40516 33068
rect 40908 33012 40964 36542
rect 40572 32956 40964 33012
rect 39676 32450 39956 32452
rect 39676 32398 39678 32450
rect 39730 32398 39956 32450
rect 39676 32396 39956 32398
rect 40012 32450 40068 32462
rect 40012 32398 40014 32450
rect 40066 32398 40068 32450
rect 39676 31780 39732 32396
rect 39676 31714 39732 31724
rect 40012 31556 40068 32398
rect 38668 30258 38724 30268
rect 38780 30492 39060 30548
rect 39676 31108 39732 31118
rect 37772 30158 37774 30210
rect 37826 30158 37828 30210
rect 37772 30146 37828 30158
rect 38780 29650 38836 30492
rect 39676 30212 39732 31052
rect 39676 30146 39732 30156
rect 39900 30882 39956 30894
rect 39900 30830 39902 30882
rect 39954 30830 39956 30882
rect 38780 29598 38782 29650
rect 38834 29598 38836 29650
rect 38780 29586 38836 29598
rect 37660 28690 37716 28700
rect 37996 29538 38052 29550
rect 37996 29486 37998 29538
rect 38050 29486 38052 29538
rect 37548 28590 37550 28642
rect 37602 28590 37604 28642
rect 37548 28578 37604 28590
rect 37324 28082 37492 28084
rect 37324 28030 37326 28082
rect 37378 28030 37492 28082
rect 37324 28028 37492 28030
rect 37324 28018 37380 28028
rect 37548 27858 37604 27870
rect 37548 27806 37550 27858
rect 37602 27806 37604 27858
rect 37436 27076 37492 27086
rect 37212 27074 37492 27076
rect 37212 27022 37438 27074
rect 37490 27022 37492 27074
rect 37212 27020 37492 27022
rect 37436 27010 37492 27020
rect 36988 24770 37044 24780
rect 37100 26964 37156 26974
rect 37100 24612 37156 26908
rect 37548 26964 37604 27806
rect 37548 26898 37604 26908
rect 37212 26404 37268 26414
rect 37212 25282 37268 26348
rect 37548 26402 37604 26414
rect 37548 26350 37550 26402
rect 37602 26350 37604 26402
rect 37212 25230 37214 25282
rect 37266 25230 37268 25282
rect 37212 25218 37268 25230
rect 37324 25394 37380 25406
rect 37324 25342 37326 25394
rect 37378 25342 37380 25394
rect 37324 25172 37380 25342
rect 37324 25106 37380 25116
rect 37548 24724 37604 26350
rect 37996 25618 38052 29486
rect 39116 29426 39172 29438
rect 39116 29374 39118 29426
rect 39170 29374 39172 29426
rect 37996 25566 37998 25618
rect 38050 25566 38052 25618
rect 37996 25554 38052 25566
rect 38668 27746 38724 27758
rect 38668 27694 38670 27746
rect 38722 27694 38724 27746
rect 38668 26852 38724 27694
rect 37772 25506 37828 25518
rect 37772 25454 37774 25506
rect 37826 25454 37828 25506
rect 37772 25172 37828 25454
rect 38444 25508 38500 25518
rect 38668 25508 38724 26796
rect 38444 25506 38724 25508
rect 38444 25454 38446 25506
rect 38498 25454 38724 25506
rect 38444 25452 38724 25454
rect 39004 25508 39060 25518
rect 37772 25106 37828 25116
rect 37884 25284 37940 25294
rect 37548 24658 37604 24668
rect 36988 24052 37044 24062
rect 36932 24050 37044 24052
rect 36932 23998 36990 24050
rect 37042 23998 37044 24050
rect 36932 23996 37044 23998
rect 36876 23958 36932 23996
rect 36988 23986 37044 23996
rect 37100 24052 37156 24556
rect 37100 23986 37156 23996
rect 37884 23938 37940 25228
rect 38444 25284 38500 25452
rect 39004 25414 39060 25452
rect 38444 25218 38500 25228
rect 38556 24836 38612 24846
rect 38556 24610 38612 24780
rect 38556 24558 38558 24610
rect 38610 24558 38612 24610
rect 38556 24546 38612 24558
rect 37884 23886 37886 23938
rect 37938 23886 37940 23938
rect 37884 23874 37940 23886
rect 38108 24500 38164 24510
rect 37100 23714 37156 23726
rect 37100 23662 37102 23714
rect 37154 23662 37156 23714
rect 37100 23378 37156 23662
rect 37100 23326 37102 23378
rect 37154 23326 37156 23378
rect 37100 23314 37156 23326
rect 38108 23266 38164 24444
rect 39116 24500 39172 29374
rect 39788 28756 39844 28766
rect 39788 26962 39844 28700
rect 39900 28418 39956 30830
rect 40012 29314 40068 31500
rect 40236 32450 40292 32462
rect 40236 32398 40238 32450
rect 40290 32398 40292 32450
rect 40236 29986 40292 32398
rect 40572 31948 40628 32956
rect 40908 32788 40964 32798
rect 40796 32676 40852 32686
rect 40236 29934 40238 29986
rect 40290 29934 40292 29986
rect 40236 29922 40292 29934
rect 40460 31892 40628 31948
rect 40684 32620 40796 32676
rect 40012 29262 40014 29314
rect 40066 29262 40068 29314
rect 40012 29250 40068 29262
rect 39900 28366 39902 28418
rect 39954 28366 39956 28418
rect 39900 28354 39956 28366
rect 39788 26910 39790 26962
rect 39842 26910 39844 26962
rect 39788 26898 39844 26910
rect 40460 26908 40516 31892
rect 40572 30660 40628 30670
rect 40572 28866 40628 30604
rect 40572 28814 40574 28866
rect 40626 28814 40628 28866
rect 40572 28802 40628 28814
rect 40572 27300 40628 27310
rect 40684 27300 40740 32620
rect 40796 32610 40852 32620
rect 40796 31220 40852 31230
rect 40796 29650 40852 31164
rect 40908 30210 40964 32732
rect 41132 32788 41188 37884
rect 41916 36596 41972 38670
rect 41356 36540 41972 36596
rect 42028 37156 42084 37166
rect 41132 32722 41188 32732
rect 41244 34018 41300 34030
rect 41244 33966 41246 34018
rect 41298 33966 41300 34018
rect 41244 33906 41300 33966
rect 41244 33854 41246 33906
rect 41298 33854 41300 33906
rect 41020 32564 41076 32574
rect 41244 32564 41300 33854
rect 41356 33346 41412 36540
rect 41916 36372 41972 36382
rect 41356 33294 41358 33346
rect 41410 33294 41412 33346
rect 41356 33282 41412 33294
rect 41580 36370 41972 36372
rect 41580 36318 41918 36370
rect 41970 36318 41972 36370
rect 41580 36316 41972 36318
rect 41580 32676 41636 36316
rect 41916 36306 41972 36316
rect 42028 36148 42084 37100
rect 41916 36092 42084 36148
rect 42252 36148 42308 39454
rect 43260 38946 43316 38958
rect 43260 38894 43262 38946
rect 43314 38894 43316 38946
rect 42364 37940 42420 37950
rect 42364 37846 42420 37884
rect 42476 37156 42532 37166
rect 42476 37062 42532 37100
rect 42252 36092 42644 36148
rect 41580 32610 41636 32620
rect 41692 35700 41748 35710
rect 41692 34132 41748 35644
rect 41804 35476 41860 35486
rect 41804 35382 41860 35420
rect 41804 34132 41860 34142
rect 41692 34130 41860 34132
rect 41692 34078 41806 34130
rect 41858 34078 41860 34130
rect 41692 34076 41860 34078
rect 41692 33906 41748 34076
rect 41804 34066 41860 34076
rect 41692 33854 41694 33906
rect 41746 33854 41748 33906
rect 41020 32562 41300 32564
rect 41020 32510 41022 32562
rect 41074 32510 41300 32562
rect 41020 32508 41300 32510
rect 41692 32562 41748 33854
rect 41692 32510 41694 32562
rect 41746 32510 41748 32562
rect 41020 32498 41076 32508
rect 40908 30158 40910 30210
rect 40962 30158 40964 30210
rect 40908 30146 40964 30158
rect 41132 31780 41188 32508
rect 41692 32498 41748 32510
rect 41916 31948 41972 36092
rect 42476 35922 42532 35934
rect 42476 35870 42478 35922
rect 42530 35870 42532 35922
rect 42140 34802 42196 34814
rect 42140 34750 42142 34802
rect 42194 34750 42196 34802
rect 42028 32564 42084 32574
rect 42028 32470 42084 32508
rect 41132 30994 41188 31724
rect 41132 30942 41134 30994
rect 41186 30942 41188 30994
rect 41132 30324 41188 30942
rect 40796 29598 40798 29650
rect 40850 29598 40852 29650
rect 40796 29586 40852 29598
rect 41132 29988 41188 30268
rect 41356 31892 41972 31948
rect 41244 29988 41300 29998
rect 41132 29986 41300 29988
rect 41132 29934 41246 29986
rect 41298 29934 41300 29986
rect 41132 29932 41300 29934
rect 40796 28644 40852 28654
rect 41132 28644 41188 29932
rect 41244 29922 41300 29932
rect 40852 28588 41188 28644
rect 41356 28642 41412 31892
rect 42028 31668 42084 31678
rect 42028 31554 42084 31612
rect 42028 31502 42030 31554
rect 42082 31502 42084 31554
rect 42028 31490 42084 31502
rect 41580 30996 41636 31006
rect 41580 30902 41636 30940
rect 42140 30660 42196 34750
rect 42364 34132 42420 34142
rect 42364 34038 42420 34076
rect 42140 30594 42196 30604
rect 42364 33572 42420 33582
rect 42140 30436 42196 30446
rect 42140 30322 42196 30380
rect 42140 30270 42142 30322
rect 42194 30270 42196 30322
rect 42140 30258 42196 30270
rect 41692 30212 41748 30222
rect 41580 30100 41636 30110
rect 41580 29650 41636 30044
rect 41580 29598 41582 29650
rect 41634 29598 41636 29650
rect 41580 29586 41636 29598
rect 41356 28590 41358 28642
rect 41410 28590 41412 28642
rect 40796 28550 40852 28588
rect 41356 28578 41412 28590
rect 40908 28420 40964 28430
rect 40908 27970 40964 28364
rect 41692 28196 41748 30156
rect 40908 27918 40910 27970
rect 40962 27918 40964 27970
rect 40908 27906 40964 27918
rect 41244 28140 41748 28196
rect 41244 27970 41300 28140
rect 41244 27918 41246 27970
rect 41298 27918 41300 27970
rect 41244 27906 41300 27918
rect 41468 27858 41524 27870
rect 41468 27806 41470 27858
rect 41522 27806 41524 27858
rect 41468 27300 41524 27806
rect 40572 27298 40740 27300
rect 40572 27246 40574 27298
rect 40626 27246 40740 27298
rect 40572 27244 40740 27246
rect 41132 27244 41524 27300
rect 42140 27858 42196 27870
rect 42140 27806 42142 27858
rect 42194 27806 42196 27858
rect 40572 27234 40628 27244
rect 40684 27074 40740 27086
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40684 26908 40740 27022
rect 41132 26908 41188 27244
rect 40236 26852 40516 26908
rect 40572 26852 41188 26908
rect 41356 27074 41412 27086
rect 41356 27022 41358 27074
rect 41410 27022 41412 27074
rect 41356 26908 41412 27022
rect 41356 26852 41748 26908
rect 39900 26290 39956 26302
rect 39900 26238 39902 26290
rect 39954 26238 39956 26290
rect 39116 24434 39172 24444
rect 39452 24722 39508 24734
rect 39452 24670 39454 24722
rect 39506 24670 39508 24722
rect 39452 24612 39508 24670
rect 39116 24276 39172 24286
rect 38108 23214 38110 23266
rect 38162 23214 38164 23266
rect 38108 23202 38164 23214
rect 38556 23938 38612 23950
rect 38556 23886 38558 23938
rect 38610 23886 38612 23938
rect 37884 22930 37940 22942
rect 37884 22878 37886 22930
rect 37938 22878 37940 22930
rect 36876 22372 36932 22382
rect 37100 22372 37156 22382
rect 36932 22370 37156 22372
rect 36932 22318 37102 22370
rect 37154 22318 37156 22370
rect 36932 22316 37156 22318
rect 36876 22306 36932 22316
rect 36652 22194 36708 22204
rect 36540 22146 36596 22158
rect 36540 22094 36542 22146
rect 36594 22094 36596 22146
rect 35980 20526 35982 20578
rect 36034 20526 36036 20578
rect 35980 20514 36036 20526
rect 36092 20690 36148 20702
rect 36092 20638 36094 20690
rect 36146 20638 36148 20690
rect 36092 20188 36148 20638
rect 36540 20580 36596 22094
rect 36988 21588 37044 21598
rect 37100 21588 37156 22316
rect 37548 22372 37604 22382
rect 37548 22370 37828 22372
rect 37548 22318 37550 22370
rect 37602 22318 37828 22370
rect 37548 22316 37828 22318
rect 37548 22306 37604 22316
rect 36988 21586 37156 21588
rect 36988 21534 36990 21586
rect 37042 21534 37156 21586
rect 36988 21532 37156 21534
rect 36988 21522 37044 21532
rect 36540 20514 36596 20524
rect 36652 21362 36708 21374
rect 36652 21310 36654 21362
rect 36706 21310 36708 21362
rect 36652 20188 36708 21310
rect 37100 20804 37156 21532
rect 37100 20710 37156 20748
rect 37324 21586 37380 21598
rect 37324 21534 37326 21586
rect 37378 21534 37380 21586
rect 36092 20132 36260 20188
rect 35868 20066 35924 20076
rect 36204 19908 36260 20132
rect 35980 19348 36036 19358
rect 35980 19254 36036 19292
rect 36092 19012 36148 19022
rect 36092 18918 36148 18956
rect 35756 17726 35758 17778
rect 35810 17726 35812 17778
rect 35756 17714 35812 17726
rect 35868 18562 35924 18574
rect 35868 18510 35870 18562
rect 35922 18510 35924 18562
rect 35756 16996 35812 17006
rect 35644 16940 35756 16996
rect 35756 16930 35812 16940
rect 34748 16594 34804 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34860 16100 34916 16110
rect 34748 15204 34804 15214
rect 34076 13766 34132 13804
rect 34300 15092 34356 15102
rect 34300 12850 34356 15036
rect 34636 14868 34692 14878
rect 34636 14642 34692 14812
rect 34636 14590 34638 14642
rect 34690 14590 34692 14642
rect 34636 14578 34692 14590
rect 34524 13860 34580 13870
rect 34524 13766 34580 13804
rect 34300 12798 34302 12850
rect 34354 12798 34356 12850
rect 34300 12786 34356 12798
rect 34412 13412 34468 13422
rect 34412 11282 34468 13356
rect 34412 11230 34414 11282
rect 34466 11230 34468 11282
rect 34412 11218 34468 11230
rect 34412 10500 34468 10510
rect 34412 10406 34468 10444
rect 33964 9662 33966 9714
rect 34018 9662 34020 9714
rect 33964 9650 34020 9662
rect 34748 8930 34804 15148
rect 34860 13858 34916 16044
rect 35868 16100 35924 18510
rect 36092 17780 36148 17790
rect 36204 17780 36260 19852
rect 36092 17778 36260 17780
rect 36092 17726 36094 17778
rect 36146 17726 36260 17778
rect 36092 17724 36260 17726
rect 36428 20132 36708 20188
rect 36092 17714 36148 17724
rect 36428 17556 36484 20132
rect 37324 18676 37380 21534
rect 37436 20972 37716 21028
rect 37436 20802 37492 20972
rect 37436 20750 37438 20802
rect 37490 20750 37492 20802
rect 37436 20738 37492 20750
rect 37548 20804 37604 20814
rect 37324 18610 37380 18620
rect 37436 20580 37492 20590
rect 36988 18452 37044 18462
rect 36988 18358 37044 18396
rect 37324 18340 37380 18350
rect 36652 18228 36708 18238
rect 35868 16034 35924 16044
rect 35980 17500 36484 17556
rect 36540 18226 36708 18228
rect 36540 18174 36654 18226
rect 36706 18174 36708 18226
rect 36540 18172 36708 18174
rect 35756 15874 35812 15886
rect 35980 15876 36036 17500
rect 35756 15822 35758 15874
rect 35810 15822 35812 15874
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35644 14756 35700 14766
rect 35420 14644 35476 14654
rect 35476 14588 35588 14644
rect 35420 14578 35476 14588
rect 35196 14420 35252 14430
rect 34860 13806 34862 13858
rect 34914 13806 34916 13858
rect 34860 13794 34916 13806
rect 35084 14364 35196 14420
rect 34860 13636 34916 13646
rect 34860 13076 34916 13580
rect 34860 12982 34916 13020
rect 35084 13074 35140 14364
rect 35196 14354 35252 14364
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13022 35086 13074
rect 35138 13022 35140 13074
rect 35084 13010 35140 13022
rect 35084 12068 35140 12078
rect 35084 11974 35140 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35532 11506 35588 14588
rect 35644 14418 35700 14700
rect 35644 14366 35646 14418
rect 35698 14366 35700 14418
rect 35644 14354 35700 14366
rect 35756 14420 35812 15822
rect 35756 14354 35812 14364
rect 35868 15820 36036 15876
rect 36092 17106 36148 17118
rect 36092 17054 36094 17106
rect 36146 17054 36148 17106
rect 35868 13300 35924 15820
rect 35980 15314 36036 15326
rect 35980 15262 35982 15314
rect 36034 15262 36036 15314
rect 35980 13524 36036 15262
rect 35980 13458 36036 13468
rect 35868 13244 36036 13300
rect 35868 13076 35924 13086
rect 35868 11508 35924 13020
rect 35980 12852 36036 13244
rect 35980 12786 36036 12796
rect 36092 12628 36148 17054
rect 36204 16996 36260 17006
rect 36204 13634 36260 16940
rect 36316 16772 36372 16782
rect 36372 16716 36484 16772
rect 36316 16706 36372 16716
rect 36204 13582 36206 13634
rect 36258 13582 36260 13634
rect 36204 13570 36260 13582
rect 36316 14308 36372 14318
rect 36204 13076 36260 13086
rect 36316 13076 36372 14252
rect 36204 13074 36372 13076
rect 36204 13022 36206 13074
rect 36258 13022 36372 13074
rect 36204 13020 36372 13022
rect 36204 13010 36260 13020
rect 36092 12572 36260 12628
rect 35532 11454 35534 11506
rect 35586 11454 35588 11506
rect 35532 11442 35588 11454
rect 35644 11506 35924 11508
rect 35644 11454 35870 11506
rect 35922 11454 35924 11506
rect 35644 11452 35924 11454
rect 35308 11394 35364 11406
rect 35308 11342 35310 11394
rect 35362 11342 35364 11394
rect 35308 11284 35364 11342
rect 35644 11284 35700 11452
rect 35868 11442 35924 11452
rect 36204 11506 36260 12572
rect 36428 12290 36484 16716
rect 36540 16100 36596 18172
rect 36652 18162 36708 18172
rect 37324 17668 37380 18284
rect 36988 17666 37380 17668
rect 36988 17614 37326 17666
rect 37378 17614 37380 17666
rect 36988 17612 37380 17614
rect 36652 16996 36708 17006
rect 36652 16902 36708 16940
rect 36540 16034 36596 16044
rect 36764 16884 36820 16894
rect 36988 16884 37044 17612
rect 37324 17602 37380 17612
rect 37324 16884 37380 16894
rect 36820 16882 37044 16884
rect 36820 16830 36990 16882
rect 37042 16830 37044 16882
rect 36820 16828 37044 16830
rect 36428 12238 36430 12290
rect 36482 12238 36484 12290
rect 36428 12226 36484 12238
rect 36540 15874 36596 15886
rect 36540 15822 36542 15874
rect 36594 15822 36596 15874
rect 36204 11454 36206 11506
rect 36258 11454 36260 11506
rect 36204 11442 36260 11454
rect 35308 11228 35700 11284
rect 35420 10724 35476 10734
rect 35420 10630 35476 10668
rect 36540 10724 36596 15822
rect 36652 15316 36708 15326
rect 36764 15316 36820 16828
rect 36988 16818 37044 16828
rect 37212 16882 37380 16884
rect 37212 16830 37326 16882
rect 37378 16830 37380 16882
rect 37212 16828 37380 16830
rect 36652 15314 36820 15316
rect 36652 15262 36654 15314
rect 36706 15262 36820 15314
rect 36652 15260 36820 15262
rect 36876 15874 36932 15886
rect 36876 15822 36878 15874
rect 36930 15822 36932 15874
rect 36652 15250 36708 15260
rect 36876 11732 36932 15822
rect 37100 13860 37156 13870
rect 36876 11666 36932 11676
rect 36988 13804 37100 13860
rect 36540 10658 36596 10668
rect 36988 10388 37044 13804
rect 37100 13794 37156 13804
rect 36428 10332 37044 10388
rect 37100 11172 37156 11182
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35644 9156 35700 9166
rect 35644 9062 35700 9100
rect 34748 8878 34750 8930
rect 34802 8878 34804 8930
rect 34748 8866 34804 8878
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 33852 6038 33908 6076
rect 34188 6804 34244 6814
rect 32844 4958 32846 5010
rect 32898 4958 32900 5010
rect 32844 4946 32900 4958
rect 33068 5906 33124 5918
rect 33068 5854 33070 5906
rect 33122 5854 33124 5906
rect 32172 4900 32228 4910
rect 32172 4898 32452 4900
rect 32172 4846 32174 4898
rect 32226 4846 32452 4898
rect 32172 4844 32452 4846
rect 32172 4834 32228 4844
rect 32172 4564 32228 4574
rect 31948 4562 32228 4564
rect 31948 4510 32174 4562
rect 32226 4510 32228 4562
rect 31948 4508 32228 4510
rect 32172 4498 32228 4508
rect 31164 4452 31220 4462
rect 31164 4358 31220 4396
rect 31388 4338 31444 4350
rect 31388 4286 31390 4338
rect 31442 4286 31444 4338
rect 31388 4004 31444 4286
rect 30940 3948 31444 4004
rect 31836 4338 31892 4350
rect 31836 4286 31838 4338
rect 31890 4286 31892 4338
rect 30492 3668 30548 3678
rect 30492 3574 30548 3612
rect 30940 800 30996 3948
rect 31612 3444 31668 3454
rect 31836 3444 31892 4286
rect 32396 3556 32452 4844
rect 33068 4452 33124 5854
rect 33068 4386 33124 4396
rect 33292 5122 33348 5134
rect 33292 5070 33294 5122
rect 33346 5070 33348 5122
rect 33180 4340 33236 4350
rect 33180 4246 33236 4284
rect 33292 4116 33348 5070
rect 33964 5122 34020 5134
rect 33964 5070 33966 5122
rect 34018 5070 34020 5122
rect 33404 5012 33460 5022
rect 33404 4562 33460 4956
rect 33404 4510 33406 4562
rect 33458 4510 33460 4562
rect 33404 4498 33460 4510
rect 33516 4898 33572 4910
rect 33516 4846 33518 4898
rect 33570 4846 33572 4898
rect 33292 4050 33348 4060
rect 33516 3780 33572 4846
rect 33852 4564 33908 4574
rect 33852 4338 33908 4508
rect 33852 4286 33854 4338
rect 33906 4286 33908 4338
rect 33852 4274 33908 4286
rect 33964 4340 34020 5070
rect 34188 4898 34244 6748
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34188 4846 34190 4898
rect 34242 4846 34244 4898
rect 34188 4834 34244 4846
rect 34748 4900 34804 4910
rect 34748 4898 35028 4900
rect 34748 4846 34750 4898
rect 34802 4846 35028 4898
rect 34748 4844 35028 4846
rect 34748 4834 34804 4844
rect 34076 4788 34132 4798
rect 34076 4562 34132 4732
rect 34076 4510 34078 4562
rect 34130 4510 34132 4562
rect 34076 4498 34132 4510
rect 34524 4450 34580 4462
rect 34524 4398 34526 4450
rect 34578 4398 34580 4450
rect 34524 4340 34580 4398
rect 33964 4284 34580 4340
rect 34748 4340 34804 4350
rect 33516 3714 33572 3724
rect 34076 4116 34132 4126
rect 32956 3668 33012 3678
rect 32620 3666 33012 3668
rect 32620 3614 32958 3666
rect 33010 3614 33012 3666
rect 32620 3612 33012 3614
rect 32508 3556 32564 3566
rect 32396 3554 32564 3556
rect 32396 3502 32510 3554
rect 32562 3502 32564 3554
rect 32396 3500 32564 3502
rect 32508 3490 32564 3500
rect 31612 3442 31892 3444
rect 31612 3390 31614 3442
rect 31666 3390 31892 3442
rect 31612 3388 31892 3390
rect 32620 3388 32676 3612
rect 32956 3602 33012 3612
rect 33628 3556 33684 3566
rect 31612 800 31668 3388
rect 32284 3332 32676 3388
rect 32956 3444 33012 3454
rect 32284 800 32340 3332
rect 32956 800 33012 3388
rect 33628 800 33684 3500
rect 33852 3444 33908 3454
rect 33852 3350 33908 3388
rect 34076 3442 34132 4060
rect 34076 3390 34078 3442
rect 34130 3390 34132 3442
rect 34076 3378 34132 3390
rect 34300 3554 34356 3566
rect 34300 3502 34302 3554
rect 34354 3502 34356 3554
rect 34300 3444 34356 3502
rect 34300 3378 34356 3388
rect 34748 3442 34804 4284
rect 34748 3390 34750 3442
rect 34802 3390 34804 3442
rect 34748 3378 34804 3390
rect 34860 4338 34916 4350
rect 34860 4286 34862 4338
rect 34914 4286 34916 4338
rect 34860 4228 34916 4286
rect 34860 1764 34916 4172
rect 34972 3556 35028 4844
rect 35644 4898 35700 4910
rect 35644 4846 35646 4898
rect 35698 4846 35700 4898
rect 35420 4564 35476 4574
rect 35420 4470 35476 4508
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34972 3490 35028 3500
rect 34300 1708 34916 1764
rect 34972 3332 35028 3342
rect 34300 800 34356 1708
rect 34972 800 35028 3276
rect 35644 3108 35700 4846
rect 36428 4564 36484 10332
rect 37100 9828 37156 11116
rect 37212 9940 37268 16828
rect 37324 16818 37380 16828
rect 37324 16100 37380 16110
rect 37324 12290 37380 16044
rect 37436 13858 37492 20524
rect 37548 18338 37604 20748
rect 37660 18564 37716 20972
rect 37660 18498 37716 18508
rect 37548 18286 37550 18338
rect 37602 18286 37604 18338
rect 37548 18274 37604 18286
rect 37660 17666 37716 17678
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 37548 15874 37604 15886
rect 37548 15822 37550 15874
rect 37602 15822 37604 15874
rect 37548 14308 37604 15822
rect 37660 15204 37716 17614
rect 37660 15138 37716 15148
rect 37772 14644 37828 22316
rect 37884 21588 37940 22878
rect 37884 21522 37940 21532
rect 37996 22260 38052 22270
rect 37996 20020 38052 22204
rect 38556 22036 38612 23886
rect 39116 23042 39172 24220
rect 39116 22990 39118 23042
rect 39170 22990 39172 23042
rect 39116 22978 39172 22990
rect 39228 23156 39284 23166
rect 38556 21970 38612 21980
rect 37996 19954 38052 19964
rect 38108 21924 38164 21934
rect 37996 14644 38052 14654
rect 37772 14642 38052 14644
rect 37772 14590 37998 14642
rect 38050 14590 38052 14642
rect 37772 14588 38052 14590
rect 37996 14578 38052 14588
rect 37548 14242 37604 14252
rect 37436 13806 37438 13858
rect 37490 13806 37492 13858
rect 37436 13794 37492 13806
rect 37324 12238 37326 12290
rect 37378 12238 37380 12290
rect 37324 12226 37380 12238
rect 37436 13524 37492 13534
rect 37436 10498 37492 13468
rect 38108 13074 38164 21868
rect 39004 21588 39060 21598
rect 38892 20132 38948 20142
rect 38892 20038 38948 20076
rect 38332 19794 38388 19806
rect 38332 19742 38334 19794
rect 38386 19742 38388 19794
rect 38332 19684 38388 19742
rect 38388 19628 38500 19684
rect 38332 19618 38388 19628
rect 38332 16660 38388 16670
rect 38332 15202 38388 16604
rect 38332 15150 38334 15202
rect 38386 15150 38388 15202
rect 38332 15138 38388 15150
rect 38444 15092 38500 19628
rect 38556 19346 38612 19358
rect 38556 19294 38558 19346
rect 38610 19294 38612 19346
rect 38556 18340 38612 19294
rect 38556 18274 38612 18284
rect 38892 18564 38948 18574
rect 38780 15540 38836 15550
rect 38444 13746 38500 15036
rect 38444 13694 38446 13746
rect 38498 13694 38500 13746
rect 38444 13682 38500 13694
rect 38556 15484 38780 15540
rect 38556 13634 38612 15484
rect 38780 15474 38836 15484
rect 38892 15148 38948 18508
rect 38556 13582 38558 13634
rect 38610 13582 38612 13634
rect 38556 13570 38612 13582
rect 38780 15092 38948 15148
rect 38108 13022 38110 13074
rect 38162 13022 38164 13074
rect 38108 13010 38164 13022
rect 38668 12068 38724 12078
rect 38780 12068 38836 15092
rect 39004 14418 39060 21532
rect 39228 20130 39284 23100
rect 39228 20078 39230 20130
rect 39282 20078 39284 20130
rect 39228 19908 39284 20078
rect 39228 19842 39284 19852
rect 39452 19234 39508 24556
rect 39676 24724 39732 24734
rect 39452 19182 39454 19234
rect 39506 19182 39508 19234
rect 39452 18452 39508 19182
rect 39452 18358 39508 18396
rect 39564 23940 39620 23950
rect 39452 16772 39508 16782
rect 39004 14366 39006 14418
rect 39058 14366 39060 14418
rect 39004 14354 39060 14366
rect 39228 15428 39284 15438
rect 39116 12852 39172 12862
rect 39116 12758 39172 12796
rect 38668 12066 38836 12068
rect 38668 12014 38670 12066
rect 38722 12014 38836 12066
rect 38668 12012 38836 12014
rect 38668 12002 38724 12012
rect 37996 11508 38052 11518
rect 37996 11414 38052 11452
rect 39228 11282 39284 15372
rect 39452 15426 39508 16716
rect 39452 15374 39454 15426
rect 39506 15374 39508 15426
rect 39452 15362 39508 15374
rect 39564 15148 39620 23884
rect 39676 23266 39732 24668
rect 39900 24164 39956 26238
rect 40236 25508 40292 26852
rect 40460 26292 40516 26302
rect 40572 26292 40628 26796
rect 40460 26290 40628 26292
rect 40460 26238 40462 26290
rect 40514 26238 40628 26290
rect 40460 26236 40628 26238
rect 41020 26292 41076 26302
rect 41132 26292 41188 26852
rect 41020 26290 41188 26292
rect 41020 26238 41022 26290
rect 41074 26238 41188 26290
rect 41020 26236 41188 26238
rect 40460 26226 40516 26236
rect 41020 26226 41076 26236
rect 40236 25442 40292 25452
rect 41020 24836 41076 24846
rect 41020 24742 41076 24780
rect 41132 24724 41188 26236
rect 41468 26292 41524 26302
rect 41468 26290 41636 26292
rect 41468 26238 41470 26290
rect 41522 26238 41636 26290
rect 41468 26236 41636 26238
rect 41468 26226 41524 26236
rect 41468 25396 41524 25406
rect 41468 25282 41524 25340
rect 41468 25230 41470 25282
rect 41522 25230 41524 25282
rect 41468 25218 41524 25230
rect 41356 24724 41412 24734
rect 41132 24722 41412 24724
rect 41132 24670 41358 24722
rect 41410 24670 41412 24722
rect 41132 24668 41412 24670
rect 41356 24658 41412 24668
rect 41580 24164 41636 26236
rect 39900 24098 39956 24108
rect 41468 24108 41636 24164
rect 40012 23716 40068 23726
rect 40796 23716 40852 23726
rect 39676 23214 39678 23266
rect 39730 23214 39732 23266
rect 39676 23202 39732 23214
rect 39900 23660 40012 23716
rect 39900 22146 39956 23660
rect 40012 23650 40068 23660
rect 40348 23714 40852 23716
rect 40348 23662 40798 23714
rect 40850 23662 40852 23714
rect 40348 23660 40852 23662
rect 40012 23156 40068 23166
rect 40012 23062 40068 23100
rect 39900 22094 39902 22146
rect 39954 22094 39956 22146
rect 39900 22082 39956 22094
rect 40012 22484 40068 22494
rect 39900 21810 39956 21822
rect 39900 21758 39902 21810
rect 39954 21758 39956 21810
rect 39788 20018 39844 20030
rect 39788 19966 39790 20018
rect 39842 19966 39844 20018
rect 39788 19684 39844 19966
rect 39788 19618 39844 19628
rect 39900 19348 39956 21758
rect 40012 20578 40068 22428
rect 40012 20526 40014 20578
rect 40066 20526 40068 20578
rect 40012 20514 40068 20526
rect 40348 20242 40404 23660
rect 40796 23650 40852 23660
rect 40908 23268 40964 23278
rect 40908 23174 40964 23212
rect 41132 23268 41188 23278
rect 41132 23154 41188 23212
rect 41132 23102 41134 23154
rect 41186 23102 41188 23154
rect 41132 23090 41188 23102
rect 40684 22540 40964 22596
rect 40572 22484 40628 22494
rect 40684 22484 40740 22540
rect 40572 22482 40740 22484
rect 40572 22430 40574 22482
rect 40626 22430 40740 22482
rect 40572 22428 40740 22430
rect 40572 22418 40628 22428
rect 40796 22372 40852 22382
rect 40796 21586 40852 22316
rect 40796 21534 40798 21586
rect 40850 21534 40852 21586
rect 40348 20190 40350 20242
rect 40402 20190 40404 20242
rect 40348 20178 40404 20190
rect 40460 21362 40516 21374
rect 40460 21310 40462 21362
rect 40514 21310 40516 21362
rect 40460 20132 40516 21310
rect 40684 20804 40740 20814
rect 40796 20804 40852 21534
rect 40740 20748 40852 20804
rect 40684 20710 40740 20748
rect 40460 20066 40516 20076
rect 40572 20578 40628 20590
rect 40572 20526 40574 20578
rect 40626 20526 40628 20578
rect 39900 19282 39956 19292
rect 40124 18676 40180 18686
rect 40012 17442 40068 17454
rect 40012 17390 40014 17442
rect 40066 17390 40068 17442
rect 39676 16994 39732 17006
rect 39676 16942 39678 16994
rect 39730 16942 39732 16994
rect 39676 15540 39732 16942
rect 39676 15474 39732 15484
rect 39900 16098 39956 16110
rect 39900 16046 39902 16098
rect 39954 16046 39956 16098
rect 39564 15092 39732 15148
rect 39228 11230 39230 11282
rect 39282 11230 39284 11282
rect 39228 11218 39284 11230
rect 39340 11732 39396 11742
rect 38668 10724 38724 10734
rect 38668 10630 38724 10668
rect 37436 10446 37438 10498
rect 37490 10446 37492 10498
rect 37436 10434 37492 10446
rect 38332 9940 38388 9950
rect 37212 9938 38388 9940
rect 37212 9886 38334 9938
rect 38386 9886 38388 9938
rect 37212 9884 38388 9886
rect 38332 9874 38388 9884
rect 37100 9762 37156 9772
rect 39340 9714 39396 11676
rect 39676 11284 39732 15092
rect 39788 15092 39844 15102
rect 39788 14530 39844 15036
rect 39788 14478 39790 14530
rect 39842 14478 39844 14530
rect 39788 14466 39844 14478
rect 39900 13524 39956 16046
rect 40012 14642 40068 17390
rect 40012 14590 40014 14642
rect 40066 14590 40068 14642
rect 40012 14578 40068 14590
rect 40012 13524 40068 13534
rect 39900 13468 40012 13524
rect 40012 13458 40068 13468
rect 40124 12068 40180 18620
rect 40348 18452 40404 18462
rect 40348 18358 40404 18396
rect 40572 17892 40628 20526
rect 40796 18228 40852 18238
rect 40348 17836 40628 17892
rect 40684 18226 40852 18228
rect 40684 18174 40798 18226
rect 40850 18174 40852 18226
rect 40684 18172 40852 18174
rect 40124 12002 40180 12012
rect 40236 15204 40292 15214
rect 39676 11218 39732 11228
rect 39340 9662 39342 9714
rect 39394 9662 39396 9714
rect 39340 9650 39396 9662
rect 38556 9604 38612 9614
rect 37100 7476 37156 7486
rect 37100 5012 37156 7420
rect 38556 6804 38612 9548
rect 40236 8370 40292 15148
rect 40348 12292 40404 17836
rect 40572 16884 40628 16894
rect 40348 12226 40404 12236
rect 40460 16658 40516 16670
rect 40460 16606 40462 16658
rect 40514 16606 40516 16658
rect 40460 8428 40516 16606
rect 40572 16098 40628 16828
rect 40572 16046 40574 16098
rect 40626 16046 40628 16098
rect 40572 16034 40628 16046
rect 40684 12852 40740 18172
rect 40796 18162 40852 18172
rect 40908 18228 40964 22540
rect 41356 22370 41412 22382
rect 41356 22318 41358 22370
rect 41410 22318 41412 22370
rect 41020 22036 41076 22046
rect 41020 18676 41076 21980
rect 41356 21924 41412 22318
rect 41356 21858 41412 21868
rect 41468 21812 41524 24108
rect 41580 23940 41636 23950
rect 41580 23846 41636 23884
rect 41692 23604 41748 26852
rect 42028 26852 42084 26862
rect 42028 25844 42084 26796
rect 42140 26068 42196 27806
rect 42364 26852 42420 33516
rect 42476 31892 42532 35870
rect 42476 31826 42532 31836
rect 42588 31890 42644 36092
rect 43260 33796 43316 38894
rect 43260 33730 43316 33740
rect 43820 37378 43876 37390
rect 43820 37326 43822 37378
rect 43874 37326 43876 37378
rect 42588 31838 42590 31890
rect 42642 31838 42644 31890
rect 42588 31826 42644 31838
rect 43596 33122 43652 33134
rect 43596 33070 43598 33122
rect 43650 33070 43652 33122
rect 43036 31778 43092 31790
rect 43036 31726 43038 31778
rect 43090 31726 43092 31778
rect 42812 31668 42868 31678
rect 42812 31574 42868 31612
rect 43036 31556 43092 31726
rect 43036 31490 43092 31500
rect 43596 30660 43652 33070
rect 43820 32564 43876 37326
rect 44044 32564 44100 32574
rect 43820 32508 44044 32564
rect 44044 32498 44100 32508
rect 44156 31948 44212 40238
rect 44380 37044 44436 37054
rect 44380 33570 44436 36988
rect 44380 33518 44382 33570
rect 44434 33518 44436 33570
rect 44380 33506 44436 33518
rect 44044 31892 44212 31948
rect 44492 32786 44548 32798
rect 44492 32734 44494 32786
rect 44546 32734 44548 32786
rect 43708 31666 43764 31678
rect 43708 31614 43710 31666
rect 43762 31614 43764 31666
rect 43708 31444 43764 31614
rect 43708 31378 43764 31388
rect 43820 31554 43876 31566
rect 43820 31502 43822 31554
rect 43874 31502 43876 31554
rect 43820 31218 43876 31502
rect 43820 31166 43822 31218
rect 43874 31166 43876 31218
rect 43820 31154 43876 31166
rect 44044 30996 44100 31892
rect 44044 30930 44100 30940
rect 44380 31556 44436 31566
rect 43596 30594 43652 30604
rect 43820 30884 43876 30894
rect 43148 30098 43204 30110
rect 43148 30046 43150 30098
rect 43202 30046 43204 30098
rect 43148 28868 43204 30046
rect 43820 29426 43876 30828
rect 44268 30884 44324 30894
rect 44044 30212 44100 30222
rect 44268 30212 44324 30828
rect 44100 30210 44324 30212
rect 44100 30158 44270 30210
rect 44322 30158 44324 30210
rect 44100 30156 44324 30158
rect 44044 30146 44100 30156
rect 44268 30146 44324 30156
rect 44380 30324 44436 31500
rect 44492 30772 44548 32734
rect 44604 31218 44660 42028
rect 44828 41074 44884 42140
rect 44828 41022 44830 41074
rect 44882 41022 44884 41074
rect 44828 41010 44884 41022
rect 44940 41858 44996 41870
rect 44940 41806 44942 41858
rect 44994 41806 44996 41858
rect 44716 38724 44772 38734
rect 44716 38630 44772 38668
rect 44940 35698 44996 41806
rect 45164 41076 45220 41086
rect 45164 40982 45220 41020
rect 45836 41076 45892 41086
rect 45836 40982 45892 41020
rect 46060 40626 46116 42364
rect 46284 41858 46340 41870
rect 46284 41806 46286 41858
rect 46338 41806 46340 41858
rect 46172 41076 46228 41086
rect 46284 41076 46340 41806
rect 46228 41020 46340 41076
rect 46508 41748 46564 41758
rect 46172 40982 46228 41020
rect 46060 40574 46062 40626
rect 46114 40574 46116 40626
rect 46060 40562 46116 40574
rect 45388 40514 45444 40526
rect 45388 40462 45390 40514
rect 45442 40462 45444 40514
rect 45388 37044 45444 40462
rect 46508 40292 46564 41692
rect 46172 40236 46564 40292
rect 46172 39506 46228 40236
rect 46172 39454 46174 39506
rect 46226 39454 46228 39506
rect 46172 39442 46228 39454
rect 45724 38948 45780 38958
rect 45724 38854 45780 38892
rect 45388 36978 45444 36988
rect 45500 36260 45556 36270
rect 44940 35646 44942 35698
rect 44994 35646 44996 35698
rect 44940 35634 44996 35646
rect 45388 35700 45444 35710
rect 45388 35606 45444 35644
rect 44940 34354 44996 34366
rect 44940 34302 44942 34354
rect 44994 34302 44996 34354
rect 44940 31948 44996 34302
rect 45500 34354 45556 36204
rect 45500 34302 45502 34354
rect 45554 34302 45556 34354
rect 45500 34290 45556 34302
rect 45164 33796 45220 33806
rect 45164 32786 45220 33740
rect 45164 32734 45166 32786
rect 45218 32734 45220 32786
rect 45164 32722 45220 32734
rect 45164 32564 45220 32574
rect 44940 31892 45108 31948
rect 44940 31556 44996 31566
rect 44940 31462 44996 31500
rect 45052 31332 45108 31892
rect 44604 31166 44606 31218
rect 44658 31166 44660 31218
rect 44604 31154 44660 31166
rect 44940 31276 45108 31332
rect 44828 30882 44884 30894
rect 44828 30830 44830 30882
rect 44882 30830 44884 30882
rect 44828 30772 44884 30830
rect 44492 30716 44884 30772
rect 43820 29374 43822 29426
rect 43874 29374 43876 29426
rect 43820 29362 43876 29374
rect 43932 30098 43988 30110
rect 43932 30046 43934 30098
rect 43986 30046 43988 30098
rect 43148 28802 43204 28812
rect 43932 28756 43988 30046
rect 44380 29428 44436 30268
rect 44828 30100 44884 30110
rect 44828 30006 44884 30044
rect 44940 29650 44996 31276
rect 44940 29598 44942 29650
rect 44994 29598 44996 29650
rect 44940 29586 44996 29598
rect 45052 30996 45108 31006
rect 45052 30210 45108 30940
rect 45052 30158 45054 30210
rect 45106 30158 45108 30210
rect 44380 29426 44996 29428
rect 44380 29374 44382 29426
rect 44434 29374 44996 29426
rect 44380 29372 44996 29374
rect 44380 29362 44436 29372
rect 43932 28690 43988 28700
rect 44940 28866 44996 29372
rect 45052 29316 45108 30158
rect 45052 29222 45108 29260
rect 44940 28814 44942 28866
rect 44994 28814 44996 28866
rect 44940 28754 44996 28814
rect 44940 28702 44942 28754
rect 44994 28702 44996 28754
rect 44940 28690 44996 28702
rect 43596 28418 43652 28430
rect 43596 28366 43598 28418
rect 43650 28366 43652 28418
rect 43596 26908 43652 28366
rect 44380 28420 44436 28430
rect 44380 28418 44996 28420
rect 44380 28366 44382 28418
rect 44434 28366 44996 28418
rect 44380 28364 44996 28366
rect 44380 28354 44436 28364
rect 44268 28196 44324 28206
rect 44268 27300 44324 28140
rect 44604 28082 44660 28094
rect 44604 28030 44606 28082
rect 44658 28030 44660 28082
rect 44380 27300 44436 27310
rect 44268 27298 44436 27300
rect 44268 27246 44382 27298
rect 44434 27246 44436 27298
rect 44268 27244 44436 27246
rect 44380 27234 44436 27244
rect 42364 26786 42420 26796
rect 43484 26852 43652 26908
rect 43820 26852 43876 26862
rect 43484 26404 43540 26852
rect 43820 26758 43876 26796
rect 43820 26514 43876 26526
rect 43820 26462 43822 26514
rect 43874 26462 43876 26514
rect 43596 26404 43652 26414
rect 43484 26348 43596 26404
rect 43596 26338 43652 26348
rect 43372 26068 43428 26078
rect 42140 26012 42756 26068
rect 42028 25788 42196 25844
rect 42028 25284 42084 25294
rect 41692 23538 41748 23548
rect 41804 25282 42084 25284
rect 41804 25230 42030 25282
rect 42082 25230 42084 25282
rect 41804 25228 42084 25230
rect 41468 21746 41524 21756
rect 41468 21588 41524 21598
rect 41468 21494 41524 21532
rect 41244 20804 41300 20814
rect 41244 20710 41300 20748
rect 41804 19684 41860 25228
rect 42028 25218 42084 25228
rect 42028 24724 42084 24734
rect 42140 24724 42196 25788
rect 42028 24722 42196 24724
rect 42028 24670 42030 24722
rect 42082 24670 42196 24722
rect 42028 24668 42196 24670
rect 42252 25394 42308 25406
rect 42252 25342 42254 25394
rect 42306 25342 42308 25394
rect 42252 25284 42308 25342
rect 42028 24658 42084 24668
rect 42252 24052 42308 25228
rect 41916 23996 42308 24052
rect 42364 25282 42420 25294
rect 42364 25230 42366 25282
rect 42418 25230 42420 25282
rect 41916 23268 41972 23996
rect 42364 23716 42420 25230
rect 42476 24276 42532 24286
rect 42476 24050 42532 24220
rect 42476 23998 42478 24050
rect 42530 23998 42532 24050
rect 42476 23986 42532 23998
rect 42364 23650 42420 23660
rect 41916 23202 41972 23212
rect 42252 23604 42308 23614
rect 42028 23154 42084 23166
rect 42028 23102 42030 23154
rect 42082 23102 42084 23154
rect 42028 22372 42084 23102
rect 42028 22306 42084 22316
rect 41916 19908 41972 19918
rect 41916 19814 41972 19852
rect 41804 19628 41972 19684
rect 41132 19346 41188 19358
rect 41132 19294 41134 19346
rect 41186 19294 41188 19346
rect 41132 19012 41188 19294
rect 41132 18946 41188 18956
rect 41020 18620 41188 18676
rect 40908 18162 40964 18172
rect 40796 17444 40852 17454
rect 40796 17350 40852 17388
rect 41132 17220 41188 18620
rect 41580 18564 41636 18574
rect 41580 18470 41636 18508
rect 40796 17164 41188 17220
rect 41356 18340 41412 18350
rect 40796 13076 40852 17164
rect 41132 16996 41188 17006
rect 41020 16884 41076 16894
rect 40908 16828 41020 16884
rect 40908 16098 40964 16828
rect 41020 16790 41076 16828
rect 40908 16046 40910 16098
rect 40962 16046 40964 16098
rect 40908 16034 40964 16046
rect 41132 15988 41188 16940
rect 41356 16884 41412 18284
rect 41356 16660 41412 16828
rect 41468 16884 41524 16894
rect 41468 16882 41860 16884
rect 41468 16830 41470 16882
rect 41522 16830 41860 16882
rect 41468 16828 41860 16830
rect 41468 16818 41524 16828
rect 41356 16604 41748 16660
rect 41356 16100 41412 16110
rect 41356 16098 41524 16100
rect 41356 16046 41358 16098
rect 41410 16046 41524 16098
rect 41356 16044 41524 16046
rect 41356 16034 41412 16044
rect 41020 15932 41188 15988
rect 41020 15538 41076 15932
rect 41020 15486 41022 15538
rect 41074 15486 41076 15538
rect 41020 15474 41076 15486
rect 41132 15316 41188 15326
rect 41468 15316 41524 16044
rect 40908 15260 41132 15316
rect 40908 15092 40964 15260
rect 41132 15222 41188 15260
rect 41356 15260 41524 15316
rect 41692 15314 41748 16604
rect 41692 15262 41694 15314
rect 41746 15262 41748 15314
rect 40908 15026 40964 15036
rect 41244 15204 41300 15214
rect 41132 13524 41188 13534
rect 41020 13076 41076 13086
rect 40796 13074 41076 13076
rect 40796 13022 41022 13074
rect 41074 13022 41076 13074
rect 40796 13020 41076 13022
rect 41020 13010 41076 13020
rect 40684 12796 41076 12852
rect 41020 9154 41076 12796
rect 41132 9938 41188 13468
rect 41244 11508 41300 15148
rect 41356 11732 41412 15260
rect 41692 15250 41748 15262
rect 41804 15148 41860 16828
rect 41356 11666 41412 11676
rect 41468 15092 41860 15148
rect 41356 11508 41412 11518
rect 41244 11452 41356 11508
rect 41356 11442 41412 11452
rect 41132 9886 41134 9938
rect 41186 9886 41188 9938
rect 41132 9874 41188 9886
rect 41020 9102 41022 9154
rect 41074 9102 41076 9154
rect 41020 9090 41076 9102
rect 40460 8372 41300 8428
rect 40236 8318 40238 8370
rect 40290 8318 40292 8370
rect 40236 8306 40292 8318
rect 41244 8146 41300 8372
rect 41244 8094 41246 8146
rect 41298 8094 41300 8146
rect 41244 8082 41300 8094
rect 41468 7362 41524 15092
rect 41916 14980 41972 19628
rect 42140 19124 42196 19134
rect 42140 19030 42196 19068
rect 41916 14914 41972 14924
rect 42028 18228 42084 18238
rect 42028 12850 42084 18172
rect 42252 17778 42308 23548
rect 42588 23156 42644 23166
rect 42476 23154 42644 23156
rect 42476 23102 42590 23154
rect 42642 23102 42644 23154
rect 42476 23100 42644 23102
rect 42476 18340 42532 23100
rect 42588 23090 42644 23100
rect 42476 18274 42532 18284
rect 42588 21588 42644 21598
rect 42252 17726 42254 17778
rect 42306 17726 42308 17778
rect 42252 17714 42308 17726
rect 42028 12798 42030 12850
rect 42082 12798 42084 12850
rect 42028 12786 42084 12798
rect 42140 17444 42196 17454
rect 41916 12068 41972 12078
rect 41916 11974 41972 12012
rect 42028 11732 42084 11742
rect 42028 8932 42084 11676
rect 42140 10388 42196 17388
rect 42364 15314 42420 15326
rect 42364 15262 42366 15314
rect 42418 15262 42420 15314
rect 42252 11508 42308 11518
rect 42252 11414 42308 11452
rect 42364 10612 42420 15262
rect 42476 13860 42532 13870
rect 42476 13766 42532 13804
rect 42588 12068 42644 21532
rect 42700 15148 42756 26012
rect 43148 25506 43204 25518
rect 43148 25454 43150 25506
rect 43202 25454 43204 25506
rect 42924 25396 42980 25406
rect 42924 25302 42980 25340
rect 43148 25396 43204 25454
rect 43148 24276 43204 25340
rect 43148 24210 43204 24220
rect 42812 24052 42868 24062
rect 42812 23958 42868 23996
rect 43372 21812 43428 26012
rect 43820 25618 43876 26462
rect 44604 26516 44660 28030
rect 44940 27074 44996 28364
rect 45164 28196 45220 32508
rect 45836 31892 45892 31902
rect 45612 30884 45668 30894
rect 45612 30790 45668 30828
rect 45724 30660 45780 30670
rect 45724 30322 45780 30604
rect 45724 30270 45726 30322
rect 45778 30270 45780 30322
rect 45724 30258 45780 30270
rect 45500 30098 45556 30110
rect 45500 30046 45502 30098
rect 45554 30046 45556 30098
rect 45500 29316 45556 30046
rect 45836 29538 45892 31836
rect 45836 29486 45838 29538
rect 45890 29486 45892 29538
rect 45836 29474 45892 29486
rect 46172 30884 46228 30894
rect 45388 28866 45444 28878
rect 45388 28814 45390 28866
rect 45442 28814 45444 28866
rect 45388 28754 45444 28814
rect 45388 28702 45390 28754
rect 45442 28702 45444 28754
rect 45388 28690 45444 28702
rect 44940 27022 44942 27074
rect 44994 27022 44996 27074
rect 44940 27010 44996 27022
rect 45052 28140 45220 28196
rect 45052 26908 45108 28140
rect 45164 27634 45220 27646
rect 45164 27582 45166 27634
rect 45218 27582 45220 27634
rect 45164 27076 45220 27582
rect 45164 27010 45220 27020
rect 44604 26450 44660 26460
rect 44828 26852 44884 26862
rect 44716 26180 44772 26190
rect 44604 26178 44772 26180
rect 44604 26126 44718 26178
rect 44770 26126 44772 26178
rect 44604 26124 44772 26126
rect 44492 26068 44548 26078
rect 44492 25974 44548 26012
rect 43820 25566 43822 25618
rect 43874 25566 43876 25618
rect 43820 25554 43876 25566
rect 43596 25396 43652 25406
rect 43596 25302 43652 25340
rect 44492 24948 44548 24958
rect 44604 24948 44660 26124
rect 44716 26114 44772 26124
rect 44828 25618 44884 26796
rect 44828 25566 44830 25618
rect 44882 25566 44884 25618
rect 44828 25554 44884 25566
rect 44940 26852 45108 26908
rect 44492 24946 44660 24948
rect 44492 24894 44494 24946
rect 44546 24894 44660 24946
rect 44492 24892 44660 24894
rect 44940 24948 44996 26852
rect 45388 26404 45444 26414
rect 45388 26310 45444 26348
rect 45052 26180 45108 26190
rect 45164 26180 45220 26190
rect 45052 26178 45164 26180
rect 45052 26126 45054 26178
rect 45106 26126 45164 26178
rect 45052 26124 45164 26126
rect 45052 26114 45108 26124
rect 45164 25394 45220 26124
rect 45164 25342 45166 25394
rect 45218 25342 45220 25394
rect 45052 24948 45108 24958
rect 44940 24946 45108 24948
rect 44940 24894 45054 24946
rect 45106 24894 45108 24946
rect 44940 24892 45108 24894
rect 44492 24882 44548 24892
rect 45052 24882 45108 24892
rect 44492 24276 44548 24286
rect 43820 23828 43876 23838
rect 43820 23734 43876 23772
rect 43820 22148 43876 22158
rect 44380 22148 44436 22158
rect 43820 22054 43876 22092
rect 43932 22146 44436 22148
rect 43932 22094 44382 22146
rect 44434 22094 44436 22146
rect 43932 22092 44436 22094
rect 43260 21756 43428 21812
rect 42924 20132 42980 20142
rect 42924 20038 42980 20076
rect 42924 19684 42980 19694
rect 42924 19234 42980 19628
rect 42924 19182 42926 19234
rect 42978 19182 42980 19234
rect 42924 19170 42980 19182
rect 43260 17554 43316 21756
rect 43708 21700 43764 21710
rect 43484 21698 43764 21700
rect 43484 21646 43710 21698
rect 43762 21646 43764 21698
rect 43484 21644 43764 21646
rect 43260 17502 43262 17554
rect 43314 17502 43316 17554
rect 43260 17490 43316 17502
rect 43372 20244 43428 20254
rect 42700 15092 42868 15148
rect 42812 14642 42868 15092
rect 42812 14590 42814 14642
rect 42866 14590 42868 14642
rect 42812 14578 42868 14590
rect 42812 13746 42868 13758
rect 42812 13694 42814 13746
rect 42866 13694 42868 13746
rect 42812 13636 42868 13694
rect 43260 13636 43316 13646
rect 42812 13634 43316 13636
rect 42812 13582 43262 13634
rect 43314 13582 43316 13634
rect 42812 13580 43316 13582
rect 43260 12852 43316 13580
rect 43260 12786 43316 12796
rect 43036 12738 43092 12750
rect 43036 12686 43038 12738
rect 43090 12686 43092 12738
rect 43036 12628 43092 12686
rect 43036 12562 43092 12572
rect 42924 12292 42980 12302
rect 42924 12198 42980 12236
rect 42588 12012 42980 12068
rect 42140 10322 42196 10332
rect 42252 10556 42420 10612
rect 42140 10052 42196 10062
rect 42140 9714 42196 9996
rect 42140 9662 42142 9714
rect 42194 9662 42196 9714
rect 42140 9650 42196 9662
rect 42140 8932 42196 8942
rect 42028 8930 42196 8932
rect 42028 8878 42142 8930
rect 42194 8878 42196 8930
rect 42028 8876 42196 8878
rect 42140 8866 42196 8876
rect 42252 8708 42308 10556
rect 42924 10498 42980 12012
rect 43260 11284 43316 11294
rect 43372 11284 43428 20188
rect 43484 19458 43540 21644
rect 43708 21634 43764 21644
rect 43820 21364 43876 21374
rect 43708 20580 43764 20590
rect 43484 19406 43486 19458
rect 43538 19406 43540 19458
rect 43484 19394 43540 19406
rect 43596 20524 43708 20580
rect 43596 15986 43652 20524
rect 43708 20514 43764 20524
rect 43820 20578 43876 21308
rect 43820 20526 43822 20578
rect 43874 20526 43876 20578
rect 43820 20514 43876 20526
rect 43820 19906 43876 19918
rect 43820 19854 43822 19906
rect 43874 19854 43876 19906
rect 43820 19794 43876 19854
rect 43820 19742 43822 19794
rect 43874 19742 43876 19794
rect 43820 19730 43876 19742
rect 43820 19348 43876 19358
rect 43820 19254 43876 19292
rect 43820 18450 43876 18462
rect 43820 18398 43822 18450
rect 43874 18398 43876 18450
rect 43820 17108 43876 18398
rect 43820 17042 43876 17052
rect 43708 16996 43764 17006
rect 43708 16902 43764 16940
rect 43596 15934 43598 15986
rect 43650 15934 43652 15986
rect 43596 15922 43652 15934
rect 43932 14418 43988 22092
rect 44380 22082 44436 22092
rect 44044 21700 44100 21710
rect 44044 18900 44100 21644
rect 44492 21588 44548 24220
rect 45052 24276 45108 24286
rect 45164 24276 45220 25342
rect 45500 25618 45556 29260
rect 45836 27972 45892 27982
rect 45836 27878 45892 27916
rect 46060 27858 46116 27870
rect 46060 27806 46062 27858
rect 46114 27806 46116 27858
rect 45612 27748 45668 27758
rect 46060 27748 46116 27806
rect 45612 27746 46116 27748
rect 45612 27694 45614 27746
rect 45666 27694 46116 27746
rect 45612 27692 46116 27694
rect 45612 27682 45668 27692
rect 45948 27076 46004 27086
rect 45724 26962 45780 26974
rect 45724 26910 45726 26962
rect 45778 26910 45780 26962
rect 45724 26908 45780 26910
rect 45724 26852 45892 26908
rect 45612 26516 45668 26526
rect 45612 25732 45668 26460
rect 45836 26292 45892 26852
rect 45836 26226 45892 26236
rect 45724 26180 45780 26190
rect 45724 26086 45780 26124
rect 45612 25676 45780 25732
rect 45500 25566 45502 25618
rect 45554 25566 45556 25618
rect 45500 24834 45556 25566
rect 45500 24782 45502 24834
rect 45554 24782 45556 24834
rect 45500 24770 45556 24782
rect 45612 25282 45668 25294
rect 45612 25230 45614 25282
rect 45666 25230 45668 25282
rect 45108 24220 45220 24276
rect 44940 24164 44996 24174
rect 44828 23826 44884 23838
rect 44828 23774 44830 23826
rect 44882 23774 44884 23826
rect 44828 22484 44884 23774
rect 44828 22418 44884 22428
rect 44828 22148 44884 22158
rect 44828 22054 44884 22092
rect 44156 21532 44548 21588
rect 44156 19906 44212 21532
rect 44492 21362 44548 21374
rect 44492 21310 44494 21362
rect 44546 21310 44548 21362
rect 44380 20578 44436 20590
rect 44380 20526 44382 20578
rect 44434 20526 44436 20578
rect 44380 20468 44436 20526
rect 44380 20402 44436 20412
rect 44492 20244 44548 21310
rect 44716 21364 44772 21374
rect 44716 21270 44772 21308
rect 44828 20580 44884 20618
rect 44828 20514 44884 20524
rect 44492 20178 44548 20188
rect 44828 20356 44884 20366
rect 44156 19854 44158 19906
rect 44210 19854 44212 19906
rect 44156 19346 44212 19854
rect 44156 19294 44158 19346
rect 44210 19294 44212 19346
rect 44156 19282 44212 19294
rect 44492 19906 44548 19918
rect 44492 19854 44494 19906
rect 44546 19854 44548 19906
rect 44044 18844 44212 18900
rect 43932 14366 43934 14418
rect 43986 14366 43988 14418
rect 43932 14354 43988 14366
rect 44044 18676 44100 18686
rect 44044 14196 44100 18620
rect 44156 15148 44212 18844
rect 44492 18676 44548 19854
rect 44492 18610 44548 18620
rect 44380 18450 44436 18462
rect 44380 18398 44382 18450
rect 44434 18398 44436 18450
rect 44268 17556 44324 17566
rect 44268 17462 44324 17500
rect 44380 16884 44436 18398
rect 44716 18340 44772 18350
rect 44380 16818 44436 16828
rect 44492 16996 44548 17006
rect 44492 16882 44548 16940
rect 44492 16830 44494 16882
rect 44546 16830 44548 16882
rect 44492 16818 44548 16830
rect 44380 15874 44436 15886
rect 44380 15822 44382 15874
rect 44434 15822 44436 15874
rect 44156 15092 44324 15148
rect 43708 14140 44100 14196
rect 43260 11282 43428 11284
rect 43260 11230 43262 11282
rect 43314 11230 43428 11282
rect 43260 11228 43428 11230
rect 43484 13860 43540 13870
rect 43260 11218 43316 11228
rect 42924 10446 42926 10498
rect 42978 10446 42980 10498
rect 42924 10434 42980 10446
rect 42476 10388 42532 10398
rect 42532 10332 42644 10388
rect 42476 10322 42532 10332
rect 41468 7310 41470 7362
rect 41522 7310 41524 7362
rect 41468 7298 41524 7310
rect 41916 8652 42308 8708
rect 42476 10164 42532 10174
rect 38556 6738 38612 6748
rect 41916 6802 41972 8652
rect 42476 8596 42532 10108
rect 41916 6750 41918 6802
rect 41970 6750 41972 6802
rect 41916 6738 41972 6750
rect 42252 8540 42532 8596
rect 38556 6468 38612 6478
rect 37660 5124 37716 5134
rect 38332 5124 38388 5134
rect 37660 5122 38164 5124
rect 37660 5070 37662 5122
rect 37714 5070 38164 5122
rect 37660 5068 38164 5070
rect 37660 5058 37716 5068
rect 37100 4946 37156 4956
rect 36428 4498 36484 4508
rect 37212 4900 37268 4910
rect 37212 4562 37268 4844
rect 37212 4510 37214 4562
rect 37266 4510 37268 4562
rect 37212 4498 37268 4510
rect 37884 4898 37940 4910
rect 37884 4846 37886 4898
rect 37938 4846 37940 4898
rect 35868 4452 35924 4462
rect 35868 4358 35924 4396
rect 36092 4338 36148 4350
rect 36092 4286 36094 4338
rect 36146 4286 36148 4338
rect 35980 3332 36036 3342
rect 35980 3238 36036 3276
rect 36092 3108 36148 4286
rect 36652 4228 36708 4238
rect 37660 4228 37716 4238
rect 36652 4134 36708 4172
rect 37436 4226 37716 4228
rect 37436 4174 37662 4226
rect 37714 4174 37716 4226
rect 37436 4172 37716 4174
rect 36540 3780 36596 3790
rect 35644 3052 36148 3108
rect 36316 3668 36372 3678
rect 35644 800 35700 3052
rect 36316 800 36372 3612
rect 36540 3554 36596 3724
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 36540 3502 36542 3554
rect 36594 3502 36596 3554
rect 36540 3490 36596 3502
rect 37436 3388 37492 4172
rect 37660 4162 37716 4172
rect 37884 4004 37940 4846
rect 37884 3938 37940 3948
rect 37884 3444 37940 3454
rect 37212 3332 37492 3388
rect 37660 3442 38052 3444
rect 37660 3390 37886 3442
rect 37938 3390 38052 3442
rect 37660 3388 38052 3390
rect 37212 980 37268 3332
rect 36988 924 37268 980
rect 36988 800 37044 924
rect 37660 800 37716 3388
rect 37884 3378 37940 3388
rect 37996 3220 38052 3388
rect 38108 3442 38164 5068
rect 38332 5122 38500 5124
rect 38332 5070 38334 5122
rect 38386 5070 38500 5122
rect 38332 5068 38500 5070
rect 38332 5058 38388 5068
rect 38444 4452 38500 5068
rect 38556 5010 38612 6412
rect 39116 5124 39172 5134
rect 39116 5122 39956 5124
rect 39116 5070 39118 5122
rect 39170 5070 39956 5122
rect 39116 5068 39956 5070
rect 39116 5058 39172 5068
rect 38556 4958 38558 5010
rect 38610 4958 38612 5010
rect 38556 4946 38612 4958
rect 39340 4900 39396 4910
rect 39340 4806 39396 4844
rect 39900 4562 39956 5068
rect 39900 4510 39902 4562
rect 39954 4510 39956 4562
rect 39900 4498 39956 4510
rect 40124 5122 40180 5134
rect 40124 5070 40126 5122
rect 40178 5070 40180 5122
rect 40124 4564 40180 5070
rect 40348 5124 40404 5134
rect 40348 5010 40404 5068
rect 40348 4958 40350 5010
rect 40402 4958 40404 5010
rect 40348 4946 40404 4958
rect 41692 5122 41748 5134
rect 41692 5070 41694 5122
rect 41746 5070 41748 5122
rect 41692 5012 41748 5070
rect 41692 4956 42196 5012
rect 40908 4900 40964 4910
rect 41356 4900 41412 4910
rect 40908 4898 41076 4900
rect 40908 4846 40910 4898
rect 40962 4846 41076 4898
rect 40908 4844 41076 4846
rect 40908 4834 40964 4844
rect 40124 4498 40180 4508
rect 40908 4564 40964 4574
rect 40908 4470 40964 4508
rect 38444 4396 38836 4452
rect 38556 4226 38612 4238
rect 38556 4174 38558 4226
rect 38610 4174 38612 4226
rect 38108 3390 38110 3442
rect 38162 3390 38164 3442
rect 38108 3378 38164 3390
rect 38444 3442 38500 3454
rect 38444 3390 38446 3442
rect 38498 3390 38500 3442
rect 38444 3388 38500 3390
rect 38220 3332 38500 3388
rect 38556 3444 38612 4174
rect 38220 3220 38276 3332
rect 37996 3164 38276 3220
rect 38556 1764 38612 3388
rect 38780 3442 38836 4396
rect 40124 4338 40180 4350
rect 40124 4286 40126 4338
rect 40178 4286 40180 4338
rect 39676 4228 39732 4238
rect 40124 4228 40180 4286
rect 41020 4340 41076 4844
rect 41132 4340 41188 4350
rect 41020 4338 41188 4340
rect 41020 4286 41134 4338
rect 41186 4286 41188 4338
rect 41020 4284 41188 4286
rect 39676 4226 40180 4228
rect 39676 4174 39678 4226
rect 39730 4174 40180 4226
rect 39676 4172 40180 4174
rect 38780 3390 38782 3442
rect 38834 3390 38836 3442
rect 38780 3378 38836 3390
rect 39004 3668 39060 3678
rect 38332 1708 38612 1764
rect 38332 800 38388 1708
rect 39004 800 39060 3612
rect 39116 3444 39172 3454
rect 39116 3350 39172 3388
rect 39676 800 39732 4172
rect 39788 4004 39844 4014
rect 39788 3554 39844 3948
rect 40236 3668 40292 3678
rect 40236 3574 40292 3612
rect 39788 3502 39790 3554
rect 39842 3502 39844 3554
rect 39788 3490 39844 3502
rect 41132 3108 41188 4284
rect 41356 3554 41412 4844
rect 41916 4450 41972 4462
rect 41916 4398 41918 4450
rect 41970 4398 41972 4450
rect 41916 4116 41972 4398
rect 41916 4050 41972 4060
rect 42140 4338 42196 4956
rect 42252 4788 42308 8540
rect 42588 8428 42644 10332
rect 43260 9602 43316 9614
rect 43260 9550 43262 9602
rect 43314 9550 43316 9602
rect 43260 9044 43316 9550
rect 43260 8978 43316 8988
rect 43484 8428 43540 13804
rect 43596 13524 43652 13534
rect 43596 13074 43652 13468
rect 43596 13022 43598 13074
rect 43650 13022 43652 13074
rect 43596 13010 43652 13022
rect 43596 12180 43652 12190
rect 43596 10052 43652 12124
rect 43596 9986 43652 9996
rect 43596 9714 43652 9726
rect 43596 9662 43598 9714
rect 43650 9662 43652 9714
rect 43596 9492 43652 9662
rect 43596 9426 43652 9436
rect 42364 8372 42644 8428
rect 42812 8372 43540 8428
rect 43708 8428 43764 14140
rect 43820 13636 43876 13646
rect 43820 10164 43876 13580
rect 44268 13634 44324 15092
rect 44380 13860 44436 15822
rect 44380 13794 44436 13804
rect 44268 13582 44270 13634
rect 44322 13582 44324 13634
rect 44268 13570 44324 13582
rect 44268 12740 44324 12750
rect 44268 12646 44324 12684
rect 44716 12066 44772 18284
rect 44828 15538 44884 20300
rect 44940 19906 44996 24108
rect 45052 23938 45108 24220
rect 45612 23940 45668 25230
rect 45724 24610 45780 25676
rect 45724 24558 45726 24610
rect 45778 24558 45780 24610
rect 45724 24546 45780 24558
rect 45052 23886 45054 23938
rect 45106 23886 45108 23938
rect 45052 23874 45108 23886
rect 45276 23884 45668 23940
rect 45724 24276 45780 24286
rect 45164 23380 45220 23390
rect 45276 23380 45332 23884
rect 45612 23716 45668 23726
rect 45724 23716 45780 24220
rect 45612 23714 45724 23716
rect 45612 23662 45614 23714
rect 45666 23662 45724 23714
rect 45612 23660 45724 23662
rect 45612 23650 45668 23660
rect 45724 23622 45780 23660
rect 45164 23378 45332 23380
rect 45164 23326 45166 23378
rect 45218 23326 45332 23378
rect 45164 23324 45332 23326
rect 45164 23314 45220 23324
rect 45724 22932 45780 22942
rect 45500 22930 45780 22932
rect 45500 22878 45726 22930
rect 45778 22878 45780 22930
rect 45500 22876 45780 22878
rect 44940 19854 44942 19906
rect 44994 19854 44996 19906
rect 44940 19842 44996 19854
rect 45052 22370 45108 22382
rect 45052 22318 45054 22370
rect 45106 22318 45108 22370
rect 45052 21588 45108 22318
rect 45052 20802 45108 21532
rect 45052 20750 45054 20802
rect 45106 20750 45108 20802
rect 45052 19684 45108 20750
rect 45052 19618 45108 19628
rect 44940 19234 44996 19246
rect 44940 19182 44942 19234
rect 44994 19182 44996 19234
rect 44940 18676 44996 19182
rect 44940 18610 44996 18620
rect 44940 18450 44996 18462
rect 44940 18398 44942 18450
rect 44994 18398 44996 18450
rect 44940 17556 44996 18398
rect 45164 17668 45220 17678
rect 45164 17666 45332 17668
rect 45164 17614 45166 17666
rect 45218 17614 45332 17666
rect 45164 17612 45332 17614
rect 45164 17602 45220 17612
rect 44940 17490 44996 17500
rect 44940 17108 44996 17118
rect 44996 17052 45220 17108
rect 44940 17042 44996 17052
rect 44828 15486 44830 15538
rect 44882 15486 44884 15538
rect 44828 15474 44884 15486
rect 44940 16882 44996 16894
rect 44940 16830 44942 16882
rect 44994 16830 44996 16882
rect 44828 14530 44884 14542
rect 44828 14478 44830 14530
rect 44882 14478 44884 14530
rect 44828 13636 44884 14478
rect 44828 13570 44884 13580
rect 44716 12014 44718 12066
rect 44770 12014 44772 12066
rect 44716 12002 44772 12014
rect 44940 11844 44996 16830
rect 45052 12964 45108 12974
rect 45052 12870 45108 12908
rect 44604 11788 44996 11844
rect 43932 11284 43988 11294
rect 43932 10722 43988 11228
rect 43932 10670 43934 10722
rect 43986 10670 43988 10722
rect 43932 10658 43988 10670
rect 44044 10836 44100 10846
rect 43820 10098 43876 10108
rect 44044 9826 44100 10780
rect 44044 9774 44046 9826
rect 44098 9774 44100 9826
rect 44044 9762 44100 9774
rect 44268 9604 44324 9614
rect 44156 9602 44324 9604
rect 44156 9550 44270 9602
rect 44322 9550 44324 9602
rect 44156 9548 44324 9550
rect 43932 9492 43988 9502
rect 43932 9266 43988 9436
rect 43932 9214 43934 9266
rect 43986 9214 43988 9266
rect 43932 9202 43988 9214
rect 43708 8372 43876 8428
rect 42364 7586 42420 8372
rect 42364 7534 42366 7586
rect 42418 7534 42420 7586
rect 42364 7522 42420 7534
rect 42812 6578 42868 8372
rect 42812 6526 42814 6578
rect 42866 6526 42868 6578
rect 42812 6514 42868 6526
rect 42252 4722 42308 4732
rect 42364 5796 42420 5806
rect 42140 4286 42142 4338
rect 42194 4286 42196 4338
rect 41804 3668 41860 3678
rect 41356 3502 41358 3554
rect 41410 3502 41412 3554
rect 41356 3490 41412 3502
rect 41468 3666 41860 3668
rect 41468 3614 41806 3666
rect 41858 3614 41860 3666
rect 41468 3612 41860 3614
rect 40348 3052 41188 3108
rect 40348 800 40404 3052
rect 41468 1764 41524 3612
rect 41804 3602 41860 3612
rect 42140 3444 42196 4286
rect 42364 4228 42420 5740
rect 43820 5684 43876 8372
rect 43932 8036 43988 8046
rect 43932 7942 43988 7980
rect 43820 5618 43876 5628
rect 44044 6580 44100 6590
rect 44044 5122 44100 6524
rect 44044 5070 44046 5122
rect 44098 5070 44100 5122
rect 44044 5058 44100 5070
rect 43596 4900 43652 4910
rect 43596 4806 43652 4844
rect 42364 4162 42420 4172
rect 43596 4450 43652 4462
rect 44044 4452 44100 4462
rect 43596 4398 43598 4450
rect 43650 4398 43652 4450
rect 43596 4116 43652 4398
rect 43596 4050 43652 4060
rect 43820 4450 44100 4452
rect 43820 4398 44046 4450
rect 44098 4398 44100 4450
rect 43820 4396 44100 4398
rect 42700 3668 42756 3678
rect 42700 3574 42756 3612
rect 43820 3556 43876 4396
rect 44044 4386 44100 4396
rect 44156 4452 44212 9548
rect 44268 9538 44324 9548
rect 44268 8820 44324 8830
rect 44268 8146 44324 8764
rect 44604 8428 44660 11788
rect 44940 11172 44996 11182
rect 44940 11078 44996 11116
rect 44828 10836 44884 10846
rect 44828 10742 44884 10780
rect 44940 9604 44996 9614
rect 44940 9510 44996 9548
rect 44716 8932 44772 8942
rect 44716 8838 44772 8876
rect 44604 8372 44772 8428
rect 44268 8094 44270 8146
rect 44322 8094 44324 8146
rect 44268 7700 44324 8094
rect 44604 7700 44660 7710
rect 44268 7698 44660 7700
rect 44268 7646 44606 7698
rect 44658 7646 44660 7698
rect 44268 7644 44660 7646
rect 44604 7634 44660 7644
rect 44380 6804 44436 6814
rect 44268 6748 44380 6804
rect 44268 5010 44324 6748
rect 44380 6738 44436 6748
rect 44268 4958 44270 5010
rect 44322 4958 44324 5010
rect 44268 4946 44324 4958
rect 44716 4562 44772 8372
rect 44940 8036 44996 8046
rect 44940 7942 44996 7980
rect 44940 7476 44996 7486
rect 44940 7382 44996 7420
rect 44940 6468 44996 6478
rect 44940 6374 44996 6412
rect 45164 5908 45220 17052
rect 45276 6804 45332 17612
rect 45500 16772 45556 22876
rect 45724 22866 45780 22876
rect 45612 21588 45668 21598
rect 45612 21494 45668 21532
rect 45724 21474 45780 21486
rect 45724 21422 45726 21474
rect 45778 21422 45780 21474
rect 45724 20356 45780 21422
rect 45724 20290 45780 20300
rect 45836 20578 45892 20590
rect 45836 20526 45838 20578
rect 45890 20526 45892 20578
rect 45724 20132 45780 20142
rect 45724 20038 45780 20076
rect 45500 16706 45556 16716
rect 45724 18564 45780 18574
rect 45500 16212 45556 16222
rect 45500 16118 45556 16156
rect 45500 15540 45556 15550
rect 45388 15428 45444 15438
rect 45388 15334 45444 15372
rect 45388 14980 45444 14990
rect 45388 13858 45444 14924
rect 45388 13806 45390 13858
rect 45442 13806 45444 13858
rect 45388 13794 45444 13806
rect 45500 13074 45556 15484
rect 45724 15538 45780 18508
rect 45724 15486 45726 15538
rect 45778 15486 45780 15538
rect 45724 15474 45780 15486
rect 45612 15316 45668 15326
rect 45612 15222 45668 15260
rect 45500 13022 45502 13074
rect 45554 13022 45556 13074
rect 45500 13010 45556 13022
rect 45724 14868 45780 14878
rect 45724 11618 45780 14812
rect 45724 11566 45726 11618
rect 45778 11566 45780 11618
rect 45724 11554 45780 11566
rect 45612 11508 45668 11518
rect 45500 10498 45556 10510
rect 45500 10446 45502 10498
rect 45554 10446 45556 10498
rect 45500 10164 45556 10446
rect 45500 10098 45556 10108
rect 45388 10052 45444 10062
rect 45388 9938 45444 9996
rect 45388 9886 45390 9938
rect 45442 9886 45444 9938
rect 45388 9874 45444 9886
rect 45612 8370 45668 11452
rect 45724 10724 45780 10734
rect 45724 10630 45780 10668
rect 45612 8318 45614 8370
rect 45666 8318 45668 8370
rect 45612 8306 45668 8318
rect 45276 6738 45332 6748
rect 45724 7476 45780 7486
rect 44940 5852 45220 5908
rect 45612 6692 45668 6702
rect 44940 5794 44996 5852
rect 44940 5742 44942 5794
rect 44994 5742 44996 5794
rect 44940 5730 44996 5742
rect 45500 5460 45556 5470
rect 44940 5124 44996 5134
rect 44940 5030 44996 5068
rect 44716 4510 44718 4562
rect 44770 4510 44772 4562
rect 44716 4498 44772 4510
rect 44156 4386 44212 4396
rect 45164 4450 45220 4462
rect 45164 4398 45166 4450
rect 45218 4398 45220 4450
rect 44492 4338 44548 4350
rect 44492 4286 44494 4338
rect 44546 4286 44548 4338
rect 44492 4228 44548 4286
rect 45164 4228 45220 4398
rect 45500 4450 45556 5404
rect 45612 5234 45668 6636
rect 45724 6690 45780 7420
rect 45724 6638 45726 6690
rect 45778 6638 45780 6690
rect 45724 6626 45780 6638
rect 45836 6580 45892 20526
rect 45948 16660 46004 27020
rect 46060 26964 46116 27692
rect 46060 26898 46116 26908
rect 46172 27186 46228 30828
rect 46172 27134 46174 27186
rect 46226 27134 46228 27186
rect 46172 26290 46228 27134
rect 46172 26238 46174 26290
rect 46226 26238 46228 26290
rect 46060 26180 46116 26190
rect 46172 26180 46228 26238
rect 46116 26124 46228 26180
rect 46060 26114 46116 26124
rect 46060 23716 46116 23726
rect 46060 23378 46116 23660
rect 46060 23326 46062 23378
rect 46114 23326 46116 23378
rect 46060 23314 46116 23326
rect 46284 22148 46340 22158
rect 46172 22146 46340 22148
rect 46172 22094 46286 22146
rect 46338 22094 46340 22146
rect 46172 22092 46340 22094
rect 46172 20690 46228 22092
rect 46284 22082 46340 22092
rect 46172 20638 46174 20690
rect 46226 20638 46228 20690
rect 46172 19572 46228 20638
rect 46172 19506 46228 19516
rect 46284 20468 46340 20478
rect 46060 19124 46116 19134
rect 46060 19030 46116 19068
rect 46060 18338 46116 18350
rect 46060 18286 46062 18338
rect 46114 18286 46116 18338
rect 46060 18228 46116 18286
rect 46060 18162 46116 18172
rect 46060 17556 46116 17566
rect 46060 17462 46116 17500
rect 46060 16884 46116 16894
rect 46060 16790 46116 16828
rect 45948 16604 46116 16660
rect 45948 16098 46004 16110
rect 45948 16046 45950 16098
rect 46002 16046 46004 16098
rect 45948 14644 46004 16046
rect 45948 14578 46004 14588
rect 45948 14420 46004 14430
rect 45948 14326 46004 14364
rect 45948 12292 46004 12302
rect 46060 12292 46116 16604
rect 46172 12964 46228 12974
rect 46172 12870 46228 12908
rect 45948 12290 46116 12292
rect 45948 12238 45950 12290
rect 46002 12238 46116 12290
rect 45948 12236 46116 12238
rect 45948 12226 46004 12236
rect 46060 10610 46116 10622
rect 46060 10558 46062 10610
rect 46114 10558 46116 10610
rect 46060 10164 46116 10558
rect 46060 10098 46116 10108
rect 46284 9940 46340 20412
rect 46060 9884 46340 9940
rect 46508 16996 46564 17006
rect 46060 9154 46116 9884
rect 46060 9102 46062 9154
rect 46114 9102 46116 9154
rect 46060 9090 46116 9102
rect 46508 9044 46564 16940
rect 46172 8988 46564 9044
rect 46620 14644 46676 14654
rect 46172 8932 46228 8988
rect 45836 6514 45892 6524
rect 45948 8876 46228 8932
rect 45948 6018 46004 8876
rect 46620 8820 46676 14588
rect 46284 8764 46676 8820
rect 46060 8148 46116 8158
rect 46060 7586 46116 8092
rect 46060 7534 46062 7586
rect 46114 7534 46116 7586
rect 46060 7522 46116 7534
rect 46172 6132 46228 6142
rect 45948 5966 45950 6018
rect 46002 5966 46004 6018
rect 45948 5954 46004 5966
rect 46060 6076 46172 6132
rect 45612 5182 45614 5234
rect 45666 5182 45668 5234
rect 45612 5170 45668 5182
rect 45500 4398 45502 4450
rect 45554 4398 45556 4450
rect 45500 4386 45556 4398
rect 45836 4452 45892 4462
rect 45836 4358 45892 4396
rect 44492 4172 45220 4228
rect 45612 4228 45668 4238
rect 45668 4172 45780 4228
rect 45612 4162 45668 4172
rect 43596 3500 43876 3556
rect 41916 3388 42196 3444
rect 43036 3444 43092 3454
rect 41916 3108 41972 3388
rect 43036 3330 43092 3388
rect 43036 3278 43038 3330
rect 43090 3278 43092 3330
rect 43036 3266 43092 3278
rect 41020 1708 41524 1764
rect 41692 3052 41972 3108
rect 41020 800 41076 1708
rect 41692 800 41748 3052
rect 43596 1428 43652 3500
rect 45724 3444 45780 4172
rect 46060 3668 46116 6076
rect 46172 6066 46228 6076
rect 46172 5460 46228 5470
rect 46172 5234 46228 5404
rect 46172 5182 46174 5234
rect 46226 5182 46228 5234
rect 46172 5170 46228 5182
rect 46172 4564 46228 4574
rect 46284 4564 46340 8764
rect 46172 4562 46340 4564
rect 46172 4510 46174 4562
rect 46226 4510 46340 4562
rect 46172 4508 46340 4510
rect 46172 4498 46228 4508
rect 46060 3554 46116 3612
rect 46060 3502 46062 3554
rect 46114 3502 46116 3554
rect 46060 3490 46116 3502
rect 45836 3444 45892 3454
rect 45724 3442 45892 3444
rect 45724 3390 45838 3442
rect 45890 3390 45892 3442
rect 45724 3388 45892 3390
rect 45836 3378 45892 3388
rect 43932 3330 43988 3342
rect 43932 3278 43934 3330
rect 43986 3278 43988 3330
rect 43932 2434 43988 3278
rect 43932 2382 43934 2434
rect 43986 2382 43988 2434
rect 43932 2370 43988 2382
rect 44380 3330 44436 3342
rect 44380 3278 44382 3330
rect 44434 3278 44436 3330
rect 44380 2100 44436 3278
rect 44380 2034 44436 2044
rect 44828 3330 44884 3342
rect 44828 3278 44830 3330
rect 44882 3278 44884 3330
rect 43596 1362 43652 1372
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
rect 40320 0 40432 800
rect 40992 0 41104 800
rect 41664 0 41776 800
rect 42336 0 42448 800
rect 43008 0 43120 800
rect 43680 0 43792 800
rect 44352 0 44464 800
rect 44828 756 44884 3278
rect 45276 3330 45332 3342
rect 45276 3278 45278 3330
rect 45330 3278 45332 3330
rect 45276 2772 45332 3278
rect 45276 2706 45332 2716
rect 45276 2434 45332 2446
rect 45276 2382 45278 2434
rect 45330 2382 45332 2434
rect 44828 690 44884 700
rect 45024 0 45136 800
rect 45276 84 45332 2382
rect 45276 18 45332 28
rect 45696 0 45808 800
rect 46368 0 46480 800
rect 47040 0 47152 800
rect 47712 0 47824 800
<< via2 >>
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 8092 44492 8148 44548
rect 9772 44492 9828 44548
rect 14812 44156 14868 44212
rect 15932 44210 15988 44212
rect 15932 44158 15934 44210
rect 15934 44158 15986 44210
rect 15986 44158 15988 44210
rect 15932 44156 15988 44158
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 7756 44044 7812 44100
rect 9324 44098 9380 44100
rect 9324 44046 9326 44098
rect 9326 44046 9378 44098
rect 9378 44046 9380 44098
rect 9324 44044 9380 44046
rect 18732 42700 18788 42756
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20860 43538 20916 43540
rect 20860 43486 20862 43538
rect 20862 43486 20914 43538
rect 20914 43486 20916 43538
rect 20860 43484 20916 43486
rect 20636 42754 20692 42756
rect 20636 42702 20638 42754
rect 20638 42702 20690 42754
rect 20690 42702 20692 42754
rect 20636 42700 20692 42702
rect 21532 43484 21588 43540
rect 21420 42700 21476 42756
rect 22092 43538 22148 43540
rect 22092 43486 22094 43538
rect 22094 43486 22146 43538
rect 22146 43486 22148 43538
rect 22092 43484 22148 43486
rect 1708 42530 1764 42532
rect 1708 42478 1710 42530
rect 1710 42478 1762 42530
rect 1762 42478 1764 42530
rect 1708 42476 1764 42478
rect 22988 43484 23044 43540
rect 23324 43596 23380 43652
rect 22428 42754 22484 42756
rect 22428 42702 22430 42754
rect 22430 42702 22482 42754
rect 22482 42702 22484 42754
rect 22428 42700 22484 42702
rect 23996 43650 24052 43652
rect 23996 43598 23998 43650
rect 23998 43598 24050 43650
rect 24050 43598 24052 43650
rect 23996 43596 24052 43598
rect 24892 44492 24948 44548
rect 25564 44546 25620 44548
rect 25564 44494 25566 44546
rect 25566 44494 25618 44546
rect 25618 44494 25620 44546
rect 25564 44492 25620 44494
rect 25340 44434 25396 44436
rect 25340 44382 25342 44434
rect 25342 44382 25394 44434
rect 25394 44382 25396 44434
rect 25340 44380 25396 44382
rect 24220 43596 24276 43652
rect 25228 43650 25284 43652
rect 25228 43598 25230 43650
rect 25230 43598 25282 43650
rect 25282 43598 25284 43650
rect 25228 43596 25284 43598
rect 23772 43538 23828 43540
rect 23772 43486 23774 43538
rect 23774 43486 23826 43538
rect 23826 43486 23828 43538
rect 23772 43484 23828 43486
rect 24332 43538 24388 43540
rect 24332 43486 24334 43538
rect 24334 43486 24386 43538
rect 24386 43486 24388 43538
rect 24332 43484 24388 43486
rect 27580 45276 27636 45332
rect 26908 44380 26964 44436
rect 28812 45276 28868 45332
rect 29596 44492 29652 44548
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 27804 43484 27860 43540
rect 27132 42194 27188 42196
rect 27132 42142 27134 42194
rect 27134 42142 27186 42194
rect 27186 42142 27188 42194
rect 27132 42140 27188 42142
rect 28476 43538 28532 43540
rect 28476 43486 28478 43538
rect 28478 43486 28530 43538
rect 28530 43486 28532 43538
rect 28476 43484 28532 43486
rect 29820 43538 29876 43540
rect 29820 43486 29822 43538
rect 29822 43486 29874 43538
rect 29874 43486 29876 43538
rect 29820 43484 29876 43486
rect 28476 42924 28532 42980
rect 27580 42028 27636 42084
rect 30380 44492 30436 44548
rect 30940 44492 30996 44548
rect 30156 43484 30212 43540
rect 29932 42140 29988 42196
rect 32620 44492 32676 44548
rect 31612 43650 31668 43652
rect 31612 43598 31614 43650
rect 31614 43598 31666 43650
rect 31666 43598 31668 43650
rect 31612 43596 31668 43598
rect 30716 43538 30772 43540
rect 30716 43486 30718 43538
rect 30718 43486 30770 43538
rect 30770 43486 30772 43538
rect 30716 43484 30772 43486
rect 30492 42194 30548 42196
rect 30492 42142 30494 42194
rect 30494 42142 30546 42194
rect 30546 42142 30548 42194
rect 30492 42140 30548 42142
rect 32060 43596 32116 43652
rect 33740 42924 33796 42980
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 36316 44492 36372 44548
rect 37100 44492 37156 44548
rect 36764 44434 36820 44436
rect 36764 44382 36766 44434
rect 36766 44382 36818 44434
rect 36818 44382 36820 44434
rect 36764 44380 36820 44382
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34860 42700 34916 42756
rect 32172 42140 32228 42196
rect 31836 42028 31892 42084
rect 39004 44492 39060 44548
rect 38780 44380 38836 44436
rect 38892 44268 38948 44324
rect 38220 42754 38276 42756
rect 38220 42702 38222 42754
rect 38222 42702 38274 42754
rect 38274 42702 38276 42754
rect 38220 42700 38276 42702
rect 38556 43484 38612 43540
rect 39004 43538 39060 43540
rect 39004 43486 39006 43538
rect 39006 43486 39058 43538
rect 39058 43486 39060 43538
rect 39004 43484 39060 43486
rect 40236 44492 40292 44548
rect 39676 42754 39732 42756
rect 39676 42702 39678 42754
rect 39678 42702 39730 42754
rect 39730 42702 39732 42754
rect 39676 42700 39732 42702
rect 39900 42642 39956 42644
rect 39900 42590 39902 42642
rect 39902 42590 39954 42642
rect 39954 42590 39956 42642
rect 39900 42588 39956 42590
rect 42364 44492 42420 44548
rect 44044 44492 44100 44548
rect 45724 44380 45780 44436
rect 43708 44322 43764 44324
rect 43708 44270 43710 44322
rect 43710 44270 43762 44322
rect 43762 44270 43764 44322
rect 43708 44268 43764 44270
rect 44044 44044 44100 44100
rect 41804 43596 41860 43652
rect 42588 43650 42644 43652
rect 42588 43598 42590 43650
rect 42590 43598 42642 43650
rect 42642 43598 42644 43650
rect 42588 43596 42644 43598
rect 43036 43596 43092 43652
rect 42812 42700 42868 42756
rect 45612 43708 45668 43764
rect 41244 42588 41300 42644
rect 45836 44098 45892 44100
rect 45836 44046 45838 44098
rect 45838 44046 45890 44098
rect 45890 44046 45892 44098
rect 45836 44044 45892 44046
rect 46172 43708 46228 43764
rect 46060 43036 46116 43092
rect 46060 42364 46116 42420
rect 35532 41916 35588 41972
rect 37100 41970 37156 41972
rect 37100 41918 37102 41970
rect 37102 41918 37154 41970
rect 37154 41918 37156 41970
rect 37100 41916 37156 41918
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 38556 39676 38612 39732
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 36316 38892 36372 38948
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 17052 37884 17108 37940
rect 12796 37324 12852 37380
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1708 34748 1764 34804
rect 2044 31500 2100 31556
rect 1596 30380 1652 30436
rect 5852 34018 5908 34020
rect 5852 33966 5854 34018
rect 5854 33966 5906 34018
rect 5906 33966 5908 34018
rect 5852 33964 5908 33966
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2940 32562 2996 32564
rect 2940 32510 2942 32562
rect 2942 32510 2994 32562
rect 2994 32510 2996 32562
rect 2940 32508 2996 32510
rect 3612 32508 3668 32564
rect 7308 34802 7364 34804
rect 7308 34750 7310 34802
rect 7310 34750 7362 34802
rect 7362 34750 7364 34802
rect 7308 34748 7364 34750
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2716 31836 2772 31892
rect 3500 31890 3556 31892
rect 3500 31838 3502 31890
rect 3502 31838 3554 31890
rect 3554 31838 3556 31890
rect 3500 31836 3556 31838
rect 6076 34188 6132 34244
rect 8540 34242 8596 34244
rect 8540 34190 8542 34242
rect 8542 34190 8594 34242
rect 8594 34190 8596 34242
rect 8540 34188 8596 34190
rect 6188 33964 6244 34020
rect 6076 31554 6132 31556
rect 6076 31502 6078 31554
rect 6078 31502 6130 31554
rect 6130 31502 6132 31554
rect 6076 31500 6132 31502
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 2380 30380 2436 30436
rect 2268 30268 2324 30324
rect 4060 30044 4116 30100
rect 4732 30156 4788 30212
rect 3052 29596 3108 29652
rect 3500 29372 3556 29428
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 2268 28028 2324 28084
rect 1932 27916 1988 27972
rect 3052 26962 3108 26964
rect 3052 26910 3054 26962
rect 3054 26910 3106 26962
rect 3106 26910 3108 26962
rect 3052 26908 3108 26910
rect 3500 28082 3556 28084
rect 3500 28030 3502 28082
rect 3502 28030 3554 28082
rect 3554 28030 3556 28082
rect 3500 28028 3556 28030
rect 3276 27970 3332 27972
rect 3276 27918 3278 27970
rect 3278 27918 3330 27970
rect 3330 27918 3332 27970
rect 3276 27916 3332 27918
rect 5068 29426 5124 29428
rect 5068 29374 5070 29426
rect 5070 29374 5122 29426
rect 5122 29374 5124 29426
rect 5068 29372 5124 29374
rect 4956 28700 5012 28756
rect 4284 28588 4340 28644
rect 4060 27804 4116 27860
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4060 27186 4116 27188
rect 4060 27134 4062 27186
rect 4062 27134 4114 27186
rect 4114 27134 4116 27186
rect 4060 27132 4116 27134
rect 5628 30828 5684 30884
rect 6188 30828 6244 30884
rect 6636 33964 6692 34020
rect 5628 30210 5684 30212
rect 5628 30158 5630 30210
rect 5630 30158 5682 30210
rect 5682 30158 5684 30210
rect 5628 30156 5684 30158
rect 6076 30044 6132 30100
rect 5628 28754 5684 28756
rect 5628 28702 5630 28754
rect 5630 28702 5682 28754
rect 5682 28702 5684 28754
rect 5628 28700 5684 28702
rect 6300 28642 6356 28644
rect 6300 28590 6302 28642
rect 6302 28590 6354 28642
rect 6354 28590 6356 28642
rect 6300 28588 6356 28590
rect 5964 28530 6020 28532
rect 5964 28478 5966 28530
rect 5966 28478 6018 28530
rect 6018 28478 6020 28530
rect 5964 28476 6020 28478
rect 5964 27916 6020 27972
rect 6076 27804 6132 27860
rect 4732 26796 4788 26852
rect 3164 26460 3220 26516
rect 3948 26460 4004 26516
rect 3052 26348 3108 26404
rect 5180 26290 5236 26292
rect 5180 26238 5182 26290
rect 5182 26238 5234 26290
rect 5234 26238 5236 26290
rect 5180 26236 5236 26238
rect 5628 26290 5684 26292
rect 5628 26238 5630 26290
rect 5630 26238 5682 26290
rect 5682 26238 5684 26290
rect 5628 26236 5684 26238
rect 7532 34018 7588 34020
rect 7532 33966 7534 34018
rect 7534 33966 7586 34018
rect 7586 33966 7588 34018
rect 7532 33964 7588 33966
rect 6748 33852 6804 33908
rect 6636 28642 6692 28644
rect 6636 28590 6638 28642
rect 6638 28590 6690 28642
rect 6690 28590 6692 28642
rect 6636 28588 6692 28590
rect 6972 32674 7028 32676
rect 6972 32622 6974 32674
rect 6974 32622 7026 32674
rect 7026 32622 7028 32674
rect 6972 32620 7028 32622
rect 7196 30882 7252 30884
rect 7196 30830 7198 30882
rect 7198 30830 7250 30882
rect 7250 30830 7252 30882
rect 7196 30828 7252 30830
rect 9996 34972 10052 35028
rect 7980 30828 8036 30884
rect 7532 29820 7588 29876
rect 8428 29820 8484 29876
rect 7196 29372 7252 29428
rect 7420 29260 7476 29316
rect 6972 28588 7028 28644
rect 8204 29650 8260 29652
rect 8204 29598 8206 29650
rect 8206 29598 8258 29650
rect 8258 29598 8260 29650
rect 8204 29596 8260 29598
rect 8316 29372 8372 29428
rect 7420 28642 7476 28644
rect 7420 28590 7422 28642
rect 7422 28590 7474 28642
rect 7474 28590 7476 28642
rect 7420 28588 7476 28590
rect 6412 26796 6468 26852
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4732 25676 4788 25732
rect 4060 25618 4116 25620
rect 4060 25566 4062 25618
rect 4062 25566 4114 25618
rect 4114 25566 4116 25618
rect 4060 25564 4116 25566
rect 4060 25228 4116 25284
rect 2044 24332 2100 24388
rect 1820 20188 1876 20244
rect 1932 19516 1988 19572
rect 1708 18508 1764 18564
rect 2492 23548 2548 23604
rect 3052 23826 3108 23828
rect 3052 23774 3054 23826
rect 3054 23774 3106 23826
rect 3106 23774 3108 23826
rect 3052 23772 3108 23774
rect 2604 23324 2660 23380
rect 2604 23154 2660 23156
rect 2604 23102 2606 23154
rect 2606 23102 2658 23154
rect 2658 23102 2660 23154
rect 2604 23100 2660 23102
rect 2828 22876 2884 22932
rect 2492 19516 2548 19572
rect 2268 19122 2324 19124
rect 2268 19070 2270 19122
rect 2270 19070 2322 19122
rect 2322 19070 2324 19122
rect 2268 19068 2324 19070
rect 2044 16940 2100 16996
rect 1596 14700 1652 14756
rect 1932 14252 1988 14308
rect 1484 12796 1540 12852
rect 1820 13468 1876 13524
rect 1596 11228 1652 11284
rect 3052 22258 3108 22260
rect 3052 22206 3054 22258
rect 3054 22206 3106 22258
rect 3106 22206 3108 22258
rect 3052 22204 3108 22206
rect 3052 20690 3108 20692
rect 3052 20638 3054 20690
rect 3054 20638 3106 20690
rect 3106 20638 3108 20690
rect 3052 20636 3108 20638
rect 3052 18172 3108 18228
rect 3500 24556 3556 24612
rect 6748 25676 6804 25732
rect 6972 26124 7028 26180
rect 8764 29314 8820 29316
rect 8764 29262 8766 29314
rect 8766 29262 8818 29314
rect 8818 29262 8820 29314
rect 8764 29260 8820 29262
rect 9212 31778 9268 31780
rect 9212 31726 9214 31778
rect 9214 31726 9266 31778
rect 9266 31726 9268 31778
rect 9212 31724 9268 31726
rect 9436 32674 9492 32676
rect 9436 32622 9438 32674
rect 9438 32622 9490 32674
rect 9490 32622 9492 32674
rect 9436 32620 9492 32622
rect 9548 31778 9604 31780
rect 9548 31726 9550 31778
rect 9550 31726 9602 31778
rect 9602 31726 9604 31778
rect 9548 31724 9604 31726
rect 9996 33292 10052 33348
rect 9996 30994 10052 30996
rect 9996 30942 9998 30994
rect 9998 30942 10050 30994
rect 10050 30942 10052 30994
rect 9996 30940 10052 30942
rect 10108 30828 10164 30884
rect 9660 29426 9716 29428
rect 9660 29374 9662 29426
rect 9662 29374 9714 29426
rect 9714 29374 9716 29426
rect 9660 29372 9716 29374
rect 10444 30882 10500 30884
rect 10444 30830 10446 30882
rect 10446 30830 10498 30882
rect 10498 30830 10500 30882
rect 10444 30828 10500 30830
rect 8652 27804 8708 27860
rect 8540 26514 8596 26516
rect 8540 26462 8542 26514
rect 8542 26462 8594 26514
rect 8594 26462 8596 26514
rect 8540 26460 8596 26462
rect 7980 26236 8036 26292
rect 5964 24556 6020 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3612 23548 3668 23604
rect 3500 23324 3556 23380
rect 3388 18508 3444 18564
rect 6860 24108 6916 24164
rect 6636 23660 6692 23716
rect 5516 23100 5572 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4060 22482 4116 22484
rect 4060 22430 4062 22482
rect 4062 22430 4114 22482
rect 4114 22430 4116 22482
rect 4060 22428 4116 22430
rect 3836 21868 3892 21924
rect 3836 20524 3892 20580
rect 3948 19292 4004 19348
rect 3500 17500 3556 17556
rect 6076 22930 6132 22932
rect 6076 22878 6078 22930
rect 6078 22878 6130 22930
rect 6130 22878 6132 22930
rect 6076 22876 6132 22878
rect 6748 22652 6804 22708
rect 5404 21420 5460 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 6076 22092 6132 22148
rect 6636 21474 6692 21476
rect 6636 21422 6638 21474
rect 6638 21422 6690 21474
rect 6690 21422 6692 21474
rect 6636 21420 6692 21422
rect 5964 19292 6020 19348
rect 6076 19628 6132 19684
rect 5964 19068 6020 19124
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 2716 14306 2772 14308
rect 2716 14254 2718 14306
rect 2718 14254 2770 14306
rect 2770 14254 2772 14306
rect 2716 14252 2772 14254
rect 2380 13916 2436 13972
rect 2380 12850 2436 12852
rect 2380 12798 2382 12850
rect 2382 12798 2434 12850
rect 2434 12798 2436 12850
rect 2380 12796 2436 12798
rect 2604 12572 2660 12628
rect 2044 11900 2100 11956
rect 2380 11282 2436 11284
rect 2380 11230 2382 11282
rect 2382 11230 2434 11282
rect 2434 11230 2436 11282
rect 2380 11228 2436 11230
rect 3164 14306 3220 14308
rect 3164 14254 3166 14306
rect 3166 14254 3218 14306
rect 3218 14254 3220 14306
rect 3164 14252 3220 14254
rect 3164 13580 3220 13636
rect 3500 12572 3556 12628
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5404 18226 5460 18228
rect 5404 18174 5406 18226
rect 5406 18174 5458 18226
rect 5458 18174 5460 18226
rect 5404 18172 5460 18174
rect 4844 16268 4900 16324
rect 4956 16828 5012 16884
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 6748 19628 6804 19684
rect 7644 24722 7700 24724
rect 7644 24670 7646 24722
rect 7646 24670 7698 24722
rect 7698 24670 7700 24722
rect 7644 24668 7700 24670
rect 8540 25676 8596 25732
rect 9884 28364 9940 28420
rect 11004 30828 11060 30884
rect 11452 33292 11508 33348
rect 12124 30994 12180 30996
rect 12124 30942 12126 30994
rect 12126 30942 12178 30994
rect 12178 30942 12180 30994
rect 12124 30940 12180 30942
rect 11452 30882 11508 30884
rect 11452 30830 11454 30882
rect 11454 30830 11506 30882
rect 11506 30830 11508 30882
rect 11452 30828 11508 30830
rect 10892 30716 10948 30772
rect 11676 29596 11732 29652
rect 11788 30716 11844 30772
rect 10444 28364 10500 28420
rect 11228 28588 11284 28644
rect 12012 28642 12068 28644
rect 12012 28590 12014 28642
rect 12014 28590 12066 28642
rect 12066 28590 12068 28642
rect 12012 28588 12068 28590
rect 12236 30828 12292 30884
rect 12348 30156 12404 30212
rect 12460 30044 12516 30100
rect 13804 37378 13860 37380
rect 13804 37326 13806 37378
rect 13806 37326 13858 37378
rect 13858 37326 13860 37378
rect 13804 37324 13860 37326
rect 13244 34300 13300 34356
rect 13468 33292 13524 33348
rect 13356 30940 13412 30996
rect 14028 35196 14084 35252
rect 14028 30604 14084 30660
rect 13468 30098 13524 30100
rect 13468 30046 13470 30098
rect 13470 30046 13522 30098
rect 13522 30046 13524 30098
rect 13468 30044 13524 30046
rect 12348 29650 12404 29652
rect 12348 29598 12350 29650
rect 12350 29598 12402 29650
rect 12402 29598 12404 29650
rect 12348 29596 12404 29598
rect 12124 28476 12180 28532
rect 10108 27858 10164 27860
rect 10108 27806 10110 27858
rect 10110 27806 10162 27858
rect 10162 27806 10164 27858
rect 10108 27804 10164 27806
rect 9772 27132 9828 27188
rect 9660 26514 9716 26516
rect 9660 26462 9662 26514
rect 9662 26462 9714 26514
rect 9714 26462 9716 26514
rect 9660 26460 9716 26462
rect 9660 26236 9716 26292
rect 9548 26178 9604 26180
rect 9548 26126 9550 26178
rect 9550 26126 9602 26178
rect 9602 26126 9604 26178
rect 9548 26124 9604 26126
rect 7980 24668 8036 24724
rect 8988 25676 9044 25732
rect 7868 23884 7924 23940
rect 8428 22146 8484 22148
rect 8428 22094 8430 22146
rect 8430 22094 8482 22146
rect 8482 22094 8484 22146
rect 8428 22092 8484 22094
rect 6972 20524 7028 20580
rect 7756 21980 7812 22036
rect 7644 19964 7700 20020
rect 6636 17388 6692 17444
rect 6972 16604 7028 16660
rect 6300 15874 6356 15876
rect 6300 15822 6302 15874
rect 6302 15822 6354 15874
rect 6354 15822 6356 15874
rect 6300 15820 6356 15822
rect 5068 15314 5124 15316
rect 5068 15262 5070 15314
rect 5070 15262 5122 15314
rect 5122 15262 5124 15314
rect 5068 15260 5124 15262
rect 4844 13970 4900 13972
rect 4844 13918 4846 13970
rect 4846 13918 4898 13970
rect 4898 13918 4900 13970
rect 4844 13916 4900 13918
rect 5740 15260 5796 15316
rect 5068 13468 5124 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4396 13132 4452 13188
rect 5852 13634 5908 13636
rect 5852 13582 5854 13634
rect 5854 13582 5906 13634
rect 5906 13582 5908 13634
rect 5852 13580 5908 13582
rect 5628 13020 5684 13076
rect 5516 12572 5572 12628
rect 4284 11900 4340 11956
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 6524 14700 6580 14756
rect 9324 24668 9380 24724
rect 11676 26962 11732 26964
rect 11676 26910 11678 26962
rect 11678 26910 11730 26962
rect 11730 26910 11732 26962
rect 11676 26908 11732 26910
rect 9884 25506 9940 25508
rect 9884 25454 9886 25506
rect 9886 25454 9938 25506
rect 9938 25454 9940 25506
rect 9884 25452 9940 25454
rect 10108 24108 10164 24164
rect 8876 22988 8932 23044
rect 9660 23042 9716 23044
rect 9660 22990 9662 23042
rect 9662 22990 9714 23042
rect 9714 22990 9716 23042
rect 9660 22988 9716 22990
rect 9212 22146 9268 22148
rect 9212 22094 9214 22146
rect 9214 22094 9266 22146
rect 9266 22094 9268 22146
rect 9212 22092 9268 22094
rect 8316 21420 8372 21476
rect 7980 18508 8036 18564
rect 9548 21532 9604 21588
rect 9324 20690 9380 20692
rect 9324 20638 9326 20690
rect 9326 20638 9378 20690
rect 9378 20638 9380 20690
rect 9324 20636 9380 20638
rect 8540 20018 8596 20020
rect 8540 19966 8542 20018
rect 8542 19966 8594 20018
rect 8594 19966 8596 20018
rect 8540 19964 8596 19966
rect 8092 17612 8148 17668
rect 8204 18844 8260 18900
rect 8652 17948 8708 18004
rect 8540 16098 8596 16100
rect 8540 16046 8542 16098
rect 8542 16046 8594 16098
rect 8594 16046 8596 16098
rect 8540 16044 8596 16046
rect 8316 15484 8372 15540
rect 7980 15148 8036 15204
rect 7868 15036 7924 15092
rect 7756 13356 7812 13412
rect 6972 13132 7028 13188
rect 6748 12572 6804 12628
rect 9212 18620 9268 18676
rect 9436 18508 9492 18564
rect 8988 17052 9044 17108
rect 9212 17666 9268 17668
rect 9212 17614 9214 17666
rect 9214 17614 9266 17666
rect 9266 17614 9268 17666
rect 9212 17612 9268 17614
rect 9100 16658 9156 16660
rect 9100 16606 9102 16658
rect 9102 16606 9154 16658
rect 9154 16606 9156 16658
rect 9100 16604 9156 16606
rect 8876 15148 8932 15204
rect 8428 14812 8484 14868
rect 8428 13634 8484 13636
rect 8428 13582 8430 13634
rect 8430 13582 8482 13634
rect 8482 13582 8484 13634
rect 8428 13580 8484 13582
rect 8988 15036 9044 15092
rect 9436 16828 9492 16884
rect 9212 16044 9268 16100
rect 9212 15484 9268 15540
rect 8764 13356 8820 13412
rect 9548 15426 9604 15428
rect 9548 15374 9550 15426
rect 9550 15374 9602 15426
rect 9602 15374 9604 15426
rect 9548 15372 9604 15374
rect 9436 13356 9492 13412
rect 12236 28700 12292 28756
rect 12236 28364 12292 28420
rect 12908 27804 12964 27860
rect 14252 30210 14308 30212
rect 14252 30158 14254 30210
rect 14254 30158 14306 30210
rect 14306 30158 14308 30210
rect 14252 30156 14308 30158
rect 15148 35196 15204 35252
rect 14700 35026 14756 35028
rect 14700 34974 14702 35026
rect 14702 34974 14754 35026
rect 14754 34974 14756 35026
rect 14700 34972 14756 34974
rect 15820 34300 15876 34356
rect 15596 33740 15652 33796
rect 15484 31612 15540 31668
rect 13692 28700 13748 28756
rect 14588 30098 14644 30100
rect 14588 30046 14590 30098
rect 14590 30046 14642 30098
rect 14642 30046 14644 30098
rect 14588 30044 14644 30046
rect 13356 28588 13412 28644
rect 13580 28476 13636 28532
rect 13468 27804 13524 27860
rect 14028 28754 14084 28756
rect 14028 28702 14030 28754
rect 14030 28702 14082 28754
rect 14082 28702 14084 28754
rect 14028 28700 14084 28702
rect 15260 30098 15316 30100
rect 15260 30046 15262 30098
rect 15262 30046 15314 30098
rect 15314 30046 15316 30098
rect 15260 30044 15316 30046
rect 14476 28754 14532 28756
rect 14476 28702 14478 28754
rect 14478 28702 14530 28754
rect 14530 28702 14532 28754
rect 14476 28700 14532 28702
rect 15148 28642 15204 28644
rect 15148 28590 15150 28642
rect 15150 28590 15202 28642
rect 15202 28590 15204 28642
rect 15148 28588 15204 28590
rect 14924 28476 14980 28532
rect 13468 27074 13524 27076
rect 13468 27022 13470 27074
rect 13470 27022 13522 27074
rect 13522 27022 13524 27074
rect 13468 27020 13524 27022
rect 11788 26290 11844 26292
rect 11788 26238 11790 26290
rect 11790 26238 11842 26290
rect 11842 26238 11844 26290
rect 11788 26236 11844 26238
rect 12348 25564 12404 25620
rect 11564 25452 11620 25508
rect 9884 21868 9940 21924
rect 12236 25228 12292 25284
rect 13020 26348 13076 26404
rect 13244 26236 13300 26292
rect 12908 25452 12964 25508
rect 12572 25340 12628 25396
rect 13692 25506 13748 25508
rect 13692 25454 13694 25506
rect 13694 25454 13746 25506
rect 13746 25454 13748 25506
rect 13692 25452 13748 25454
rect 14364 25506 14420 25508
rect 14364 25454 14366 25506
rect 14366 25454 14418 25506
rect 14418 25454 14420 25506
rect 14364 25452 14420 25454
rect 13468 25394 13524 25396
rect 13468 25342 13470 25394
rect 13470 25342 13522 25394
rect 13522 25342 13524 25394
rect 13468 25340 13524 25342
rect 14140 25228 14196 25284
rect 13132 23772 13188 23828
rect 12572 22988 12628 23044
rect 11564 22092 11620 22148
rect 11676 22876 11732 22932
rect 9884 21420 9940 21476
rect 10556 21474 10612 21476
rect 10556 21422 10558 21474
rect 10558 21422 10610 21474
rect 10610 21422 10612 21474
rect 10556 21420 10612 21422
rect 15820 31724 15876 31780
rect 16044 33628 16100 33684
rect 16380 35196 16436 35252
rect 16604 34690 16660 34692
rect 16604 34638 16606 34690
rect 16606 34638 16658 34690
rect 16658 34638 16660 34690
rect 16604 34636 16660 34638
rect 16828 33628 16884 33684
rect 16492 32284 16548 32340
rect 18844 37938 18900 37940
rect 18844 37886 18846 37938
rect 18846 37886 18898 37938
rect 18898 37886 18900 37938
rect 18844 37884 18900 37886
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 17836 35196 17892 35252
rect 17276 33516 17332 33572
rect 16156 30044 16212 30100
rect 16828 30044 16884 30100
rect 15932 29932 15988 29988
rect 16268 29708 16324 29764
rect 16380 29650 16436 29652
rect 16380 29598 16382 29650
rect 16382 29598 16434 29650
rect 16434 29598 16436 29650
rect 16380 29596 16436 29598
rect 17500 33292 17556 33348
rect 17388 32284 17444 32340
rect 17948 34636 18004 34692
rect 17612 31724 17668 31780
rect 18396 34018 18452 34020
rect 18396 33966 18398 34018
rect 18398 33966 18450 34018
rect 18450 33966 18452 34018
rect 18396 33964 18452 33966
rect 17164 30156 17220 30212
rect 16940 29372 16996 29428
rect 17388 30604 17444 30660
rect 18060 32060 18116 32116
rect 17836 31836 17892 31892
rect 17612 30044 17668 30100
rect 17164 28588 17220 28644
rect 18396 30716 18452 30772
rect 18172 29708 18228 29764
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 19516 33740 19572 33796
rect 21196 36316 21252 36372
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 34242 19796 34244
rect 19740 34190 19742 34242
rect 19742 34190 19794 34242
rect 19794 34190 19796 34242
rect 19740 34188 19796 34190
rect 19628 33516 19684 33572
rect 18732 31836 18788 31892
rect 18732 30716 18788 30772
rect 18284 29372 18340 29428
rect 18284 28476 18340 28532
rect 17388 27020 17444 27076
rect 17052 26460 17108 26516
rect 17500 26796 17556 26852
rect 19068 30210 19124 30212
rect 19068 30158 19070 30210
rect 19070 30158 19122 30210
rect 19122 30158 19124 30210
rect 19068 30156 19124 30158
rect 18396 27916 18452 27972
rect 18284 26796 18340 26852
rect 18844 26460 18900 26516
rect 15484 26236 15540 26292
rect 15372 24892 15428 24948
rect 14924 24444 14980 24500
rect 15148 23996 15204 24052
rect 14028 23884 14084 23940
rect 13916 23436 13972 23492
rect 15260 23436 15316 23492
rect 13132 22930 13188 22932
rect 13132 22878 13134 22930
rect 13134 22878 13186 22930
rect 13186 22878 13188 22930
rect 13132 22876 13188 22878
rect 12796 22652 12852 22708
rect 12572 22316 12628 22372
rect 12684 22428 12740 22484
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 13804 22370 13860 22372
rect 13804 22318 13806 22370
rect 13806 22318 13858 22370
rect 13858 22318 13860 22370
rect 13804 22316 13860 22318
rect 13020 22258 13076 22260
rect 13020 22206 13022 22258
rect 13022 22206 13074 22258
rect 13074 22206 13076 22258
rect 13020 22204 13076 22206
rect 13356 21756 13412 21812
rect 15036 22204 15092 22260
rect 14476 22146 14532 22148
rect 14476 22094 14478 22146
rect 14478 22094 14530 22146
rect 14530 22094 14532 22146
rect 14476 22092 14532 22094
rect 13916 21644 13972 21700
rect 10220 19852 10276 19908
rect 10668 19964 10724 20020
rect 9884 17948 9940 18004
rect 10220 17612 10276 17668
rect 9772 17388 9828 17444
rect 8652 12460 8708 12516
rect 9324 13020 9380 13076
rect 10108 17052 10164 17108
rect 9996 15484 10052 15540
rect 9884 15202 9940 15204
rect 9884 15150 9886 15202
rect 9886 15150 9938 15202
rect 9938 15150 9940 15202
rect 9884 15148 9940 15150
rect 9884 14812 9940 14868
rect 10220 16994 10276 16996
rect 10220 16942 10222 16994
rect 10222 16942 10274 16994
rect 10274 16942 10276 16994
rect 10220 16940 10276 16942
rect 10444 16268 10500 16324
rect 10332 15538 10388 15540
rect 10332 15486 10334 15538
rect 10334 15486 10386 15538
rect 10386 15486 10388 15538
rect 10332 15484 10388 15486
rect 11452 19068 11508 19124
rect 11228 18620 11284 18676
rect 10668 16828 10724 16884
rect 9660 12012 9716 12068
rect 10556 12460 10612 12516
rect 10780 15202 10836 15204
rect 10780 15150 10782 15202
rect 10782 15150 10834 15202
rect 10834 15150 10836 15202
rect 10780 15148 10836 15150
rect 11452 17500 11508 17556
rect 12460 20018 12516 20020
rect 12460 19966 12462 20018
rect 12462 19966 12514 20018
rect 12514 19966 12516 20018
rect 12460 19964 12516 19966
rect 12236 19122 12292 19124
rect 12236 19070 12238 19122
rect 12238 19070 12290 19122
rect 12290 19070 12292 19122
rect 12236 19068 12292 19070
rect 12572 19122 12628 19124
rect 12572 19070 12574 19122
rect 12574 19070 12626 19122
rect 12626 19070 12628 19122
rect 12572 19068 12628 19070
rect 12124 18508 12180 18564
rect 12460 16882 12516 16884
rect 12460 16830 12462 16882
rect 12462 16830 12514 16882
rect 12514 16830 12516 16882
rect 12460 16828 12516 16830
rect 11788 13356 11844 13412
rect 12348 15874 12404 15876
rect 12348 15822 12350 15874
rect 12350 15822 12402 15874
rect 12402 15822 12404 15874
rect 12348 15820 12404 15822
rect 12348 15148 12404 15204
rect 12684 15596 12740 15652
rect 13468 18508 13524 18564
rect 13692 19068 13748 19124
rect 13020 17388 13076 17444
rect 13468 17612 13524 17668
rect 14140 19122 14196 19124
rect 14140 19070 14142 19122
rect 14142 19070 14194 19122
rect 14194 19070 14196 19122
rect 14140 19068 14196 19070
rect 13580 17554 13636 17556
rect 13580 17502 13582 17554
rect 13582 17502 13634 17554
rect 13634 17502 13636 17554
rect 13580 17500 13636 17502
rect 12908 15874 12964 15876
rect 12908 15822 12910 15874
rect 12910 15822 12962 15874
rect 12962 15822 12964 15874
rect 12908 15820 12964 15822
rect 13692 16716 13748 16772
rect 14140 16828 14196 16884
rect 14028 16156 14084 16212
rect 13692 15820 13748 15876
rect 14028 15874 14084 15876
rect 14028 15822 14030 15874
rect 14030 15822 14082 15874
rect 14082 15822 14084 15874
rect 14028 15820 14084 15822
rect 13020 15484 13076 15540
rect 13580 15596 13636 15652
rect 14812 19404 14868 19460
rect 14364 19234 14420 19236
rect 14364 19182 14366 19234
rect 14366 19182 14418 19234
rect 14418 19182 14420 19234
rect 14364 19180 14420 19182
rect 14364 17442 14420 17444
rect 14364 17390 14366 17442
rect 14366 17390 14418 17442
rect 14418 17390 14420 17442
rect 14364 17388 14420 17390
rect 14924 19234 14980 19236
rect 14924 19182 14926 19234
rect 14926 19182 14978 19234
rect 14978 19182 14980 19234
rect 14924 19180 14980 19182
rect 14924 17612 14980 17668
rect 14812 16716 14868 16772
rect 14588 16044 14644 16100
rect 15820 25452 15876 25508
rect 16828 26178 16884 26180
rect 16828 26126 16830 26178
rect 16830 26126 16882 26178
rect 16882 26126 16884 26178
rect 16828 26124 16884 26126
rect 17948 26178 18004 26180
rect 17948 26126 17950 26178
rect 17950 26126 18002 26178
rect 18002 26126 18004 26178
rect 17948 26124 18004 26126
rect 18620 26124 18676 26180
rect 17500 24722 17556 24724
rect 17500 24670 17502 24722
rect 17502 24670 17554 24722
rect 17554 24670 17556 24722
rect 17500 24668 17556 24670
rect 16380 24332 16436 24388
rect 16268 23714 16324 23716
rect 16268 23662 16270 23714
rect 16270 23662 16322 23714
rect 16322 23662 16324 23714
rect 16268 23660 16324 23662
rect 17052 23714 17108 23716
rect 17052 23662 17054 23714
rect 17054 23662 17106 23714
rect 17106 23662 17108 23714
rect 17052 23660 17108 23662
rect 15820 19404 15876 19460
rect 16380 22258 16436 22260
rect 16380 22206 16382 22258
rect 16382 22206 16434 22258
rect 16434 22206 16436 22258
rect 16380 22204 16436 22206
rect 16380 21698 16436 21700
rect 16380 21646 16382 21698
rect 16382 21646 16434 21698
rect 16434 21646 16436 21698
rect 16380 21644 16436 21646
rect 15708 18284 15764 18340
rect 15148 16828 15204 16884
rect 15036 16268 15092 16324
rect 15484 16156 15540 16212
rect 15260 16098 15316 16100
rect 15260 16046 15262 16098
rect 15262 16046 15314 16098
rect 15314 16046 15316 16098
rect 15260 16044 15316 16046
rect 14364 13020 14420 13076
rect 15932 19010 15988 19012
rect 15932 18958 15934 19010
rect 15934 18958 15986 19010
rect 15986 18958 15988 19010
rect 15932 18956 15988 18958
rect 16380 19292 16436 19348
rect 16268 18396 16324 18452
rect 16716 22988 16772 23044
rect 16716 22092 16772 22148
rect 17164 21868 17220 21924
rect 16716 18284 16772 18340
rect 16380 17052 16436 17108
rect 16268 16380 16324 16436
rect 16940 17666 16996 17668
rect 16940 17614 16942 17666
rect 16942 17614 16994 17666
rect 16994 17614 16996 17666
rect 16940 17612 16996 17614
rect 16828 16268 16884 16324
rect 17164 15484 17220 15540
rect 17500 24444 17556 24500
rect 17836 24220 17892 24276
rect 17388 23042 17444 23044
rect 17388 22990 17390 23042
rect 17390 22990 17442 23042
rect 17442 22990 17444 23042
rect 17388 22988 17444 22990
rect 18060 22988 18116 23044
rect 17724 21980 17780 22036
rect 17948 20748 18004 20804
rect 18172 21980 18228 22036
rect 18508 21868 18564 21924
rect 17836 20018 17892 20020
rect 17836 19966 17838 20018
rect 17838 19966 17890 20018
rect 17890 19966 17892 20018
rect 17836 19964 17892 19966
rect 17836 18450 17892 18452
rect 17836 18398 17838 18450
rect 17838 18398 17890 18450
rect 17890 18398 17892 18450
rect 17836 18396 17892 18398
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 17724 17052 17780 17108
rect 18284 17164 18340 17220
rect 19068 29596 19124 29652
rect 19068 27916 19124 27972
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20636 34972 20692 35028
rect 20860 31948 20916 32004
rect 22316 35026 22372 35028
rect 22316 34974 22318 35026
rect 22318 34974 22370 35026
rect 22370 34974 22372 35026
rect 22316 34972 22372 34974
rect 21308 34524 21364 34580
rect 23548 36370 23604 36372
rect 23548 36318 23550 36370
rect 23550 36318 23602 36370
rect 23602 36318 23604 36370
rect 23548 36316 23604 36318
rect 22428 34524 22484 34580
rect 21532 32060 21588 32116
rect 21644 33068 21700 33124
rect 20636 30156 20692 30212
rect 20748 30098 20804 30100
rect 20748 30046 20750 30098
rect 20750 30046 20802 30098
rect 20802 30046 20804 30098
rect 20748 30044 20804 30046
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 27916 19796 27972
rect 19740 26908 19796 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20524 28812 20580 28868
rect 20748 28642 20804 28644
rect 20748 28590 20750 28642
rect 20750 28590 20802 28642
rect 20802 28590 20804 28642
rect 20748 28588 20804 28590
rect 19068 26124 19124 26180
rect 20300 25228 20356 25284
rect 21756 32956 21812 33012
rect 21644 30044 21700 30100
rect 21644 28812 21700 28868
rect 21532 28700 21588 28756
rect 21196 26908 21252 26964
rect 20748 25282 20804 25284
rect 20748 25230 20750 25282
rect 20750 25230 20802 25282
rect 20802 25230 20804 25282
rect 20748 25228 20804 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19964 24668 20020 24724
rect 18620 18396 18676 18452
rect 18060 16994 18116 16996
rect 18060 16942 18062 16994
rect 18062 16942 18114 16994
rect 18114 16942 18116 16994
rect 18060 16940 18116 16942
rect 17500 16380 17556 16436
rect 17836 15932 17892 15988
rect 16828 13916 16884 13972
rect 18620 15986 18676 15988
rect 18620 15934 18622 15986
rect 18622 15934 18674 15986
rect 18674 15934 18676 15986
rect 18620 15932 18676 15934
rect 20188 24332 20244 24388
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19404 23266 19460 23268
rect 19404 23214 19406 23266
rect 19406 23214 19458 23266
rect 19458 23214 19460 23266
rect 19404 23212 19460 23214
rect 19068 23042 19124 23044
rect 19068 22990 19070 23042
rect 19070 22990 19122 23042
rect 19122 22990 19124 23042
rect 19068 22988 19124 22990
rect 19404 22204 19460 22260
rect 18844 18620 18900 18676
rect 19180 18956 19236 19012
rect 20972 24946 21028 24948
rect 20972 24894 20974 24946
rect 20974 24894 21026 24946
rect 21026 24894 21028 24946
rect 20972 24892 21028 24894
rect 22764 31948 22820 32004
rect 23212 33180 23268 33236
rect 22204 31388 22260 31444
rect 21980 29986 22036 29988
rect 21980 29934 21982 29986
rect 21982 29934 22034 29986
rect 22034 29934 22036 29986
rect 21980 29932 22036 29934
rect 22764 29986 22820 29988
rect 22764 29934 22766 29986
rect 22766 29934 22818 29986
rect 22818 29934 22820 29986
rect 22764 29932 22820 29934
rect 22652 27244 22708 27300
rect 23324 33068 23380 33124
rect 23548 31388 23604 31444
rect 34636 35420 34692 35476
rect 24332 34748 24388 34804
rect 24220 31052 24276 31108
rect 23772 30828 23828 30884
rect 24892 33068 24948 33124
rect 24780 31778 24836 31780
rect 24780 31726 24782 31778
rect 24782 31726 24834 31778
rect 24834 31726 24836 31778
rect 24780 31724 24836 31726
rect 26124 34802 26180 34804
rect 26124 34750 26126 34802
rect 26126 34750 26178 34802
rect 26178 34750 26180 34802
rect 26124 34748 26180 34750
rect 25788 33292 25844 33348
rect 25676 33234 25732 33236
rect 25676 33182 25678 33234
rect 25678 33182 25730 33234
rect 25730 33182 25732 33234
rect 25676 33180 25732 33182
rect 25116 32956 25172 33012
rect 25116 31836 25172 31892
rect 23772 28476 23828 28532
rect 23660 27804 23716 27860
rect 25228 31778 25284 31780
rect 25228 31726 25230 31778
rect 25230 31726 25282 31778
rect 25282 31726 25284 31778
rect 25228 31724 25284 31726
rect 28924 34188 28980 34244
rect 27244 33068 27300 33124
rect 26236 31836 26292 31892
rect 26012 31724 26068 31780
rect 25228 31106 25284 31108
rect 25228 31054 25230 31106
rect 25230 31054 25282 31106
rect 25282 31054 25284 31106
rect 25228 31052 25284 31054
rect 26572 31724 26628 31780
rect 25228 30828 25284 30884
rect 24892 30044 24948 30100
rect 24444 28812 24500 28868
rect 24220 28754 24276 28756
rect 24220 28702 24222 28754
rect 24222 28702 24274 28754
rect 24274 28702 24276 28754
rect 24220 28700 24276 28702
rect 24108 27692 24164 27748
rect 25676 30210 25732 30212
rect 25676 30158 25678 30210
rect 25678 30158 25730 30210
rect 25730 30158 25732 30210
rect 25676 30156 25732 30158
rect 26684 30994 26740 30996
rect 26684 30942 26686 30994
rect 26686 30942 26738 30994
rect 26738 30942 26740 30994
rect 26684 30940 26740 30942
rect 28700 33180 28756 33236
rect 28252 32508 28308 32564
rect 28140 32396 28196 32452
rect 27244 30828 27300 30884
rect 26012 30156 26068 30212
rect 26012 29932 26068 29988
rect 25452 28812 25508 28868
rect 25004 28476 25060 28532
rect 26572 28642 26628 28644
rect 26572 28590 26574 28642
rect 26574 28590 26626 28642
rect 26626 28590 26628 28642
rect 26572 28588 26628 28590
rect 25228 27746 25284 27748
rect 25228 27694 25230 27746
rect 25230 27694 25282 27746
rect 25282 27694 25284 27746
rect 25228 27692 25284 27694
rect 25004 27580 25060 27636
rect 25004 27298 25060 27300
rect 25004 27246 25006 27298
rect 25006 27246 25058 27298
rect 25058 27246 25060 27298
rect 25004 27244 25060 27246
rect 24444 27132 24500 27188
rect 25116 27132 25172 27188
rect 25004 26908 25060 26964
rect 22204 26236 22260 26292
rect 22092 24892 22148 24948
rect 21196 24722 21252 24724
rect 21196 24670 21198 24722
rect 21198 24670 21250 24722
rect 21250 24670 21252 24722
rect 21196 24668 21252 24670
rect 21644 23996 21700 24052
rect 23100 26236 23156 26292
rect 23660 25116 23716 25172
rect 22204 24050 22260 24052
rect 22204 23998 22206 24050
rect 22206 23998 22258 24050
rect 22258 23998 22260 24050
rect 22204 23996 22260 23998
rect 23324 23996 23380 24052
rect 23212 23884 23268 23940
rect 20748 23826 20804 23828
rect 20748 23774 20750 23826
rect 20750 23774 20802 23826
rect 20802 23774 20804 23826
rect 20748 23772 20804 23774
rect 21308 23660 21364 23716
rect 21644 23826 21700 23828
rect 21644 23774 21646 23826
rect 21646 23774 21698 23826
rect 21698 23774 21700 23826
rect 21644 23772 21700 23774
rect 20748 23212 20804 23268
rect 21196 22988 21252 23044
rect 19628 21868 19684 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19852 19292 19908 19348
rect 18956 18338 19012 18340
rect 18956 18286 18958 18338
rect 18958 18286 19010 18338
rect 19010 18286 19012 18338
rect 18956 18284 19012 18286
rect 19180 17612 19236 17668
rect 19068 17164 19124 17220
rect 18956 16940 19012 16996
rect 18396 13916 18452 13972
rect 12012 12066 12068 12068
rect 12012 12014 12014 12066
rect 12014 12014 12066 12066
rect 12066 12014 12068 12066
rect 12012 12012 12068 12014
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18396 19684 18452
rect 19852 18284 19908 18340
rect 20300 20524 20356 20580
rect 20412 20748 20468 20804
rect 20300 19516 20356 19572
rect 21420 22370 21476 22372
rect 21420 22318 21422 22370
rect 21422 22318 21474 22370
rect 21474 22318 21476 22370
rect 21420 22316 21476 22318
rect 21532 20914 21588 20916
rect 21532 20862 21534 20914
rect 21534 20862 21586 20914
rect 21586 20862 21588 20914
rect 21532 20860 21588 20862
rect 20748 19516 20804 19572
rect 20860 19964 20916 20020
rect 21420 20524 21476 20580
rect 20300 18620 20356 18676
rect 20524 18956 20580 19012
rect 20188 17612 20244 17668
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19740 15484 19796 15540
rect 20300 15148 20356 15204
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19292 13074 19348 13076
rect 19292 13022 19294 13074
rect 19294 13022 19346 13074
rect 19346 13022 19348 13074
rect 19292 13020 19348 13022
rect 20860 18396 20916 18452
rect 22428 23826 22484 23828
rect 22428 23774 22430 23826
rect 22430 23774 22482 23826
rect 22482 23774 22484 23826
rect 22428 23772 22484 23774
rect 23660 23548 23716 23604
rect 23548 23042 23604 23044
rect 23548 22990 23550 23042
rect 23550 22990 23602 23042
rect 23602 22990 23604 23042
rect 23548 22988 23604 22990
rect 21868 22204 21924 22260
rect 23436 21586 23492 21588
rect 23436 21534 23438 21586
rect 23438 21534 23490 21586
rect 23490 21534 23492 21586
rect 23436 21532 23492 21534
rect 24556 25506 24612 25508
rect 24556 25454 24558 25506
rect 24558 25454 24610 25506
rect 24610 25454 24612 25506
rect 24556 25452 24612 25454
rect 28140 30156 28196 30212
rect 27916 30098 27972 30100
rect 27916 30046 27918 30098
rect 27918 30046 27970 30098
rect 27970 30046 27972 30098
rect 27916 30044 27972 30046
rect 27580 29538 27636 29540
rect 27580 29486 27582 29538
rect 27582 29486 27634 29538
rect 27634 29486 27636 29538
rect 27580 29484 27636 29486
rect 27020 28588 27076 28644
rect 27132 28700 27188 28756
rect 27356 28028 27412 28084
rect 27468 27858 27524 27860
rect 27468 27806 27470 27858
rect 27470 27806 27522 27858
rect 27522 27806 27524 27858
rect 27468 27804 27524 27806
rect 26796 26908 26852 26964
rect 27580 27132 27636 27188
rect 25676 26290 25732 26292
rect 25676 26238 25678 26290
rect 25678 26238 25730 26290
rect 25730 26238 25732 26290
rect 25676 26236 25732 26238
rect 25116 25452 25172 25508
rect 25676 25452 25732 25508
rect 24780 24946 24836 24948
rect 24780 24894 24782 24946
rect 24782 24894 24834 24946
rect 24834 24894 24836 24946
rect 24780 24892 24836 24894
rect 23884 23772 23940 23828
rect 24332 23548 24388 23604
rect 23884 23266 23940 23268
rect 23884 23214 23886 23266
rect 23886 23214 23938 23266
rect 23938 23214 23940 23266
rect 23884 23212 23940 23214
rect 24556 23212 24612 23268
rect 24444 22316 24500 22372
rect 23884 20860 23940 20916
rect 23660 20802 23716 20804
rect 23660 20750 23662 20802
rect 23662 20750 23714 20802
rect 23714 20750 23716 20802
rect 23660 20748 23716 20750
rect 26012 25340 26068 25396
rect 26348 23996 26404 24052
rect 26572 24108 26628 24164
rect 27244 24108 27300 24164
rect 26796 23548 26852 23604
rect 26012 23266 26068 23268
rect 26012 23214 26014 23266
rect 26014 23214 26066 23266
rect 26066 23214 26068 23266
rect 26012 23212 26068 23214
rect 26684 23154 26740 23156
rect 26684 23102 26686 23154
rect 26686 23102 26738 23154
rect 26738 23102 26740 23154
rect 26684 23100 26740 23102
rect 25004 22370 25060 22372
rect 25004 22318 25006 22370
rect 25006 22318 25058 22370
rect 25058 22318 25060 22370
rect 25004 22316 25060 22318
rect 24892 22146 24948 22148
rect 24892 22094 24894 22146
rect 24894 22094 24946 22146
rect 24946 22094 24948 22146
rect 24892 22092 24948 22094
rect 25340 21644 25396 21700
rect 25676 21196 25732 21252
rect 25788 21644 25844 21700
rect 21084 17612 21140 17668
rect 23100 19852 23156 19908
rect 22316 19010 22372 19012
rect 22316 18958 22318 19010
rect 22318 18958 22370 19010
rect 22370 18958 22372 19010
rect 22316 18956 22372 18958
rect 22540 18396 22596 18452
rect 21868 17778 21924 17780
rect 21868 17726 21870 17778
rect 21870 17726 21922 17778
rect 21922 17726 21924 17778
rect 21868 17724 21924 17726
rect 23660 18450 23716 18452
rect 23660 18398 23662 18450
rect 23662 18398 23714 18450
rect 23714 18398 23716 18450
rect 23660 18396 23716 18398
rect 24332 18450 24388 18452
rect 24332 18398 24334 18450
rect 24334 18398 24386 18450
rect 24386 18398 24388 18450
rect 24332 18396 24388 18398
rect 22540 17778 22596 17780
rect 22540 17726 22542 17778
rect 22542 17726 22594 17778
rect 22594 17726 22596 17778
rect 22540 17724 22596 17726
rect 22764 17666 22820 17668
rect 22764 17614 22766 17666
rect 22766 17614 22818 17666
rect 22818 17614 22820 17666
rect 22764 17612 22820 17614
rect 21532 17500 21588 17556
rect 21756 15932 21812 15988
rect 22428 17500 22484 17556
rect 20860 13580 20916 13636
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 22876 16604 22932 16660
rect 22652 15932 22708 15988
rect 23436 15820 23492 15876
rect 23660 16604 23716 16660
rect 23996 16044 24052 16100
rect 22876 15036 22932 15092
rect 22988 13580 23044 13636
rect 23884 15090 23940 15092
rect 23884 15038 23886 15090
rect 23886 15038 23938 15090
rect 23938 15038 23940 15090
rect 23884 15036 23940 15038
rect 23884 14588 23940 14644
rect 25228 19906 25284 19908
rect 25228 19854 25230 19906
rect 25230 19854 25282 19906
rect 25282 19854 25284 19906
rect 25228 19852 25284 19854
rect 25116 19516 25172 19572
rect 29036 33292 29092 33348
rect 29036 33068 29092 33124
rect 29820 32956 29876 33012
rect 29708 32620 29764 32676
rect 30044 31724 30100 31780
rect 28252 29484 28308 29540
rect 28476 30604 28532 30660
rect 29820 31276 29876 31332
rect 29708 31106 29764 31108
rect 29708 31054 29710 31106
rect 29710 31054 29762 31106
rect 29762 31054 29764 31106
rect 29708 31052 29764 31054
rect 29260 30210 29316 30212
rect 29260 30158 29262 30210
rect 29262 30158 29314 30210
rect 29314 30158 29316 30210
rect 29260 30156 29316 30158
rect 30044 31218 30100 31220
rect 30044 31166 30046 31218
rect 30046 31166 30098 31218
rect 30098 31166 30100 31218
rect 30044 31164 30100 31166
rect 30268 33068 30324 33124
rect 30492 32674 30548 32676
rect 30492 32622 30494 32674
rect 30494 32622 30546 32674
rect 30546 32622 30548 32674
rect 30492 32620 30548 32622
rect 31164 33234 31220 33236
rect 31164 33182 31166 33234
rect 31166 33182 31218 33234
rect 31218 33182 31220 33234
rect 31164 33180 31220 33182
rect 31052 32956 31108 33012
rect 30716 32562 30772 32564
rect 30716 32510 30718 32562
rect 30718 32510 30770 32562
rect 30770 32510 30772 32562
rect 30716 32508 30772 32510
rect 31388 32562 31444 32564
rect 31388 32510 31390 32562
rect 31390 32510 31442 32562
rect 31442 32510 31444 32562
rect 31388 32508 31444 32510
rect 31836 32562 31892 32564
rect 31836 32510 31838 32562
rect 31838 32510 31890 32562
rect 31890 32510 31892 32562
rect 31836 32508 31892 32510
rect 31164 32450 31220 32452
rect 31164 32398 31166 32450
rect 31166 32398 31218 32450
rect 31218 32398 31220 32450
rect 31164 32396 31220 32398
rect 31500 31164 31556 31220
rect 30940 30882 30996 30884
rect 30940 30830 30942 30882
rect 30942 30830 30994 30882
rect 30994 30830 30996 30882
rect 30940 30828 30996 30830
rect 30156 30604 30212 30660
rect 30940 30604 30996 30660
rect 30604 29708 30660 29764
rect 29820 29260 29876 29316
rect 28140 28754 28196 28756
rect 28140 28702 28142 28754
rect 28142 28702 28194 28754
rect 28194 28702 28196 28754
rect 28140 28700 28196 28702
rect 29820 28082 29876 28084
rect 29820 28030 29822 28082
rect 29822 28030 29874 28082
rect 29874 28030 29876 28082
rect 29820 28028 29876 28030
rect 31948 31106 32004 31108
rect 31948 31054 31950 31106
rect 31950 31054 32002 31106
rect 32002 31054 32004 31106
rect 31948 31052 32004 31054
rect 31612 29596 31668 29652
rect 32396 31388 32452 31444
rect 32396 30604 32452 30660
rect 32396 30268 32452 30324
rect 32060 29596 32116 29652
rect 31724 29314 31780 29316
rect 31724 29262 31726 29314
rect 31726 29262 31778 29314
rect 31778 29262 31780 29314
rect 31724 29260 31780 29262
rect 32508 30156 32564 30212
rect 32956 32620 33012 32676
rect 32844 30716 32900 30772
rect 30268 27804 30324 27860
rect 27916 27020 27972 27076
rect 28700 27074 28756 27076
rect 28700 27022 28702 27074
rect 28702 27022 28754 27074
rect 28754 27022 28756 27074
rect 28700 27020 28756 27022
rect 31836 27858 31892 27860
rect 31836 27806 31838 27858
rect 31838 27806 31890 27858
rect 31890 27806 31892 27858
rect 31836 27804 31892 27806
rect 31836 27580 31892 27636
rect 29372 26908 29428 26964
rect 28140 25564 28196 25620
rect 28588 25394 28644 25396
rect 28588 25342 28590 25394
rect 28590 25342 28642 25394
rect 28642 25342 28644 25394
rect 28588 25340 28644 25342
rect 28028 24444 28084 24500
rect 28812 23772 28868 23828
rect 30156 25564 30212 25620
rect 29596 25394 29652 25396
rect 29596 25342 29598 25394
rect 29598 25342 29650 25394
rect 29650 25342 29652 25394
rect 29596 25340 29652 25342
rect 30044 24220 30100 24276
rect 28588 23212 28644 23268
rect 29036 23660 29092 23716
rect 31388 27020 31444 27076
rect 31836 27074 31892 27076
rect 31836 27022 31838 27074
rect 31838 27022 31890 27074
rect 31890 27022 31892 27074
rect 31836 27020 31892 27022
rect 33068 31388 33124 31444
rect 33292 32562 33348 32564
rect 33292 32510 33294 32562
rect 33294 32510 33346 32562
rect 33346 32510 33348 32562
rect 33292 32508 33348 32510
rect 33292 31836 33348 31892
rect 33180 31276 33236 31332
rect 33852 32674 33908 32676
rect 33852 32622 33854 32674
rect 33854 32622 33906 32674
rect 33906 32622 33908 32674
rect 33852 32620 33908 32622
rect 33516 30828 33572 30884
rect 33180 29596 33236 29652
rect 33068 29372 33124 29428
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35644 32620 35700 32676
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 34636 31724 34692 31780
rect 34076 31164 34132 31220
rect 33964 30268 34020 30324
rect 34300 29820 34356 29876
rect 33852 29372 33908 29428
rect 33516 28700 33572 28756
rect 32172 26236 32228 26292
rect 30380 24556 30436 24612
rect 30828 24220 30884 24276
rect 30604 23548 30660 23604
rect 32284 25506 32340 25508
rect 32284 25454 32286 25506
rect 32286 25454 32338 25506
rect 32338 25454 32340 25506
rect 32284 25452 32340 25454
rect 32956 25228 33012 25284
rect 33964 27916 34020 27972
rect 33740 26402 33796 26404
rect 33740 26350 33742 26402
rect 33742 26350 33794 26402
rect 33794 26350 33796 26402
rect 33740 26348 33796 26350
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34972 29708 35028 29764
rect 35308 30156 35364 30212
rect 35532 29820 35588 29876
rect 35756 31890 35812 31892
rect 35756 31838 35758 31890
rect 35758 31838 35810 31890
rect 35810 31838 35812 31890
rect 35756 31836 35812 31838
rect 35980 30940 36036 30996
rect 35308 29426 35364 29428
rect 35308 29374 35310 29426
rect 35310 29374 35362 29426
rect 35362 29374 35364 29426
rect 35308 29372 35364 29374
rect 35756 30380 35812 30436
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34524 27186 34580 27188
rect 34524 27134 34526 27186
rect 34526 27134 34578 27186
rect 34578 27134 34580 27186
rect 34524 27132 34580 27134
rect 35980 28418 36036 28420
rect 35980 28366 35982 28418
rect 35982 28366 36034 28418
rect 36034 28366 36036 28418
rect 35980 28364 36036 28366
rect 37212 34972 37268 35028
rect 36652 33516 36708 33572
rect 36764 33404 36820 33460
rect 36540 31052 36596 31108
rect 36540 30210 36596 30212
rect 36540 30158 36542 30210
rect 36542 30158 36594 30210
rect 36594 30158 36596 30210
rect 36540 30156 36596 30158
rect 36428 28140 36484 28196
rect 33964 26236 34020 26292
rect 34076 27020 34132 27076
rect 31052 24610 31108 24612
rect 31052 24558 31054 24610
rect 31054 24558 31106 24610
rect 31106 24558 31108 24610
rect 31052 24556 31108 24558
rect 31052 23884 31108 23940
rect 32060 23884 32116 23940
rect 31164 23826 31220 23828
rect 31164 23774 31166 23826
rect 31166 23774 31218 23826
rect 31218 23774 31220 23826
rect 31164 23772 31220 23774
rect 31052 23100 31108 23156
rect 32508 23100 32564 23156
rect 26908 21644 26964 21700
rect 27356 21868 27412 21924
rect 26796 20860 26852 20916
rect 27132 21196 27188 21252
rect 26012 19852 26068 19908
rect 25340 18396 25396 18452
rect 25340 17500 25396 17556
rect 25788 19234 25844 19236
rect 25788 19182 25790 19234
rect 25790 19182 25842 19234
rect 25842 19182 25844 19234
rect 25788 19180 25844 19182
rect 25676 18172 25732 18228
rect 24780 16658 24836 16660
rect 24780 16606 24782 16658
rect 24782 16606 24834 16658
rect 24834 16606 24836 16658
rect 24780 16604 24836 16606
rect 24892 16098 24948 16100
rect 24892 16046 24894 16098
rect 24894 16046 24946 16098
rect 24946 16046 24948 16098
rect 24892 16044 24948 16046
rect 24668 15596 24724 15652
rect 24220 14588 24276 14644
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 24892 15036 24948 15092
rect 25116 16098 25172 16100
rect 25116 16046 25118 16098
rect 25118 16046 25170 16098
rect 25170 16046 25172 16098
rect 25116 16044 25172 16046
rect 25004 13356 25060 13412
rect 25116 15820 25172 15876
rect 26012 15596 26068 15652
rect 25900 15484 25956 15540
rect 26908 18396 26964 18452
rect 26236 16604 26292 16660
rect 26236 15202 26292 15204
rect 26236 15150 26238 15202
rect 26238 15150 26290 15202
rect 26290 15150 26292 15202
rect 26236 15148 26292 15150
rect 26124 13804 26180 13860
rect 26460 15372 26516 15428
rect 27020 17554 27076 17556
rect 27020 17502 27022 17554
rect 27022 17502 27074 17554
rect 27074 17502 27076 17554
rect 27020 17500 27076 17502
rect 27804 20860 27860 20916
rect 27580 19292 27636 19348
rect 28140 20076 28196 20132
rect 32172 22988 32228 23044
rect 28588 20914 28644 20916
rect 28588 20862 28590 20914
rect 28590 20862 28642 20914
rect 28642 20862 28644 20914
rect 28588 20860 28644 20862
rect 28476 19964 28532 20020
rect 28028 19740 28084 19796
rect 28588 19180 28644 19236
rect 28252 18172 28308 18228
rect 27580 17500 27636 17556
rect 29036 21868 29092 21924
rect 29820 21756 29876 21812
rect 32172 21698 32228 21700
rect 32172 21646 32174 21698
rect 32174 21646 32226 21698
rect 32226 21646 32228 21698
rect 32172 21644 32228 21646
rect 33964 24444 34020 24500
rect 32956 24050 33012 24052
rect 32956 23998 32958 24050
rect 32958 23998 33010 24050
rect 33010 23998 33012 24050
rect 32956 23996 33012 23998
rect 33068 23266 33124 23268
rect 33068 23214 33070 23266
rect 33070 23214 33122 23266
rect 33122 23214 33124 23266
rect 33068 23212 33124 23214
rect 33292 23154 33348 23156
rect 33292 23102 33294 23154
rect 33294 23102 33346 23154
rect 33346 23102 33348 23154
rect 33292 23100 33348 23102
rect 33180 22316 33236 22372
rect 30268 20860 30324 20916
rect 29148 19404 29204 19460
rect 29260 19180 29316 19236
rect 28924 18620 28980 18676
rect 30044 19404 30100 19460
rect 29820 18732 29876 18788
rect 29708 18508 29764 18564
rect 28140 15538 28196 15540
rect 28140 15486 28142 15538
rect 28142 15486 28194 15538
rect 28194 15486 28196 15538
rect 28140 15484 28196 15486
rect 27916 15148 27972 15204
rect 27244 15036 27300 15092
rect 27468 12236 27524 12292
rect 27580 13356 27636 13412
rect 28028 13858 28084 13860
rect 28028 13806 28030 13858
rect 28030 13806 28082 13858
rect 28082 13806 28084 13858
rect 28028 13804 28084 13806
rect 28924 16882 28980 16884
rect 28924 16830 28926 16882
rect 28926 16830 28978 16882
rect 28978 16830 28980 16882
rect 28924 16828 28980 16830
rect 28924 16044 28980 16100
rect 28252 12012 28308 12068
rect 28476 12684 28532 12740
rect 24444 10444 24500 10500
rect 26572 10498 26628 10500
rect 26572 10446 26574 10498
rect 26574 10446 26626 10498
rect 26626 10446 26628 10498
rect 26572 10444 26628 10446
rect 24108 9996 24164 10052
rect 5292 9660 5348 9716
rect 9212 9714 9268 9716
rect 9212 9662 9214 9714
rect 9214 9662 9266 9714
rect 9266 9662 9268 9714
rect 9212 9660 9268 9662
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 2828 7980 2884 8036
rect 3388 8034 3444 8036
rect 3388 7982 3390 8034
rect 3390 7982 3442 8034
rect 3442 7982 3444 8034
rect 3388 7980 3444 7982
rect 18396 7980 18452 8036
rect 2044 7420 2100 7476
rect 2940 7308 2996 7364
rect 3500 7362 3556 7364
rect 3500 7310 3502 7362
rect 3502 7310 3554 7362
rect 3554 7310 3556 7362
rect 3500 7308 3556 7310
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 1932 6748 1988 6804
rect 2940 6690 2996 6692
rect 2940 6638 2942 6690
rect 2942 6638 2994 6690
rect 2994 6638 2996 6690
rect 2940 6636 2996 6638
rect 16604 6636 16660 6692
rect 2044 6076 2100 6132
rect 2156 6300 2212 6356
rect 2940 5906 2996 5908
rect 2940 5854 2942 5906
rect 2942 5854 2994 5906
rect 2994 5854 2996 5906
rect 2940 5852 2996 5854
rect 1932 5404 1988 5460
rect 8876 5628 8932 5684
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 2156 4956 2212 5012
rect 1708 4732 1764 4788
rect 2492 4732 2548 4788
rect 10556 5516 10612 5572
rect 10108 5292 10164 5348
rect 1708 4060 1764 4116
rect 2044 4172 2100 4228
rect 1708 3442 1764 3444
rect 1708 3390 1710 3442
rect 1710 3390 1762 3442
rect 1762 3390 1764 3442
rect 1708 3388 1764 3390
rect 2492 4060 2548 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 7196 3724 7252 3780
rect 2940 3442 2996 3444
rect 2940 3390 2942 3442
rect 2942 3390 2994 3442
rect 2994 3390 2996 3442
rect 2940 3388 2996 3390
rect 2380 2716 2436 2772
rect 8764 3554 8820 3556
rect 8764 3502 8766 3554
rect 8766 3502 8818 3554
rect 8818 3502 8820 3554
rect 8764 3500 8820 3502
rect 12572 5180 12628 5236
rect 11788 4956 11844 5012
rect 11004 3612 11060 3668
rect 11900 3724 11956 3780
rect 12236 3554 12292 3556
rect 12236 3502 12238 3554
rect 12238 3502 12290 3554
rect 12290 3502 12292 3554
rect 12236 3500 12292 3502
rect 14700 5180 14756 5236
rect 13692 5122 13748 5124
rect 13692 5070 13694 5122
rect 13694 5070 13746 5122
rect 13746 5070 13748 5122
rect 13692 5068 13748 5070
rect 14812 5068 14868 5124
rect 13468 3500 13524 3556
rect 15596 5122 15652 5124
rect 15596 5070 15598 5122
rect 15598 5070 15650 5122
rect 15650 5070 15652 5122
rect 15596 5068 15652 5070
rect 16380 5068 16436 5124
rect 18284 5740 18340 5796
rect 17500 5122 17556 5124
rect 17500 5070 17502 5122
rect 17502 5070 17554 5122
rect 17554 5070 17556 5122
rect 17500 5068 17556 5070
rect 18060 5122 18116 5124
rect 18060 5070 18062 5122
rect 18062 5070 18114 5122
rect 18114 5070 18116 5122
rect 18060 5068 18116 5070
rect 17724 4562 17780 4564
rect 17724 4510 17726 4562
rect 17726 4510 17778 4562
rect 17778 4510 17780 4562
rect 17724 4508 17780 4510
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 22204 7308 22260 7364
rect 18620 6300 18676 6356
rect 18508 5180 18564 5236
rect 18284 4172 18340 4228
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 23884 6076 23940 6132
rect 20748 6018 20804 6020
rect 20748 5966 20750 6018
rect 20750 5966 20802 6018
rect 20802 5966 20804 6018
rect 20748 5964 20804 5966
rect 20412 5794 20468 5796
rect 20412 5742 20414 5794
rect 20414 5742 20466 5794
rect 20466 5742 20468 5794
rect 20412 5740 20468 5742
rect 20972 5740 21028 5796
rect 21644 5852 21700 5908
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20076 4450 20132 4452
rect 20076 4398 20078 4450
rect 20078 4398 20130 4450
rect 20130 4398 20132 4450
rect 20076 4396 20132 4398
rect 20412 4396 20468 4452
rect 21196 3388 21252 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22428 5906 22484 5908
rect 22428 5854 22430 5906
rect 22430 5854 22482 5906
rect 22482 5854 22484 5906
rect 22428 5852 22484 5854
rect 22204 5516 22260 5572
rect 21756 5010 21812 5012
rect 21756 4958 21758 5010
rect 21758 4958 21810 5010
rect 21810 4958 21812 5010
rect 21756 4956 21812 4958
rect 22988 5180 23044 5236
rect 23100 5292 23156 5348
rect 22764 5122 22820 5124
rect 22764 5070 22766 5122
rect 22766 5070 22818 5122
rect 22818 5070 22820 5122
rect 22764 5068 22820 5070
rect 22652 4956 22708 5012
rect 23660 5628 23716 5684
rect 23436 5068 23492 5124
rect 23212 4508 23268 4564
rect 22092 3388 22148 3444
rect 23548 3612 23604 3668
rect 23324 3500 23380 3556
rect 25228 7980 25284 8036
rect 24444 6130 24500 6132
rect 24444 6078 24446 6130
rect 24446 6078 24498 6130
rect 24498 6078 24500 6130
rect 24444 6076 24500 6078
rect 25228 6076 25284 6132
rect 24444 5122 24500 5124
rect 24444 5070 24446 5122
rect 24446 5070 24498 5122
rect 24498 5070 24500 5122
rect 24444 5068 24500 5070
rect 24220 4338 24276 4340
rect 24220 4286 24222 4338
rect 24222 4286 24274 4338
rect 24274 4286 24276 4338
rect 24220 4284 24276 4286
rect 24444 3500 24500 3556
rect 26236 4508 26292 4564
rect 28252 5740 28308 5796
rect 27020 5628 27076 5684
rect 26460 4732 26516 4788
rect 28588 12572 28644 12628
rect 28924 15314 28980 15316
rect 28924 15262 28926 15314
rect 28926 15262 28978 15314
rect 28978 15262 28980 15314
rect 28924 15260 28980 15262
rect 29596 16828 29652 16884
rect 29708 15260 29764 15316
rect 29372 12066 29428 12068
rect 29372 12014 29374 12066
rect 29374 12014 29426 12066
rect 29426 12014 29428 12066
rect 29372 12012 29428 12014
rect 29260 11676 29316 11732
rect 29820 13580 29876 13636
rect 31276 20860 31332 20916
rect 32060 20130 32116 20132
rect 32060 20078 32062 20130
rect 32062 20078 32114 20130
rect 32114 20078 32116 20130
rect 32060 20076 32116 20078
rect 31052 19906 31108 19908
rect 31052 19854 31054 19906
rect 31054 19854 31106 19906
rect 31106 19854 31108 19906
rect 31052 19852 31108 19854
rect 31052 19292 31108 19348
rect 30604 18508 30660 18564
rect 30268 17778 30324 17780
rect 30268 17726 30270 17778
rect 30270 17726 30322 17778
rect 30322 17726 30324 17778
rect 30268 17724 30324 17726
rect 30492 16828 30548 16884
rect 30156 15484 30212 15540
rect 31948 19292 32004 19348
rect 31276 18620 31332 18676
rect 31164 14700 31220 14756
rect 30380 13132 30436 13188
rect 31724 18450 31780 18452
rect 31724 18398 31726 18450
rect 31726 18398 31778 18450
rect 31778 18398 31780 18450
rect 31724 18396 31780 18398
rect 32508 19180 32564 19236
rect 32284 19010 32340 19012
rect 32284 18958 32286 19010
rect 32286 18958 32338 19010
rect 32338 18958 32340 19010
rect 32284 18956 32340 18958
rect 32172 18844 32228 18900
rect 31388 18338 31444 18340
rect 31388 18286 31390 18338
rect 31390 18286 31442 18338
rect 31442 18286 31444 18338
rect 31388 18284 31444 18286
rect 31948 18284 32004 18340
rect 33068 20018 33124 20020
rect 33068 19966 33070 20018
rect 33070 19966 33122 20018
rect 33122 19966 33124 20018
rect 33068 19964 33124 19966
rect 33292 20018 33348 20020
rect 33292 19966 33294 20018
rect 33294 19966 33346 20018
rect 33346 19966 33348 20018
rect 33292 19964 33348 19966
rect 33292 19292 33348 19348
rect 33628 20076 33684 20132
rect 32732 19068 32788 19124
rect 32508 18172 32564 18228
rect 31724 17276 31780 17332
rect 31612 15538 31668 15540
rect 31612 15486 31614 15538
rect 31614 15486 31666 15538
rect 31666 15486 31668 15538
rect 31612 15484 31668 15486
rect 30380 12290 30436 12292
rect 30380 12238 30382 12290
rect 30382 12238 30434 12290
rect 30434 12238 30436 12290
rect 30380 12236 30436 12238
rect 29596 11452 29652 11508
rect 30492 11506 30548 11508
rect 30492 11454 30494 11506
rect 30494 11454 30546 11506
rect 30546 11454 30548 11506
rect 30492 11452 30548 11454
rect 28588 9996 28644 10052
rect 33180 16882 33236 16884
rect 33180 16830 33182 16882
rect 33182 16830 33234 16882
rect 33234 16830 33236 16882
rect 33180 16828 33236 16830
rect 32396 15090 32452 15092
rect 32396 15038 32398 15090
rect 32398 15038 32450 15090
rect 32450 15038 32452 15090
rect 32396 15036 32452 15038
rect 32172 14588 32228 14644
rect 32396 14700 32452 14756
rect 32508 13858 32564 13860
rect 32508 13806 32510 13858
rect 32510 13806 32562 13858
rect 32562 13806 32564 13858
rect 32508 13804 32564 13806
rect 32732 14924 32788 14980
rect 32844 14306 32900 14308
rect 32844 14254 32846 14306
rect 32846 14254 32898 14306
rect 32898 14254 32900 14306
rect 32844 14252 32900 14254
rect 32620 13356 32676 13412
rect 32396 11564 32452 11620
rect 32732 13132 32788 13188
rect 33740 19906 33796 19908
rect 33740 19854 33742 19906
rect 33742 19854 33794 19906
rect 33794 19854 33796 19906
rect 33740 19852 33796 19854
rect 33516 19234 33572 19236
rect 33516 19182 33518 19234
rect 33518 19182 33570 19234
rect 33570 19182 33572 19234
rect 33516 19180 33572 19182
rect 33964 21532 34020 21588
rect 35532 26962 35588 26964
rect 35532 26910 35534 26962
rect 35534 26910 35586 26962
rect 35586 26910 35588 26962
rect 35532 26908 35588 26910
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34300 25452 34356 25508
rect 36876 33180 36932 33236
rect 36428 26962 36484 26964
rect 36428 26910 36430 26962
rect 36430 26910 36482 26962
rect 36482 26910 36484 26962
rect 36428 26908 36484 26910
rect 36988 30156 37044 30212
rect 36988 28642 37044 28644
rect 36988 28590 36990 28642
rect 36990 28590 37042 28642
rect 37042 28590 37044 28642
rect 36988 28588 37044 28590
rect 36652 25228 36708 25284
rect 35868 25116 35924 25172
rect 36876 25116 36932 25172
rect 35532 24444 35588 24500
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34748 23324 34804 23380
rect 34972 24108 35028 24164
rect 34412 22316 34468 22372
rect 35420 23938 35476 23940
rect 35420 23886 35422 23938
rect 35422 23886 35474 23938
rect 35474 23886 35476 23938
rect 35420 23884 35476 23886
rect 34972 22988 35028 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34860 21868 34916 21924
rect 34972 21644 35028 21700
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34076 20076 34132 20132
rect 33964 20018 34020 20020
rect 33964 19966 33966 20018
rect 33966 19966 34018 20018
rect 34018 19966 34020 20018
rect 33964 19964 34020 19966
rect 34636 19292 34692 19348
rect 33852 18508 33908 18564
rect 33628 17500 33684 17556
rect 33516 15148 33572 15204
rect 33404 14812 33460 14868
rect 33292 14700 33348 14756
rect 33068 14588 33124 14644
rect 33404 13858 33460 13860
rect 33404 13806 33406 13858
rect 33406 13806 33458 13858
rect 33458 13806 33460 13858
rect 33404 13804 33460 13806
rect 33292 13580 33348 13636
rect 33404 11506 33460 11508
rect 33404 11454 33406 11506
rect 33406 11454 33458 11506
rect 33458 11454 33460 11506
rect 33404 11452 33460 11454
rect 32956 10668 33012 10724
rect 33404 9772 33460 9828
rect 31724 8316 31780 8372
rect 32844 8316 32900 8372
rect 30268 7868 30324 7924
rect 28812 5794 28868 5796
rect 28812 5742 28814 5794
rect 28814 5742 28866 5794
rect 28866 5742 28868 5794
rect 28812 5740 28868 5742
rect 28588 4732 28644 4788
rect 28028 4562 28084 4564
rect 28028 4510 28030 4562
rect 28030 4510 28082 4562
rect 28082 4510 28084 4562
rect 28028 4508 28084 4510
rect 26236 4226 26292 4228
rect 26236 4174 26238 4226
rect 26238 4174 26290 4226
rect 26290 4174 26292 4226
rect 26236 4172 26292 4174
rect 27132 4060 27188 4116
rect 25116 3554 25172 3556
rect 25116 3502 25118 3554
rect 25118 3502 25170 3554
rect 25170 3502 25172 3554
rect 25116 3500 25172 3502
rect 25676 3500 25732 3556
rect 26460 3554 26516 3556
rect 26460 3502 26462 3554
rect 26462 3502 26514 3554
rect 26514 3502 26516 3554
rect 26460 3500 26516 3502
rect 26236 3388 26292 3444
rect 26908 3554 26964 3556
rect 26908 3502 26910 3554
rect 26910 3502 26962 3554
rect 26962 3502 26964 3554
rect 26908 3500 26964 3502
rect 27132 3500 27188 3556
rect 27244 3388 27300 3444
rect 27692 3554 27748 3556
rect 27692 3502 27694 3554
rect 27694 3502 27746 3554
rect 27746 3502 27748 3554
rect 27692 3500 27748 3502
rect 28252 3388 28308 3444
rect 29372 4396 29428 4452
rect 31276 6972 31332 7028
rect 32620 6076 32676 6132
rect 29596 3612 29652 3668
rect 29260 3442 29316 3444
rect 29260 3390 29262 3442
rect 29262 3390 29314 3442
rect 29314 3390 29316 3442
rect 29260 3388 29316 3390
rect 31500 4898 31556 4900
rect 31500 4846 31502 4898
rect 31502 4846 31554 4898
rect 31554 4846 31556 4898
rect 31500 4844 31556 4846
rect 33740 14588 33796 14644
rect 33740 14252 33796 14308
rect 34076 17724 34132 17780
rect 33852 12012 33908 12068
rect 33964 14924 34020 14980
rect 33852 10780 33908 10836
rect 33740 10444 33796 10500
rect 33516 9100 33572 9156
rect 33628 8988 33684 9044
rect 33628 6972 33684 7028
rect 34412 18844 34468 18900
rect 34188 16716 34244 16772
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35644 18508 35700 18564
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35308 17724 35364 17780
rect 35084 17554 35140 17556
rect 35084 17502 35086 17554
rect 35086 17502 35138 17554
rect 35138 17502 35140 17554
rect 35084 17500 35140 17502
rect 36204 24050 36260 24052
rect 36204 23998 36206 24050
rect 36206 23998 36258 24050
rect 36258 23998 36260 24050
rect 36204 23996 36260 23998
rect 38108 36204 38164 36260
rect 37772 35532 37828 35588
rect 37436 31164 37492 31220
rect 37324 31052 37380 31108
rect 37324 30210 37380 30212
rect 37324 30158 37326 30210
rect 37326 30158 37378 30210
rect 37378 30158 37380 30210
rect 37324 30156 37380 30158
rect 37548 30268 37604 30324
rect 37324 28588 37380 28644
rect 37436 28812 37492 28868
rect 37996 33458 38052 33460
rect 37996 33406 37998 33458
rect 37998 33406 38050 33458
rect 38050 33406 38052 33458
rect 37996 33404 38052 33406
rect 43036 39730 43092 39732
rect 43036 39678 43038 39730
rect 43038 39678 43090 39730
rect 43090 39678 43092 39730
rect 43036 39676 43092 39678
rect 40236 38668 40292 38724
rect 39452 38108 39508 38164
rect 39116 35756 39172 35812
rect 38892 35586 38948 35588
rect 38892 35534 38894 35586
rect 38894 35534 38946 35586
rect 38946 35534 38948 35586
rect 38892 35532 38948 35534
rect 38780 34076 38836 34132
rect 38108 30940 38164 30996
rect 37884 30882 37940 30884
rect 37884 30830 37886 30882
rect 37886 30830 37938 30882
rect 37938 30830 37940 30882
rect 37884 30828 37940 30830
rect 38556 30828 38612 30884
rect 39004 33516 39060 33572
rect 39004 33234 39060 33236
rect 39004 33182 39006 33234
rect 39006 33182 39058 33234
rect 39058 33182 39060 33234
rect 39004 33180 39060 33182
rect 38780 32674 38836 32676
rect 38780 32622 38782 32674
rect 38782 32622 38834 32674
rect 38834 32622 38836 32674
rect 38780 32620 38836 32622
rect 38780 31052 38836 31108
rect 38892 30716 38948 30772
rect 39228 32508 39284 32564
rect 39116 31778 39172 31780
rect 39116 31726 39118 31778
rect 39118 31726 39170 31778
rect 39170 31726 39172 31778
rect 39116 31724 39172 31726
rect 39900 35810 39956 35812
rect 39900 35758 39902 35810
rect 39902 35758 39954 35810
rect 39954 35758 39956 35810
rect 39900 35756 39956 35758
rect 41356 38162 41412 38164
rect 41356 38110 41358 38162
rect 41358 38110 41410 38162
rect 41410 38110 41412 38162
rect 41356 38108 41412 38110
rect 41132 37884 41188 37940
rect 40796 35026 40852 35028
rect 40796 34974 40798 35026
rect 40798 34974 40850 35026
rect 40850 34974 40852 35026
rect 40796 34972 40852 34974
rect 40236 33516 40292 33572
rect 39676 31724 39732 31780
rect 40012 31500 40068 31556
rect 38668 30268 38724 30324
rect 39676 31106 39732 31108
rect 39676 31054 39678 31106
rect 39678 31054 39730 31106
rect 39730 31054 39732 31106
rect 39676 31052 39732 31054
rect 39676 30156 39732 30212
rect 37660 28700 37716 28756
rect 36988 24780 37044 24836
rect 37100 26908 37156 26964
rect 37548 26908 37604 26964
rect 37212 26348 37268 26404
rect 37324 25116 37380 25172
rect 38668 26796 38724 26852
rect 39004 25506 39060 25508
rect 39004 25454 39006 25506
rect 39006 25454 39058 25506
rect 39058 25454 39060 25506
rect 39004 25452 39060 25454
rect 37772 25116 37828 25172
rect 37884 25228 37940 25284
rect 37548 24668 37604 24724
rect 37100 24610 37156 24612
rect 37100 24558 37102 24610
rect 37102 24558 37154 24610
rect 37154 24558 37156 24610
rect 37100 24556 37156 24558
rect 36876 23996 36932 24052
rect 37100 23996 37156 24052
rect 38444 25228 38500 25284
rect 38556 24780 38612 24836
rect 38108 24444 38164 24500
rect 39788 28700 39844 28756
rect 40908 32732 40964 32788
rect 40796 32620 40852 32676
rect 40572 30604 40628 30660
rect 40796 31164 40852 31220
rect 42028 37100 42084 37156
rect 41132 32732 41188 32788
rect 42364 37938 42420 37940
rect 42364 37886 42366 37938
rect 42366 37886 42418 37938
rect 42418 37886 42420 37938
rect 42364 37884 42420 37886
rect 42476 37154 42532 37156
rect 42476 37102 42478 37154
rect 42478 37102 42530 37154
rect 42530 37102 42532 37154
rect 42476 37100 42532 37102
rect 41580 32620 41636 32676
rect 41692 35698 41748 35700
rect 41692 35646 41694 35698
rect 41694 35646 41746 35698
rect 41746 35646 41748 35698
rect 41692 35644 41748 35646
rect 41804 35474 41860 35476
rect 41804 35422 41806 35474
rect 41806 35422 41858 35474
rect 41858 35422 41860 35474
rect 41804 35420 41860 35422
rect 42028 32562 42084 32564
rect 42028 32510 42030 32562
rect 42030 32510 42082 32562
rect 42082 32510 42084 32562
rect 42028 32508 42084 32510
rect 41132 31724 41188 31780
rect 41132 30268 41188 30324
rect 40796 28642 40852 28644
rect 40796 28590 40798 28642
rect 40798 28590 40850 28642
rect 40850 28590 40852 28642
rect 40796 28588 40852 28590
rect 42028 31612 42084 31668
rect 41580 30994 41636 30996
rect 41580 30942 41582 30994
rect 41582 30942 41634 30994
rect 41634 30942 41636 30994
rect 41580 30940 41636 30942
rect 42364 34130 42420 34132
rect 42364 34078 42366 34130
rect 42366 34078 42418 34130
rect 42418 34078 42420 34130
rect 42364 34076 42420 34078
rect 42140 30604 42196 30660
rect 42364 33516 42420 33572
rect 42140 30380 42196 30436
rect 41692 30210 41748 30212
rect 41692 30158 41694 30210
rect 41694 30158 41746 30210
rect 41746 30158 41748 30210
rect 41692 30156 41748 30158
rect 41580 30044 41636 30100
rect 40908 28364 40964 28420
rect 39116 24444 39172 24500
rect 39452 24556 39508 24612
rect 39116 24220 39172 24276
rect 36876 22316 36932 22372
rect 36652 22204 36708 22260
rect 36540 20524 36596 20580
rect 37100 20802 37156 20804
rect 37100 20750 37102 20802
rect 37102 20750 37154 20802
rect 37154 20750 37156 20802
rect 37100 20748 37156 20750
rect 35868 20076 35924 20132
rect 36204 19852 36260 19908
rect 35980 19346 36036 19348
rect 35980 19294 35982 19346
rect 35982 19294 36034 19346
rect 36034 19294 36036 19346
rect 35980 19292 36036 19294
rect 36092 19010 36148 19012
rect 36092 18958 36094 19010
rect 36094 18958 36146 19010
rect 36146 18958 36148 19010
rect 36092 18956 36148 18958
rect 35756 16940 35812 16996
rect 34748 16604 34804 16660
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34860 16044 34916 16100
rect 34748 15148 34804 15204
rect 34076 13858 34132 13860
rect 34076 13806 34078 13858
rect 34078 13806 34130 13858
rect 34130 13806 34132 13858
rect 34076 13804 34132 13806
rect 34300 15036 34356 15092
rect 34636 14812 34692 14868
rect 34524 13858 34580 13860
rect 34524 13806 34526 13858
rect 34526 13806 34578 13858
rect 34578 13806 34580 13858
rect 34524 13804 34580 13806
rect 34412 13356 34468 13412
rect 34412 10498 34468 10500
rect 34412 10446 34414 10498
rect 34414 10446 34466 10498
rect 34466 10446 34468 10498
rect 34412 10444 34468 10446
rect 37548 20748 37604 20804
rect 37324 18620 37380 18676
rect 37436 20524 37492 20580
rect 36988 18450 37044 18452
rect 36988 18398 36990 18450
rect 36990 18398 37042 18450
rect 37042 18398 37044 18450
rect 36988 18396 37044 18398
rect 37324 18284 37380 18340
rect 35868 16044 35924 16100
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35644 14700 35700 14756
rect 35420 14588 35476 14644
rect 35196 14364 35252 14420
rect 34860 13580 34916 13636
rect 34860 13074 34916 13076
rect 34860 13022 34862 13074
rect 34862 13022 34914 13074
rect 34914 13022 34916 13074
rect 34860 13020 34916 13022
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35084 12066 35140 12068
rect 35084 12014 35086 12066
rect 35086 12014 35138 12066
rect 35138 12014 35140 12066
rect 35084 12012 35140 12014
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35756 14364 35812 14420
rect 35980 13468 36036 13524
rect 35868 13074 35924 13076
rect 35868 13022 35870 13074
rect 35870 13022 35922 13074
rect 35922 13022 35924 13074
rect 35868 13020 35924 13022
rect 35980 12796 36036 12852
rect 36204 16940 36260 16996
rect 36316 16716 36372 16772
rect 36316 14252 36372 14308
rect 36652 16994 36708 16996
rect 36652 16942 36654 16994
rect 36654 16942 36706 16994
rect 36706 16942 36708 16994
rect 36652 16940 36708 16942
rect 36540 16044 36596 16100
rect 36764 16828 36820 16884
rect 35420 10722 35476 10724
rect 35420 10670 35422 10722
rect 35422 10670 35474 10722
rect 35474 10670 35476 10722
rect 35420 10668 35476 10670
rect 36876 11676 36932 11732
rect 37100 13804 37156 13860
rect 36540 10668 36596 10724
rect 37100 11116 37156 11172
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35644 9154 35700 9156
rect 35644 9102 35646 9154
rect 35646 9102 35698 9154
rect 35698 9102 35700 9154
rect 35644 9100 35700 9102
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 33852 6130 33908 6132
rect 33852 6078 33854 6130
rect 33854 6078 33906 6130
rect 33906 6078 33908 6130
rect 33852 6076 33908 6078
rect 34188 6748 34244 6804
rect 31164 4450 31220 4452
rect 31164 4398 31166 4450
rect 31166 4398 31218 4450
rect 31218 4398 31220 4450
rect 31164 4396 31220 4398
rect 30492 3666 30548 3668
rect 30492 3614 30494 3666
rect 30494 3614 30546 3666
rect 30546 3614 30548 3666
rect 30492 3612 30548 3614
rect 33068 4396 33124 4452
rect 33180 4338 33236 4340
rect 33180 4286 33182 4338
rect 33182 4286 33234 4338
rect 33234 4286 33236 4338
rect 33180 4284 33236 4286
rect 33404 4956 33460 5012
rect 33292 4060 33348 4116
rect 33852 4508 33908 4564
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34076 4732 34132 4788
rect 34748 4284 34804 4340
rect 33516 3724 33572 3780
rect 34076 4060 34132 4116
rect 33628 3500 33684 3556
rect 32956 3388 33012 3444
rect 33852 3442 33908 3444
rect 33852 3390 33854 3442
rect 33854 3390 33906 3442
rect 33906 3390 33908 3442
rect 33852 3388 33908 3390
rect 34300 3388 34356 3444
rect 34860 4172 34916 4228
rect 35420 4562 35476 4564
rect 35420 4510 35422 4562
rect 35422 4510 35474 4562
rect 35474 4510 35476 4562
rect 35420 4508 35476 4510
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34972 3554 35028 3556
rect 34972 3502 34974 3554
rect 34974 3502 35026 3554
rect 35026 3502 35028 3554
rect 34972 3500 35028 3502
rect 34972 3276 35028 3332
rect 37324 16044 37380 16100
rect 37660 18508 37716 18564
rect 37660 15148 37716 15204
rect 37884 21532 37940 21588
rect 37996 22204 38052 22260
rect 39228 23100 39284 23156
rect 38556 21980 38612 22036
rect 37996 19964 38052 20020
rect 38108 21868 38164 21924
rect 37548 14252 37604 14308
rect 37436 13468 37492 13524
rect 39004 21532 39060 21588
rect 38892 20130 38948 20132
rect 38892 20078 38894 20130
rect 38894 20078 38946 20130
rect 38946 20078 38948 20130
rect 38892 20076 38948 20078
rect 38332 19628 38388 19684
rect 38332 16604 38388 16660
rect 38556 18284 38612 18340
rect 38892 18508 38948 18564
rect 38444 15036 38500 15092
rect 38780 15484 38836 15540
rect 39228 19852 39284 19908
rect 39676 24668 39732 24724
rect 39452 18450 39508 18452
rect 39452 18398 39454 18450
rect 39454 18398 39506 18450
rect 39506 18398 39508 18450
rect 39452 18396 39508 18398
rect 39564 23884 39620 23940
rect 39452 16716 39508 16772
rect 39228 15372 39284 15428
rect 39116 12850 39172 12852
rect 39116 12798 39118 12850
rect 39118 12798 39170 12850
rect 39170 12798 39172 12850
rect 39116 12796 39172 12798
rect 37996 11506 38052 11508
rect 37996 11454 37998 11506
rect 37998 11454 38050 11506
rect 38050 11454 38052 11506
rect 37996 11452 38052 11454
rect 40572 26796 40628 26852
rect 40236 25452 40292 25508
rect 41020 24834 41076 24836
rect 41020 24782 41022 24834
rect 41022 24782 41074 24834
rect 41074 24782 41076 24834
rect 41020 24780 41076 24782
rect 41468 25340 41524 25396
rect 39900 24108 39956 24164
rect 40012 23660 40068 23716
rect 40012 23154 40068 23156
rect 40012 23102 40014 23154
rect 40014 23102 40066 23154
rect 40066 23102 40068 23154
rect 40012 23100 40068 23102
rect 40012 22428 40068 22484
rect 39788 19628 39844 19684
rect 40908 23266 40964 23268
rect 40908 23214 40910 23266
rect 40910 23214 40962 23266
rect 40962 23214 40964 23266
rect 40908 23212 40964 23214
rect 41132 23212 41188 23268
rect 40796 22370 40852 22372
rect 40796 22318 40798 22370
rect 40798 22318 40850 22370
rect 40850 22318 40852 22370
rect 40796 22316 40852 22318
rect 40684 20802 40740 20804
rect 40684 20750 40686 20802
rect 40686 20750 40738 20802
rect 40738 20750 40740 20802
rect 40684 20748 40740 20750
rect 40460 20076 40516 20132
rect 39900 19292 39956 19348
rect 40124 18620 40180 18676
rect 39676 15484 39732 15540
rect 39340 11676 39396 11732
rect 38668 10722 38724 10724
rect 38668 10670 38670 10722
rect 38670 10670 38722 10722
rect 38722 10670 38724 10722
rect 38668 10668 38724 10670
rect 37100 9772 37156 9828
rect 39788 15036 39844 15092
rect 40012 13468 40068 13524
rect 40348 18450 40404 18452
rect 40348 18398 40350 18450
rect 40350 18398 40402 18450
rect 40402 18398 40404 18450
rect 40348 18396 40404 18398
rect 40124 12012 40180 12068
rect 40236 15148 40292 15204
rect 39676 11228 39732 11284
rect 38556 9548 38612 9604
rect 37100 7420 37156 7476
rect 40572 16828 40628 16884
rect 40348 12236 40404 12292
rect 41020 21980 41076 22036
rect 41356 21868 41412 21924
rect 41580 23938 41636 23940
rect 41580 23886 41582 23938
rect 41582 23886 41634 23938
rect 41634 23886 41636 23938
rect 41580 23884 41636 23886
rect 42028 26796 42084 26852
rect 42476 31836 42532 31892
rect 43260 33740 43316 33796
rect 42812 31666 42868 31668
rect 42812 31614 42814 31666
rect 42814 31614 42866 31666
rect 42866 31614 42868 31666
rect 42812 31612 42868 31614
rect 43036 31500 43092 31556
rect 44044 32508 44100 32564
rect 44380 36988 44436 37044
rect 43708 31388 43764 31444
rect 44044 30940 44100 30996
rect 44380 31500 44436 31556
rect 43596 30604 43652 30660
rect 43820 30828 43876 30884
rect 44268 30828 44324 30884
rect 44044 30156 44100 30212
rect 44716 38722 44772 38724
rect 44716 38670 44718 38722
rect 44718 38670 44770 38722
rect 44770 38670 44772 38722
rect 44716 38668 44772 38670
rect 45164 41074 45220 41076
rect 45164 41022 45166 41074
rect 45166 41022 45218 41074
rect 45218 41022 45220 41074
rect 45164 41020 45220 41022
rect 45836 41074 45892 41076
rect 45836 41022 45838 41074
rect 45838 41022 45890 41074
rect 45890 41022 45892 41074
rect 45836 41020 45892 41022
rect 46172 41074 46228 41076
rect 46172 41022 46174 41074
rect 46174 41022 46226 41074
rect 46226 41022 46228 41074
rect 46172 41020 46228 41022
rect 46508 41692 46564 41748
rect 45724 38946 45780 38948
rect 45724 38894 45726 38946
rect 45726 38894 45778 38946
rect 45778 38894 45780 38946
rect 45724 38892 45780 38894
rect 45388 36988 45444 37044
rect 45500 36204 45556 36260
rect 45388 35698 45444 35700
rect 45388 35646 45390 35698
rect 45390 35646 45442 35698
rect 45442 35646 45444 35698
rect 45388 35644 45444 35646
rect 45164 33740 45220 33796
rect 45164 32508 45220 32564
rect 44940 31554 44996 31556
rect 44940 31502 44942 31554
rect 44942 31502 44994 31554
rect 44994 31502 44996 31554
rect 44940 31500 44996 31502
rect 44380 30268 44436 30324
rect 43148 28812 43204 28868
rect 44828 30098 44884 30100
rect 44828 30046 44830 30098
rect 44830 30046 44882 30098
rect 44882 30046 44884 30098
rect 44828 30044 44884 30046
rect 45052 30994 45108 30996
rect 45052 30942 45054 30994
rect 45054 30942 45106 30994
rect 45106 30942 45108 30994
rect 45052 30940 45108 30942
rect 43932 28700 43988 28756
rect 45052 29314 45108 29316
rect 45052 29262 45054 29314
rect 45054 29262 45106 29314
rect 45106 29262 45108 29314
rect 45052 29260 45108 29262
rect 44268 28140 44324 28196
rect 42364 26796 42420 26852
rect 43820 26850 43876 26852
rect 43820 26798 43822 26850
rect 43822 26798 43874 26850
rect 43874 26798 43876 26850
rect 43820 26796 43876 26798
rect 43596 26348 43652 26404
rect 41692 23548 41748 23604
rect 41468 21756 41524 21812
rect 41468 21586 41524 21588
rect 41468 21534 41470 21586
rect 41470 21534 41522 21586
rect 41522 21534 41524 21586
rect 41468 21532 41524 21534
rect 41244 20802 41300 20804
rect 41244 20750 41246 20802
rect 41246 20750 41298 20802
rect 41298 20750 41300 20802
rect 41244 20748 41300 20750
rect 42252 25228 42308 25284
rect 42476 24220 42532 24276
rect 42364 23660 42420 23716
rect 41916 23212 41972 23268
rect 42252 23548 42308 23604
rect 42028 22316 42084 22372
rect 41916 19906 41972 19908
rect 41916 19854 41918 19906
rect 41918 19854 41970 19906
rect 41970 19854 41972 19906
rect 41916 19852 41972 19854
rect 41132 18956 41188 19012
rect 40908 18172 40964 18228
rect 40796 17442 40852 17444
rect 40796 17390 40798 17442
rect 40798 17390 40850 17442
rect 40850 17390 40852 17442
rect 40796 17388 40852 17390
rect 41580 18562 41636 18564
rect 41580 18510 41582 18562
rect 41582 18510 41634 18562
rect 41634 18510 41636 18562
rect 41580 18508 41636 18510
rect 41356 18284 41412 18340
rect 41132 16940 41188 16996
rect 41020 16882 41076 16884
rect 41020 16830 41022 16882
rect 41022 16830 41074 16882
rect 41074 16830 41076 16882
rect 41020 16828 41076 16830
rect 41356 16828 41412 16884
rect 41132 15314 41188 15316
rect 41132 15262 41134 15314
rect 41134 15262 41186 15314
rect 41186 15262 41188 15314
rect 41132 15260 41188 15262
rect 40908 15036 40964 15092
rect 41244 15148 41300 15204
rect 41132 13468 41188 13524
rect 41356 11676 41412 11732
rect 41356 11452 41412 11508
rect 42140 19122 42196 19124
rect 42140 19070 42142 19122
rect 42142 19070 42194 19122
rect 42194 19070 42196 19122
rect 42140 19068 42196 19070
rect 41916 14924 41972 14980
rect 42028 18172 42084 18228
rect 42476 18284 42532 18340
rect 42588 21532 42644 21588
rect 42140 17388 42196 17444
rect 41916 12066 41972 12068
rect 41916 12014 41918 12066
rect 41918 12014 41970 12066
rect 41970 12014 41972 12066
rect 41916 12012 41972 12014
rect 42028 11676 42084 11732
rect 42252 11506 42308 11508
rect 42252 11454 42254 11506
rect 42254 11454 42306 11506
rect 42306 11454 42308 11506
rect 42252 11452 42308 11454
rect 42476 13858 42532 13860
rect 42476 13806 42478 13858
rect 42478 13806 42530 13858
rect 42530 13806 42532 13858
rect 42476 13804 42532 13806
rect 43372 26012 43428 26068
rect 42924 25394 42980 25396
rect 42924 25342 42926 25394
rect 42926 25342 42978 25394
rect 42978 25342 42980 25394
rect 42924 25340 42980 25342
rect 43148 25340 43204 25396
rect 43148 24220 43204 24276
rect 42812 24050 42868 24052
rect 42812 23998 42814 24050
rect 42814 23998 42866 24050
rect 42866 23998 42868 24050
rect 42812 23996 42868 23998
rect 45836 31836 45892 31892
rect 45612 30882 45668 30884
rect 45612 30830 45614 30882
rect 45614 30830 45666 30882
rect 45666 30830 45668 30882
rect 45612 30828 45668 30830
rect 45724 30604 45780 30660
rect 46172 30828 46228 30884
rect 45500 29314 45556 29316
rect 45500 29262 45502 29314
rect 45502 29262 45554 29314
rect 45554 29262 45556 29314
rect 45500 29260 45556 29262
rect 45164 27020 45220 27076
rect 44604 26460 44660 26516
rect 44828 26796 44884 26852
rect 44492 26066 44548 26068
rect 44492 26014 44494 26066
rect 44494 26014 44546 26066
rect 44546 26014 44548 26066
rect 44492 26012 44548 26014
rect 43596 25394 43652 25396
rect 43596 25342 43598 25394
rect 43598 25342 43650 25394
rect 43650 25342 43652 25394
rect 43596 25340 43652 25342
rect 45388 26402 45444 26404
rect 45388 26350 45390 26402
rect 45390 26350 45442 26402
rect 45442 26350 45444 26402
rect 45388 26348 45444 26350
rect 45164 26124 45220 26180
rect 44492 24220 44548 24276
rect 43820 23826 43876 23828
rect 43820 23774 43822 23826
rect 43822 23774 43874 23826
rect 43874 23774 43876 23826
rect 43820 23772 43876 23774
rect 43820 22146 43876 22148
rect 43820 22094 43822 22146
rect 43822 22094 43874 22146
rect 43874 22094 43876 22146
rect 43820 22092 43876 22094
rect 42924 20130 42980 20132
rect 42924 20078 42926 20130
rect 42926 20078 42978 20130
rect 42978 20078 42980 20130
rect 42924 20076 42980 20078
rect 42924 19628 42980 19684
rect 43372 20188 43428 20244
rect 43260 12796 43316 12852
rect 43036 12572 43092 12628
rect 42924 12290 42980 12292
rect 42924 12238 42926 12290
rect 42926 12238 42978 12290
rect 42978 12238 42980 12290
rect 42924 12236 42980 12238
rect 42140 10332 42196 10388
rect 42140 9996 42196 10052
rect 43820 21308 43876 21364
rect 43708 20524 43764 20580
rect 43820 19346 43876 19348
rect 43820 19294 43822 19346
rect 43822 19294 43874 19346
rect 43874 19294 43876 19346
rect 43820 19292 43876 19294
rect 43820 17052 43876 17108
rect 43708 16994 43764 16996
rect 43708 16942 43710 16994
rect 43710 16942 43762 16994
rect 43762 16942 43764 16994
rect 43708 16940 43764 16942
rect 44044 21644 44100 21700
rect 45836 27970 45892 27972
rect 45836 27918 45838 27970
rect 45838 27918 45890 27970
rect 45890 27918 45892 27970
rect 45836 27916 45892 27918
rect 45948 27020 46004 27076
rect 45612 26460 45668 26516
rect 45836 26236 45892 26292
rect 45724 26178 45780 26180
rect 45724 26126 45726 26178
rect 45726 26126 45778 26178
rect 45778 26126 45780 26178
rect 45724 26124 45780 26126
rect 45052 24220 45108 24276
rect 44940 24108 44996 24164
rect 44828 22428 44884 22484
rect 44828 22146 44884 22148
rect 44828 22094 44830 22146
rect 44830 22094 44882 22146
rect 44882 22094 44884 22146
rect 44828 22092 44884 22094
rect 44380 20412 44436 20468
rect 44716 21362 44772 21364
rect 44716 21310 44718 21362
rect 44718 21310 44770 21362
rect 44770 21310 44772 21362
rect 44716 21308 44772 21310
rect 44828 20578 44884 20580
rect 44828 20526 44830 20578
rect 44830 20526 44882 20578
rect 44882 20526 44884 20578
rect 44828 20524 44884 20526
rect 44492 20188 44548 20244
rect 44828 20300 44884 20356
rect 44044 18620 44100 18676
rect 44492 18620 44548 18676
rect 44268 17554 44324 17556
rect 44268 17502 44270 17554
rect 44270 17502 44322 17554
rect 44322 17502 44324 17554
rect 44268 17500 44324 17502
rect 44716 18284 44772 18340
rect 44380 16828 44436 16884
rect 44492 16940 44548 16996
rect 43484 13804 43540 13860
rect 42476 10332 42532 10388
rect 42476 10108 42532 10164
rect 38556 6748 38612 6804
rect 38556 6412 38612 6468
rect 37100 4956 37156 5012
rect 36428 4508 36484 4564
rect 37212 4844 37268 4900
rect 35868 4450 35924 4452
rect 35868 4398 35870 4450
rect 35870 4398 35922 4450
rect 35922 4398 35924 4450
rect 35868 4396 35924 4398
rect 35980 3330 36036 3332
rect 35980 3278 35982 3330
rect 35982 3278 36034 3330
rect 36034 3278 36036 3330
rect 35980 3276 36036 3278
rect 36652 4226 36708 4228
rect 36652 4174 36654 4226
rect 36654 4174 36706 4226
rect 36706 4174 36708 4226
rect 36652 4172 36708 4174
rect 36540 3724 36596 3780
rect 36316 3612 36372 3668
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 37884 3948 37940 4004
rect 39340 4898 39396 4900
rect 39340 4846 39342 4898
rect 39342 4846 39394 4898
rect 39394 4846 39396 4898
rect 39340 4844 39396 4846
rect 40348 5068 40404 5124
rect 40124 4508 40180 4564
rect 40908 4562 40964 4564
rect 40908 4510 40910 4562
rect 40910 4510 40962 4562
rect 40962 4510 40964 4562
rect 40908 4508 40964 4510
rect 38556 3388 38612 3444
rect 41356 4844 41412 4900
rect 39004 3612 39060 3668
rect 39116 3442 39172 3444
rect 39116 3390 39118 3442
rect 39118 3390 39170 3442
rect 39170 3390 39172 3442
rect 39116 3388 39172 3390
rect 39788 3948 39844 4004
rect 40236 3666 40292 3668
rect 40236 3614 40238 3666
rect 40238 3614 40290 3666
rect 40290 3614 40292 3666
rect 40236 3612 40292 3614
rect 41916 4060 41972 4116
rect 43260 8988 43316 9044
rect 43596 13468 43652 13524
rect 43596 12124 43652 12180
rect 43596 9996 43652 10052
rect 43596 9436 43652 9492
rect 43820 13634 43876 13636
rect 43820 13582 43822 13634
rect 43822 13582 43874 13634
rect 43874 13582 43876 13634
rect 43820 13580 43876 13582
rect 44380 13804 44436 13860
rect 44268 12738 44324 12740
rect 44268 12686 44270 12738
rect 44270 12686 44322 12738
rect 44322 12686 44324 12738
rect 44268 12684 44324 12686
rect 45724 24220 45780 24276
rect 45724 23660 45780 23716
rect 45052 21586 45108 21588
rect 45052 21534 45054 21586
rect 45054 21534 45106 21586
rect 45106 21534 45108 21586
rect 45052 21532 45108 21534
rect 45052 19628 45108 19684
rect 44940 18620 44996 18676
rect 44940 17500 44996 17556
rect 44940 17052 44996 17108
rect 44828 13580 44884 13636
rect 45052 12962 45108 12964
rect 45052 12910 45054 12962
rect 45054 12910 45106 12962
rect 45106 12910 45108 12962
rect 45052 12908 45108 12910
rect 43932 11228 43988 11284
rect 44044 10780 44100 10836
rect 43820 10108 43876 10164
rect 43932 9436 43988 9492
rect 42252 4732 42308 4788
rect 42364 5740 42420 5796
rect 43932 8034 43988 8036
rect 43932 7982 43934 8034
rect 43934 7982 43986 8034
rect 43986 7982 43988 8034
rect 43932 7980 43988 7982
rect 43820 5628 43876 5684
rect 44044 6524 44100 6580
rect 43596 4898 43652 4900
rect 43596 4846 43598 4898
rect 43598 4846 43650 4898
rect 43650 4846 43652 4898
rect 43596 4844 43652 4846
rect 42364 4172 42420 4228
rect 43596 4060 43652 4116
rect 42700 3666 42756 3668
rect 42700 3614 42702 3666
rect 42702 3614 42754 3666
rect 42754 3614 42756 3666
rect 42700 3612 42756 3614
rect 44268 8764 44324 8820
rect 44940 11170 44996 11172
rect 44940 11118 44942 11170
rect 44942 11118 44994 11170
rect 44994 11118 44996 11170
rect 44940 11116 44996 11118
rect 44828 10834 44884 10836
rect 44828 10782 44830 10834
rect 44830 10782 44882 10834
rect 44882 10782 44884 10834
rect 44828 10780 44884 10782
rect 44940 9602 44996 9604
rect 44940 9550 44942 9602
rect 44942 9550 44994 9602
rect 44994 9550 44996 9602
rect 44940 9548 44996 9550
rect 44716 8930 44772 8932
rect 44716 8878 44718 8930
rect 44718 8878 44770 8930
rect 44770 8878 44772 8930
rect 44716 8876 44772 8878
rect 44380 6748 44436 6804
rect 44940 8034 44996 8036
rect 44940 7982 44942 8034
rect 44942 7982 44994 8034
rect 44994 7982 44996 8034
rect 44940 7980 44996 7982
rect 44940 7474 44996 7476
rect 44940 7422 44942 7474
rect 44942 7422 44994 7474
rect 44994 7422 44996 7474
rect 44940 7420 44996 7422
rect 44940 6466 44996 6468
rect 44940 6414 44942 6466
rect 44942 6414 44994 6466
rect 44994 6414 44996 6466
rect 44940 6412 44996 6414
rect 45612 21586 45668 21588
rect 45612 21534 45614 21586
rect 45614 21534 45666 21586
rect 45666 21534 45668 21586
rect 45612 21532 45668 21534
rect 45724 20300 45780 20356
rect 45724 20130 45780 20132
rect 45724 20078 45726 20130
rect 45726 20078 45778 20130
rect 45778 20078 45780 20130
rect 45724 20076 45780 20078
rect 45500 16716 45556 16772
rect 45724 18508 45780 18564
rect 45500 16210 45556 16212
rect 45500 16158 45502 16210
rect 45502 16158 45554 16210
rect 45554 16158 45556 16210
rect 45500 16156 45556 16158
rect 45500 15484 45556 15540
rect 45388 15426 45444 15428
rect 45388 15374 45390 15426
rect 45390 15374 45442 15426
rect 45442 15374 45444 15426
rect 45388 15372 45444 15374
rect 45388 14924 45444 14980
rect 45612 15314 45668 15316
rect 45612 15262 45614 15314
rect 45614 15262 45666 15314
rect 45666 15262 45668 15314
rect 45612 15260 45668 15262
rect 45724 14812 45780 14868
rect 45612 11452 45668 11508
rect 45500 10108 45556 10164
rect 45388 9996 45444 10052
rect 45724 10722 45780 10724
rect 45724 10670 45726 10722
rect 45726 10670 45778 10722
rect 45778 10670 45780 10722
rect 45724 10668 45780 10670
rect 45276 6748 45332 6804
rect 45724 7420 45780 7476
rect 45612 6636 45668 6692
rect 45500 5404 45556 5460
rect 44940 5122 44996 5124
rect 44940 5070 44942 5122
rect 44942 5070 44994 5122
rect 44994 5070 44996 5122
rect 44940 5068 44996 5070
rect 44156 4396 44212 4452
rect 46060 26908 46116 26964
rect 46060 26124 46116 26180
rect 46060 23714 46116 23716
rect 46060 23662 46062 23714
rect 46062 23662 46114 23714
rect 46114 23662 46116 23714
rect 46060 23660 46116 23662
rect 46172 19516 46228 19572
rect 46284 20412 46340 20468
rect 46060 19122 46116 19124
rect 46060 19070 46062 19122
rect 46062 19070 46114 19122
rect 46114 19070 46116 19122
rect 46060 19068 46116 19070
rect 46060 18172 46116 18228
rect 46060 17554 46116 17556
rect 46060 17502 46062 17554
rect 46062 17502 46114 17554
rect 46114 17502 46116 17554
rect 46060 17500 46116 17502
rect 46060 16882 46116 16884
rect 46060 16830 46062 16882
rect 46062 16830 46114 16882
rect 46114 16830 46116 16882
rect 46060 16828 46116 16830
rect 45948 14588 46004 14644
rect 45948 14418 46004 14420
rect 45948 14366 45950 14418
rect 45950 14366 46002 14418
rect 46002 14366 46004 14418
rect 45948 14364 46004 14366
rect 46172 12962 46228 12964
rect 46172 12910 46174 12962
rect 46174 12910 46226 12962
rect 46226 12910 46228 12962
rect 46172 12908 46228 12910
rect 46060 10108 46116 10164
rect 46508 16940 46564 16996
rect 46620 14588 46676 14644
rect 45836 6524 45892 6580
rect 46060 8092 46116 8148
rect 46172 6076 46228 6132
rect 45836 4450 45892 4452
rect 45836 4398 45838 4450
rect 45838 4398 45890 4450
rect 45890 4398 45892 4450
rect 45836 4396 45892 4398
rect 45612 4172 45668 4228
rect 43036 3388 43092 3444
rect 46172 5404 46228 5460
rect 46060 3612 46116 3668
rect 44380 2044 44436 2100
rect 43596 1372 43652 1428
rect 45276 2716 45332 2772
rect 44828 700 44884 756
rect 45276 28 45332 84
<< metal3 >>
rect 27570 45276 27580 45332
rect 27636 45276 28812 45332
rect 28868 45276 28878 45332
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 8082 44492 8092 44548
rect 8148 44492 9772 44548
rect 9828 44492 9838 44548
rect 24882 44492 24892 44548
rect 24948 44492 25564 44548
rect 25620 44492 25630 44548
rect 29586 44492 29596 44548
rect 29652 44492 30380 44548
rect 30436 44492 30446 44548
rect 30930 44492 30940 44548
rect 30996 44492 32620 44548
rect 32676 44492 32686 44548
rect 36306 44492 36316 44548
rect 36372 44492 37100 44548
rect 37156 44492 37166 44548
rect 38994 44492 39004 44548
rect 39060 44492 40236 44548
rect 40292 44492 40302 44548
rect 42354 44492 42364 44548
rect 42420 44492 44044 44548
rect 44100 44492 44110 44548
rect 47200 44436 48000 44464
rect 25330 44380 25340 44436
rect 25396 44380 26908 44436
rect 26964 44380 26974 44436
rect 36754 44380 36764 44436
rect 36820 44380 38780 44436
rect 38836 44380 38846 44436
rect 45714 44380 45724 44436
rect 45780 44380 48000 44436
rect 47200 44352 48000 44380
rect 38882 44268 38892 44324
rect 38948 44268 43708 44324
rect 43764 44268 43774 44324
rect 14802 44156 14812 44212
rect 14868 44156 15932 44212
rect 15988 44156 15998 44212
rect 7746 44044 7756 44100
rect 7812 44044 9324 44100
rect 9380 44044 9390 44100
rect 44034 44044 44044 44100
rect 44100 44044 45836 44100
rect 45892 44044 45902 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 47200 43764 48000 43792
rect 45602 43708 45612 43764
rect 45668 43708 46172 43764
rect 46228 43708 48000 43764
rect 47200 43680 48000 43708
rect 23314 43596 23324 43652
rect 23380 43596 23996 43652
rect 24052 43596 24062 43652
rect 24210 43596 24220 43652
rect 24276 43596 25228 43652
rect 25284 43596 25294 43652
rect 31602 43596 31612 43652
rect 31668 43596 32060 43652
rect 32116 43596 32126 43652
rect 41794 43596 41804 43652
rect 41860 43596 42588 43652
rect 42644 43596 43036 43652
rect 43092 43596 43102 43652
rect 20850 43484 20860 43540
rect 20916 43484 21532 43540
rect 21588 43484 22092 43540
rect 22148 43484 22158 43540
rect 22978 43484 22988 43540
rect 23044 43484 23772 43540
rect 23828 43484 24332 43540
rect 24388 43484 24398 43540
rect 27794 43484 27804 43540
rect 27860 43484 28476 43540
rect 28532 43484 28542 43540
rect 29810 43484 29820 43540
rect 29876 43484 30156 43540
rect 30212 43484 30716 43540
rect 30772 43484 30782 43540
rect 38546 43484 38556 43540
rect 38612 43484 39004 43540
rect 39060 43484 39070 43540
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 47200 43092 48000 43120
rect 46050 43036 46060 43092
rect 46116 43036 48000 43092
rect 47200 43008 48000 43036
rect 28466 42924 28476 42980
rect 28532 42924 33740 42980
rect 33796 42924 33806 42980
rect 18722 42700 18732 42756
rect 18788 42700 20636 42756
rect 20692 42700 20702 42756
rect 21410 42700 21420 42756
rect 21476 42700 22428 42756
rect 22484 42700 22494 42756
rect 34850 42700 34860 42756
rect 34916 42700 38220 42756
rect 38276 42700 38286 42756
rect 39666 42700 39676 42756
rect 39732 42700 42812 42756
rect 42868 42700 42878 42756
rect 39890 42588 39900 42644
rect 39956 42588 41244 42644
rect 41300 42588 41310 42644
rect 1698 42476 1708 42532
rect 1764 42476 1774 42532
rect 0 42420 800 42448
rect 1708 42420 1764 42476
rect 47200 42420 48000 42448
rect 0 42364 1764 42420
rect 46050 42364 46060 42420
rect 46116 42364 48000 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 47200 42336 48000 42364
rect 27122 42140 27132 42196
rect 27188 42140 29932 42196
rect 29988 42140 29998 42196
rect 30482 42140 30492 42196
rect 30548 42140 32172 42196
rect 32228 42140 32238 42196
rect 27570 42028 27580 42084
rect 27636 42028 31836 42084
rect 31892 42028 31902 42084
rect 35522 41916 35532 41972
rect 35588 41916 37100 41972
rect 37156 41916 37166 41972
rect 47200 41748 48000 41776
rect 46498 41692 46508 41748
rect 46564 41692 48000 41748
rect 47200 41664 48000 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 47200 41076 48000 41104
rect 45154 41020 45164 41076
rect 45220 41020 45836 41076
rect 45892 41020 45902 41076
rect 46162 41020 46172 41076
rect 46228 41020 48000 41076
rect 47200 40992 48000 41020
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 38546 39676 38556 39732
rect 38612 39676 43036 39732
rect 43092 39676 43102 39732
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 36306 38892 36316 38948
rect 36372 38892 45724 38948
rect 45780 38892 45790 38948
rect 40226 38668 40236 38724
rect 40292 38668 44716 38724
rect 44772 38668 44782 38724
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 39442 38108 39452 38164
rect 39508 38108 41356 38164
rect 41412 38108 41422 38164
rect 17042 37884 17052 37940
rect 17108 37884 18844 37940
rect 18900 37884 18910 37940
rect 41122 37884 41132 37940
rect 41188 37884 42364 37940
rect 42420 37884 42430 37940
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 12786 37324 12796 37380
rect 12852 37324 13804 37380
rect 13860 37324 13870 37380
rect 42018 37100 42028 37156
rect 42084 37100 42476 37156
rect 42532 37100 42542 37156
rect 44370 36988 44380 37044
rect 44436 36988 45388 37044
rect 45444 36988 45454 37044
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 21186 36316 21196 36372
rect 21252 36316 23548 36372
rect 23604 36316 23614 36372
rect 38098 36204 38108 36260
rect 38164 36204 45500 36260
rect 45556 36204 45566 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 39106 35756 39116 35812
rect 39172 35756 39900 35812
rect 39956 35756 39966 35812
rect 41682 35644 41692 35700
rect 41748 35644 45388 35700
rect 45444 35644 45454 35700
rect 37762 35532 37772 35588
rect 37828 35532 38892 35588
rect 38948 35532 38958 35588
rect 34626 35420 34636 35476
rect 34692 35420 41804 35476
rect 41860 35420 41870 35476
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 14018 35196 14028 35252
rect 14084 35196 15148 35252
rect 15204 35196 15214 35252
rect 16370 35196 16380 35252
rect 16436 35196 17836 35252
rect 17892 35196 17902 35252
rect 9986 34972 9996 35028
rect 10052 34972 14700 35028
rect 14756 34972 14766 35028
rect 20626 34972 20636 35028
rect 20692 34972 22316 35028
rect 22372 34972 22382 35028
rect 37202 34972 37212 35028
rect 37268 34972 40796 35028
rect 40852 34972 40862 35028
rect 1698 34748 1708 34804
rect 1764 34748 7308 34804
rect 7364 34748 7374 34804
rect 24322 34748 24332 34804
rect 24388 34748 26124 34804
rect 26180 34748 26190 34804
rect 16594 34636 16604 34692
rect 16660 34636 17948 34692
rect 18004 34636 18014 34692
rect 21298 34524 21308 34580
rect 21364 34524 22428 34580
rect 22484 34524 22494 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 13234 34300 13244 34356
rect 13300 34300 15820 34356
rect 15876 34300 15886 34356
rect 6066 34188 6076 34244
rect 6132 34188 8540 34244
rect 8596 34188 8606 34244
rect 19730 34188 19740 34244
rect 19796 34188 28924 34244
rect 28980 34188 28990 34244
rect 38770 34076 38780 34132
rect 38836 34076 42364 34132
rect 42420 34076 42430 34132
rect 5842 33964 5852 34020
rect 5908 33964 6188 34020
rect 6244 33964 6254 34020
rect 6626 33964 6636 34020
rect 6692 33964 7532 34020
rect 7588 33964 7598 34020
rect 15092 33964 18396 34020
rect 18452 33964 18462 34020
rect 15092 33908 15148 33964
rect 6738 33852 6748 33908
rect 6804 33852 15148 33908
rect 15586 33740 15596 33796
rect 15652 33740 19516 33796
rect 19572 33740 19582 33796
rect 43250 33740 43260 33796
rect 43316 33740 45164 33796
rect 45220 33740 45230 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 16034 33628 16044 33684
rect 16100 33628 16828 33684
rect 16884 33628 16894 33684
rect 17266 33516 17276 33572
rect 17332 33516 19628 33572
rect 19684 33516 19694 33572
rect 36642 33516 36652 33572
rect 36708 33516 39004 33572
rect 39060 33516 39070 33572
rect 40226 33516 40236 33572
rect 40292 33516 42364 33572
rect 42420 33516 42430 33572
rect 36754 33404 36764 33460
rect 36820 33404 37996 33460
rect 38052 33404 38062 33460
rect 9986 33292 9996 33348
rect 10052 33292 11452 33348
rect 11508 33292 11518 33348
rect 13458 33292 13468 33348
rect 13524 33292 17500 33348
rect 17556 33292 17566 33348
rect 25778 33292 25788 33348
rect 25844 33292 29036 33348
rect 29092 33292 29102 33348
rect 23202 33180 23212 33236
rect 23268 33180 25676 33236
rect 25732 33180 25742 33236
rect 28690 33180 28700 33236
rect 28756 33180 31164 33236
rect 31220 33180 31230 33236
rect 36866 33180 36876 33236
rect 36932 33180 39004 33236
rect 39060 33180 39070 33236
rect 21634 33068 21644 33124
rect 21700 33068 23324 33124
rect 23380 33068 23390 33124
rect 24882 33068 24892 33124
rect 24948 33068 27244 33124
rect 27300 33068 27310 33124
rect 29026 33068 29036 33124
rect 29092 33068 30268 33124
rect 30324 33068 30334 33124
rect 21746 32956 21756 33012
rect 21812 32956 25116 33012
rect 25172 32956 25182 33012
rect 29810 32956 29820 33012
rect 29876 32956 31052 33012
rect 31108 32956 31118 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 40898 32732 40908 32788
rect 40964 32732 41132 32788
rect 41188 32732 41198 32788
rect 6962 32620 6972 32676
rect 7028 32620 9436 32676
rect 9492 32620 9502 32676
rect 29698 32620 29708 32676
rect 29764 32620 30492 32676
rect 30548 32620 30558 32676
rect 32946 32620 32956 32676
rect 33012 32620 33852 32676
rect 33908 32620 33918 32676
rect 35634 32620 35644 32676
rect 35700 32620 38780 32676
rect 38836 32620 38846 32676
rect 40786 32620 40796 32676
rect 40852 32620 41580 32676
rect 41636 32620 41646 32676
rect 2930 32508 2940 32564
rect 2996 32508 3612 32564
rect 3668 32508 3678 32564
rect 28242 32508 28252 32564
rect 28308 32508 30716 32564
rect 30772 32508 31388 32564
rect 31444 32508 31836 32564
rect 31892 32508 33292 32564
rect 33348 32508 33358 32564
rect 39218 32508 39228 32564
rect 39284 32508 42028 32564
rect 42084 32508 42094 32564
rect 44034 32508 44044 32564
rect 44100 32508 45164 32564
rect 45220 32508 45230 32564
rect 28130 32396 28140 32452
rect 28196 32396 31164 32452
rect 31220 32396 31230 32452
rect 16482 32284 16492 32340
rect 16548 32284 17388 32340
rect 17444 32284 17454 32340
rect 47200 32256 48000 32368
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 18050 32060 18060 32116
rect 18116 32060 21532 32116
rect 21588 32060 21598 32116
rect 20850 31948 20860 32004
rect 20916 31948 22764 32004
rect 22820 31948 22830 32004
rect 2706 31836 2716 31892
rect 2772 31836 3500 31892
rect 3556 31836 3566 31892
rect 17826 31836 17836 31892
rect 17892 31836 18732 31892
rect 18788 31836 18798 31892
rect 25106 31836 25116 31892
rect 25172 31836 26236 31892
rect 26292 31836 26302 31892
rect 33282 31836 33292 31892
rect 33348 31836 35756 31892
rect 35812 31836 35822 31892
rect 42466 31836 42476 31892
rect 42532 31836 45836 31892
rect 45892 31836 45902 31892
rect 9202 31724 9212 31780
rect 9268 31724 9548 31780
rect 9604 31724 9614 31780
rect 15810 31724 15820 31780
rect 15876 31724 17612 31780
rect 17668 31724 17678 31780
rect 24770 31724 24780 31780
rect 24836 31724 25228 31780
rect 25284 31724 26012 31780
rect 26068 31724 26572 31780
rect 26628 31724 26638 31780
rect 30034 31724 30044 31780
rect 30100 31724 34636 31780
rect 34692 31724 34702 31780
rect 39106 31724 39116 31780
rect 39172 31724 39676 31780
rect 39732 31724 41132 31780
rect 41188 31724 41198 31780
rect 0 31668 800 31696
rect 0 31612 15484 31668
rect 15540 31612 15550 31668
rect 42018 31612 42028 31668
rect 42084 31612 42812 31668
rect 42868 31612 42878 31668
rect 0 31584 800 31612
rect 47200 31584 48000 31696
rect 2034 31500 2044 31556
rect 2100 31500 6076 31556
rect 6132 31500 6142 31556
rect 40002 31500 40012 31556
rect 40068 31500 43036 31556
rect 43092 31500 43102 31556
rect 44370 31500 44380 31556
rect 44436 31500 44940 31556
rect 44996 31500 45006 31556
rect 43036 31444 43092 31500
rect 22194 31388 22204 31444
rect 22260 31388 23548 31444
rect 23604 31388 23614 31444
rect 32386 31388 32396 31444
rect 32452 31388 33068 31444
rect 33124 31388 33134 31444
rect 43036 31388 43708 31444
rect 43764 31388 45108 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 29810 31276 29820 31332
rect 29876 31276 33180 31332
rect 33236 31276 33246 31332
rect 26852 31164 30044 31220
rect 30100 31164 30110 31220
rect 31490 31164 31500 31220
rect 31556 31164 32900 31220
rect 34066 31164 34076 31220
rect 34132 31164 34142 31220
rect 37426 31164 37436 31220
rect 37492 31164 40796 31220
rect 40852 31164 40862 31220
rect 24210 31052 24220 31108
rect 24276 31052 25228 31108
rect 25284 31052 25294 31108
rect 26852 30996 26908 31164
rect 32844 31108 32900 31164
rect 34076 31108 34132 31164
rect 29698 31052 29708 31108
rect 29764 31052 31948 31108
rect 32004 31052 32014 31108
rect 32844 31052 34132 31108
rect 36530 31052 36540 31108
rect 36596 31052 37324 31108
rect 37380 31052 37390 31108
rect 38770 31052 38780 31108
rect 38836 31052 39676 31108
rect 39732 31052 39742 31108
rect 45052 30996 45108 31388
rect 9986 30940 9996 30996
rect 10052 30940 12124 30996
rect 12180 30940 13356 30996
rect 13412 30940 13422 30996
rect 26674 30940 26684 30996
rect 26740 30940 26908 30996
rect 35970 30940 35980 30996
rect 36036 30940 38108 30996
rect 38164 30940 38174 30996
rect 41570 30940 41580 30996
rect 41636 30940 44044 30996
rect 44100 30940 44110 30996
rect 45042 30940 45052 30996
rect 45108 30940 45118 30996
rect 47200 30912 48000 31024
rect 5618 30828 5628 30884
rect 5684 30828 6188 30884
rect 6244 30828 7196 30884
rect 7252 30828 7262 30884
rect 7970 30828 7980 30884
rect 8036 30828 10108 30884
rect 10164 30828 10174 30884
rect 10434 30828 10444 30884
rect 10500 30828 11004 30884
rect 11060 30828 11452 30884
rect 11508 30828 12236 30884
rect 12292 30828 12302 30884
rect 23762 30828 23772 30884
rect 23828 30828 25228 30884
rect 25284 30828 25294 30884
rect 27234 30828 27244 30884
rect 27300 30828 30940 30884
rect 30996 30828 31006 30884
rect 33506 30828 33516 30884
rect 33572 30828 37884 30884
rect 37940 30828 37950 30884
rect 38546 30828 38556 30884
rect 38612 30828 43820 30884
rect 43876 30828 43886 30884
rect 44258 30828 44268 30884
rect 44324 30828 45612 30884
rect 45668 30828 46172 30884
rect 46228 30828 46238 30884
rect 10882 30716 10892 30772
rect 10948 30716 11788 30772
rect 11844 30716 11854 30772
rect 18386 30716 18396 30772
rect 18452 30716 18732 30772
rect 18788 30716 18798 30772
rect 32834 30716 32844 30772
rect 32900 30716 38892 30772
rect 38948 30716 38958 30772
rect 14018 30604 14028 30660
rect 14084 30604 17388 30660
rect 17444 30604 17454 30660
rect 28466 30604 28476 30660
rect 28532 30604 30156 30660
rect 30212 30604 30222 30660
rect 30930 30604 30940 30660
rect 30996 30604 32396 30660
rect 32452 30604 32462 30660
rect 40562 30604 40572 30660
rect 40628 30604 42140 30660
rect 42196 30604 42206 30660
rect 43586 30604 43596 30660
rect 43652 30604 45724 30660
rect 45780 30604 45790 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 1586 30380 1596 30436
rect 1652 30380 2380 30436
rect 2436 30380 2446 30436
rect 35746 30380 35756 30436
rect 35812 30380 42140 30436
rect 42196 30380 42206 30436
rect 2258 30268 2268 30324
rect 2324 30268 3388 30324
rect 32386 30268 32396 30324
rect 32452 30268 33964 30324
rect 34020 30268 34030 30324
rect 37538 30268 37548 30324
rect 37604 30268 38668 30324
rect 38724 30268 38734 30324
rect 41122 30268 41132 30324
rect 41188 30268 44380 30324
rect 44436 30268 44446 30324
rect 3332 30212 3388 30268
rect 47200 30240 48000 30352
rect 3332 30156 4732 30212
rect 4788 30156 5628 30212
rect 5684 30156 5694 30212
rect 12338 30156 12348 30212
rect 12404 30156 14252 30212
rect 14308 30156 14318 30212
rect 17154 30156 17164 30212
rect 17220 30156 19068 30212
rect 19124 30156 20636 30212
rect 20692 30156 20702 30212
rect 25666 30156 25676 30212
rect 25732 30156 26012 30212
rect 26068 30156 28140 30212
rect 28196 30156 29260 30212
rect 29316 30156 32508 30212
rect 32564 30156 32574 30212
rect 35298 30156 35308 30212
rect 35364 30156 36540 30212
rect 36596 30156 36988 30212
rect 37044 30156 37324 30212
rect 37380 30156 37390 30212
rect 39666 30156 39676 30212
rect 39732 30156 41692 30212
rect 41748 30156 44044 30212
rect 44100 30156 44110 30212
rect 4050 30044 4060 30100
rect 4116 30044 6076 30100
rect 6132 30044 6142 30100
rect 12450 30044 12460 30100
rect 12516 30044 13468 30100
rect 13524 30044 13534 30100
rect 14578 30044 14588 30100
rect 14644 30044 15260 30100
rect 15316 30044 16156 30100
rect 16212 30044 16828 30100
rect 16884 30044 17612 30100
rect 17668 30044 17678 30100
rect 20738 30044 20748 30100
rect 20804 30044 21644 30100
rect 21700 30044 21710 30100
rect 24882 30044 24892 30100
rect 24948 30044 27916 30100
rect 27972 30044 27982 30100
rect 41570 30044 41580 30100
rect 41636 30044 44828 30100
rect 44884 30044 44894 30100
rect 15922 29932 15932 29988
rect 15988 29932 21980 29988
rect 22036 29932 22046 29988
rect 22754 29932 22764 29988
rect 22820 29932 26012 29988
rect 26068 29932 26078 29988
rect 7522 29820 7532 29876
rect 7588 29820 8428 29876
rect 8484 29820 8494 29876
rect 34290 29820 34300 29876
rect 34356 29820 35532 29876
rect 35588 29820 35598 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 16258 29708 16268 29764
rect 16324 29708 18172 29764
rect 18228 29708 18238 29764
rect 30594 29708 30604 29764
rect 30660 29708 34972 29764
rect 35028 29708 35038 29764
rect 3042 29596 3052 29652
rect 3108 29596 8204 29652
rect 8260 29596 8270 29652
rect 11666 29596 11676 29652
rect 11732 29596 12348 29652
rect 12404 29596 12414 29652
rect 16370 29596 16380 29652
rect 16436 29596 19068 29652
rect 19124 29596 19134 29652
rect 31602 29596 31612 29652
rect 31668 29596 32060 29652
rect 32116 29596 33180 29652
rect 33236 29596 33246 29652
rect 47200 29568 48000 29680
rect 27570 29484 27580 29540
rect 27636 29484 28252 29540
rect 28308 29484 28318 29540
rect 3490 29372 3500 29428
rect 3556 29372 5068 29428
rect 5124 29372 5134 29428
rect 7186 29372 7196 29428
rect 7252 29372 8316 29428
rect 8372 29372 9660 29428
rect 9716 29372 9726 29428
rect 16930 29372 16940 29428
rect 16996 29372 18284 29428
rect 18340 29372 18350 29428
rect 33058 29372 33068 29428
rect 33124 29372 33852 29428
rect 33908 29372 35308 29428
rect 35364 29372 35374 29428
rect 7410 29260 7420 29316
rect 7476 29260 8764 29316
rect 8820 29260 8830 29316
rect 29810 29260 29820 29316
rect 29876 29260 31724 29316
rect 31780 29260 31790 29316
rect 45042 29260 45052 29316
rect 45108 29260 45500 29316
rect 45556 29260 45566 29316
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 47200 28896 48000 29008
rect 20514 28812 20524 28868
rect 20580 28812 21644 28868
rect 21700 28812 24444 28868
rect 24500 28812 25452 28868
rect 25508 28812 25518 28868
rect 37426 28812 37436 28868
rect 37492 28812 43148 28868
rect 43204 28812 43214 28868
rect 4946 28700 4956 28756
rect 5012 28700 5628 28756
rect 5684 28700 5694 28756
rect 12226 28700 12236 28756
rect 12292 28700 13692 28756
rect 13748 28700 14028 28756
rect 14084 28700 14476 28756
rect 14532 28700 14542 28756
rect 21522 28700 21532 28756
rect 21588 28700 24220 28756
rect 24276 28700 24286 28756
rect 27122 28700 27132 28756
rect 27188 28700 28140 28756
rect 28196 28700 28206 28756
rect 33506 28700 33516 28756
rect 33572 28700 37660 28756
rect 37716 28700 37726 28756
rect 39778 28700 39788 28756
rect 39844 28700 43932 28756
rect 43988 28700 43998 28756
rect 4274 28588 4284 28644
rect 4340 28588 6300 28644
rect 6356 28588 6366 28644
rect 6626 28588 6636 28644
rect 6692 28588 6972 28644
rect 7028 28588 7420 28644
rect 7476 28588 7486 28644
rect 11218 28588 11228 28644
rect 11284 28588 12012 28644
rect 12068 28588 12078 28644
rect 13346 28588 13356 28644
rect 13412 28588 15148 28644
rect 15204 28588 17164 28644
rect 17220 28588 17230 28644
rect 20188 28588 20748 28644
rect 20804 28588 26572 28644
rect 26628 28588 27020 28644
rect 27076 28588 27086 28644
rect 36978 28588 36988 28644
rect 37044 28588 37324 28644
rect 37380 28588 40796 28644
rect 40852 28588 40862 28644
rect 6636 28532 6692 28588
rect 20188 28532 20244 28588
rect 5954 28476 5964 28532
rect 6020 28476 6692 28532
rect 12114 28476 12124 28532
rect 12180 28476 13580 28532
rect 13636 28476 14924 28532
rect 14980 28476 14990 28532
rect 18274 28476 18284 28532
rect 18340 28476 20244 28532
rect 23762 28476 23772 28532
rect 23828 28476 25004 28532
rect 25060 28476 25070 28532
rect 9874 28364 9884 28420
rect 9940 28364 10444 28420
rect 10500 28364 12236 28420
rect 12292 28364 12302 28420
rect 35970 28364 35980 28420
rect 36036 28364 40908 28420
rect 40964 28364 40974 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 47200 28224 48000 28336
rect 36418 28140 36428 28196
rect 36484 28140 44268 28196
rect 44324 28140 44334 28196
rect 2258 28028 2268 28084
rect 2324 28028 3500 28084
rect 3556 28028 3566 28084
rect 27346 28028 27356 28084
rect 27412 28028 29820 28084
rect 29876 28028 29886 28084
rect 1922 27916 1932 27972
rect 1988 27916 3276 27972
rect 3332 27916 5964 27972
rect 6020 27916 6030 27972
rect 18386 27916 18396 27972
rect 18452 27916 19068 27972
rect 19124 27916 19740 27972
rect 19796 27916 19806 27972
rect 33954 27916 33964 27972
rect 34020 27916 45836 27972
rect 45892 27916 45902 27972
rect 4050 27804 4060 27860
rect 4116 27804 6076 27860
rect 6132 27804 6142 27860
rect 8642 27804 8652 27860
rect 8708 27804 10108 27860
rect 10164 27804 12908 27860
rect 12964 27804 13468 27860
rect 13524 27804 13534 27860
rect 23650 27804 23660 27860
rect 23716 27804 27468 27860
rect 27524 27804 27534 27860
rect 30258 27804 30268 27860
rect 30324 27804 31836 27860
rect 31892 27804 31902 27860
rect 24098 27692 24108 27748
rect 24164 27692 25228 27748
rect 25284 27692 25294 27748
rect 24994 27580 25004 27636
rect 25060 27580 31836 27636
rect 31892 27580 31902 27636
rect 47200 27552 48000 27664
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 22642 27244 22652 27300
rect 22708 27244 25004 27300
rect 25060 27244 25070 27300
rect 4050 27132 4060 27188
rect 4116 27132 9772 27188
rect 9828 27132 9838 27188
rect 24434 27132 24444 27188
rect 24500 27132 25116 27188
rect 25172 27132 26908 27188
rect 27570 27132 27580 27188
rect 27636 27132 34524 27188
rect 34580 27132 34590 27188
rect 26852 27076 26908 27132
rect 13458 27020 13468 27076
rect 13524 27020 17388 27076
rect 17444 27020 17454 27076
rect 26852 27020 27916 27076
rect 27972 27020 28700 27076
rect 28756 27020 31388 27076
rect 31444 27020 31454 27076
rect 31826 27020 31836 27076
rect 31892 27020 34076 27076
rect 34132 27020 34142 27076
rect 45154 27020 45164 27076
rect 45220 27020 45948 27076
rect 46004 27020 46014 27076
rect 47200 26964 48000 26992
rect 3042 26908 3052 26964
rect 3108 26908 11676 26964
rect 11732 26908 11742 26964
rect 19730 26908 19740 26964
rect 19796 26908 21196 26964
rect 21252 26908 21262 26964
rect 24994 26908 25004 26964
rect 25060 26908 26796 26964
rect 26852 26908 26862 26964
rect 29362 26908 29372 26964
rect 29428 26908 35532 26964
rect 35588 26908 35598 26964
rect 36418 26908 36428 26964
rect 36484 26908 37100 26964
rect 37156 26908 37548 26964
rect 37604 26908 37614 26964
rect 46050 26908 46060 26964
rect 46116 26908 48000 26964
rect 47200 26880 48000 26908
rect 4722 26796 4732 26852
rect 4788 26796 6412 26852
rect 6468 26796 6478 26852
rect 17490 26796 17500 26852
rect 17556 26796 18284 26852
rect 18340 26796 18350 26852
rect 38658 26796 38668 26852
rect 38724 26796 40572 26852
rect 40628 26796 40638 26852
rect 42018 26796 42028 26852
rect 42084 26796 42364 26852
rect 42420 26796 42430 26852
rect 43810 26796 43820 26852
rect 43876 26796 44828 26852
rect 44884 26796 44894 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 3154 26460 3164 26516
rect 3220 26460 3948 26516
rect 4004 26460 4014 26516
rect 8530 26460 8540 26516
rect 8596 26460 9660 26516
rect 9716 26460 9726 26516
rect 17042 26460 17052 26516
rect 17108 26460 18844 26516
rect 18900 26460 18910 26516
rect 44594 26460 44604 26516
rect 44660 26460 45612 26516
rect 45668 26460 45678 26516
rect 3042 26348 3052 26404
rect 3108 26348 13020 26404
rect 13076 26348 13086 26404
rect 33730 26348 33740 26404
rect 33796 26348 37212 26404
rect 37268 26348 37278 26404
rect 43586 26348 43596 26404
rect 43652 26348 45388 26404
rect 45444 26348 45454 26404
rect 47200 26292 48000 26320
rect 5170 26236 5180 26292
rect 5236 26236 5628 26292
rect 5684 26236 7980 26292
rect 8036 26236 8046 26292
rect 9650 26236 9660 26292
rect 9716 26236 11788 26292
rect 11844 26236 13244 26292
rect 13300 26236 13310 26292
rect 15474 26236 15484 26292
rect 15540 26236 22204 26292
rect 22260 26236 22270 26292
rect 23090 26236 23100 26292
rect 23156 26236 25676 26292
rect 25732 26236 25742 26292
rect 32162 26236 32172 26292
rect 32228 26236 33964 26292
rect 34020 26236 34030 26292
rect 45826 26236 45836 26292
rect 45892 26236 48000 26292
rect 47200 26208 48000 26236
rect 6962 26124 6972 26180
rect 7028 26124 9548 26180
rect 9604 26124 9614 26180
rect 16818 26124 16828 26180
rect 16884 26124 17948 26180
rect 18004 26124 18620 26180
rect 18676 26124 19068 26180
rect 19124 26124 19134 26180
rect 45154 26124 45164 26180
rect 45220 26124 45724 26180
rect 45780 26124 46060 26180
rect 46116 26124 46126 26180
rect 43362 26012 43372 26068
rect 43428 26012 44492 26068
rect 44548 26012 44558 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 4722 25676 4732 25732
rect 4788 25676 6748 25732
rect 6804 25676 6814 25732
rect 8530 25676 8540 25732
rect 8596 25676 8988 25732
rect 9044 25676 9054 25732
rect 4050 25564 4060 25620
rect 4116 25564 12348 25620
rect 12404 25564 12414 25620
rect 28130 25564 28140 25620
rect 28196 25564 30156 25620
rect 30212 25564 30222 25620
rect 47200 25536 48000 25648
rect 8372 25452 9884 25508
rect 9940 25452 9950 25508
rect 11554 25452 11564 25508
rect 11620 25452 12908 25508
rect 12964 25452 13692 25508
rect 13748 25452 14364 25508
rect 14420 25452 15820 25508
rect 15876 25452 15886 25508
rect 24546 25452 24556 25508
rect 24612 25452 25116 25508
rect 25172 25452 25676 25508
rect 25732 25452 25742 25508
rect 32274 25452 32284 25508
rect 32340 25452 34300 25508
rect 34356 25452 34366 25508
rect 38994 25452 39004 25508
rect 39060 25452 40236 25508
rect 40292 25452 40302 25508
rect 8372 25284 8428 25452
rect 12562 25340 12572 25396
rect 12628 25340 13468 25396
rect 13524 25340 13534 25396
rect 26002 25340 26012 25396
rect 26068 25340 28588 25396
rect 28644 25340 29596 25396
rect 29652 25340 29662 25396
rect 41458 25340 41468 25396
rect 41524 25340 42924 25396
rect 42980 25340 42990 25396
rect 43138 25340 43148 25396
rect 43204 25340 43596 25396
rect 43652 25340 43662 25396
rect 4050 25228 4060 25284
rect 4116 25228 8428 25284
rect 12226 25228 12236 25284
rect 12292 25228 14140 25284
rect 14196 25228 14206 25284
rect 20290 25228 20300 25284
rect 20356 25228 20748 25284
rect 20804 25228 22596 25284
rect 32946 25228 32956 25284
rect 33012 25228 36652 25284
rect 36708 25228 37884 25284
rect 37940 25228 38444 25284
rect 38500 25228 38510 25284
rect 38612 25228 42252 25284
rect 42308 25228 42318 25284
rect 22540 25172 22596 25228
rect 38612 25172 38668 25228
rect 22540 25116 23660 25172
rect 23716 25116 23726 25172
rect 35858 25116 35868 25172
rect 35924 25116 36876 25172
rect 36932 25116 37324 25172
rect 37380 25116 37772 25172
rect 37828 25116 38668 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 15362 24892 15372 24948
rect 15428 24892 20972 24948
rect 21028 24892 21038 24948
rect 22082 24892 22092 24948
rect 22148 24892 24780 24948
rect 24836 24892 24846 24948
rect 47200 24864 48000 24976
rect 36978 24780 36988 24836
rect 37044 24780 38556 24836
rect 38612 24780 41020 24836
rect 41076 24780 41086 24836
rect 7634 24668 7644 24724
rect 7700 24668 7980 24724
rect 8036 24668 9324 24724
rect 9380 24668 9390 24724
rect 17490 24668 17500 24724
rect 17556 24668 19964 24724
rect 20020 24668 21196 24724
rect 21252 24668 21262 24724
rect 37538 24668 37548 24724
rect 37604 24668 39676 24724
rect 39732 24668 39742 24724
rect 3490 24556 3500 24612
rect 3556 24556 5964 24612
rect 6020 24556 6030 24612
rect 30370 24556 30380 24612
rect 30436 24556 31052 24612
rect 31108 24556 31118 24612
rect 37090 24556 37100 24612
rect 37156 24556 39452 24612
rect 39508 24556 39518 24612
rect 3500 24388 3556 24556
rect 14914 24444 14924 24500
rect 14980 24444 17500 24500
rect 17556 24444 17566 24500
rect 28018 24444 28028 24500
rect 28084 24444 33964 24500
rect 34020 24444 34030 24500
rect 35522 24444 35532 24500
rect 35588 24444 38108 24500
rect 38164 24444 39116 24500
rect 39172 24444 39182 24500
rect 2034 24332 2044 24388
rect 2100 24332 3556 24388
rect 16370 24332 16380 24388
rect 16436 24332 20188 24388
rect 20244 24332 20254 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 10332 24220 17836 24276
rect 17892 24220 17902 24276
rect 30034 24220 30044 24276
rect 30100 24220 30828 24276
rect 30884 24220 30894 24276
rect 39106 24220 39116 24276
rect 39172 24220 42476 24276
rect 42532 24220 43148 24276
rect 43204 24220 44492 24276
rect 44548 24220 45052 24276
rect 45108 24220 45724 24276
rect 45780 24220 45790 24276
rect 6850 24108 6860 24164
rect 6916 24108 10108 24164
rect 10164 24108 10174 24164
rect 10332 23940 10388 24220
rect 47200 24192 48000 24304
rect 26562 24108 26572 24164
rect 26628 24108 27244 24164
rect 27300 24108 27310 24164
rect 34962 24108 34972 24164
rect 35028 24108 37380 24164
rect 39890 24108 39900 24164
rect 39956 24108 44940 24164
rect 44996 24108 45006 24164
rect 37324 24052 37380 24108
rect 15138 23996 15148 24052
rect 15204 23996 21644 24052
rect 21700 23996 21710 24052
rect 22194 23996 22204 24052
rect 22260 23996 23324 24052
rect 23380 23996 23390 24052
rect 26338 23996 26348 24052
rect 26404 23996 32956 24052
rect 33012 23996 33022 24052
rect 36194 23996 36204 24052
rect 36260 23996 36876 24052
rect 36932 23996 36942 24052
rect 37090 23996 37100 24052
rect 37156 23996 37166 24052
rect 37324 23996 42812 24052
rect 42868 23996 42878 24052
rect 7858 23884 7868 23940
rect 7924 23884 10388 23940
rect 14018 23884 14028 23940
rect 14084 23884 23212 23940
rect 23268 23884 23278 23940
rect 31042 23884 31052 23940
rect 31108 23884 32060 23940
rect 32116 23884 35420 23940
rect 35476 23884 35486 23940
rect 3042 23772 3052 23828
rect 3108 23772 13132 23828
rect 13188 23772 13198 23828
rect 20738 23772 20748 23828
rect 20804 23772 21644 23828
rect 21700 23772 22428 23828
rect 22484 23772 23884 23828
rect 23940 23772 23950 23828
rect 28802 23772 28812 23828
rect 28868 23772 31164 23828
rect 31220 23772 31230 23828
rect 37100 23716 37156 23996
rect 39554 23884 39564 23940
rect 39620 23884 41580 23940
rect 41636 23884 41646 23940
rect 6626 23660 6636 23716
rect 6692 23660 16268 23716
rect 16324 23660 16334 23716
rect 17042 23660 17052 23716
rect 17108 23660 21308 23716
rect 21364 23660 21374 23716
rect 29026 23660 29036 23716
rect 29092 23660 37156 23716
rect 38612 23772 43820 23828
rect 43876 23772 43886 23828
rect 38612 23604 38668 23772
rect 40002 23660 40012 23716
rect 40068 23660 42364 23716
rect 42420 23660 42430 23716
rect 45714 23660 45724 23716
rect 45780 23660 46060 23716
rect 46116 23660 46126 23716
rect 2482 23548 2492 23604
rect 2548 23548 3612 23604
rect 3668 23548 3678 23604
rect 23650 23548 23660 23604
rect 23716 23548 24332 23604
rect 24388 23548 26796 23604
rect 26852 23548 26862 23604
rect 30594 23548 30604 23604
rect 30660 23548 38668 23604
rect 41682 23548 41692 23604
rect 41748 23548 42252 23604
rect 42308 23548 42318 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 47200 23520 48000 23632
rect 13906 23436 13916 23492
rect 13972 23436 15260 23492
rect 15316 23436 15326 23492
rect 2594 23324 2604 23380
rect 2660 23324 3500 23380
rect 3556 23324 3566 23380
rect 34738 23324 34748 23380
rect 34804 23324 38668 23380
rect 38612 23268 38668 23324
rect 19394 23212 19404 23268
rect 19460 23212 20748 23268
rect 20804 23212 20814 23268
rect 23874 23212 23884 23268
rect 23940 23212 24556 23268
rect 24612 23212 26012 23268
rect 26068 23212 26078 23268
rect 28578 23212 28588 23268
rect 28644 23212 33068 23268
rect 33124 23212 33134 23268
rect 38612 23212 40908 23268
rect 40964 23212 40974 23268
rect 41122 23212 41132 23268
rect 41188 23212 41916 23268
rect 41972 23212 41982 23268
rect 41132 23156 41188 23212
rect 2594 23100 2604 23156
rect 2660 23100 5516 23156
rect 5572 23100 5582 23156
rect 26674 23100 26684 23156
rect 26740 23100 31052 23156
rect 31108 23100 32508 23156
rect 32564 23100 33292 23156
rect 33348 23100 33358 23156
rect 39218 23100 39228 23156
rect 39284 23100 40012 23156
rect 40068 23100 41188 23156
rect 8866 22988 8876 23044
rect 8932 22988 9660 23044
rect 9716 22988 12572 23044
rect 12628 22988 12638 23044
rect 16706 22988 16716 23044
rect 16772 22988 17388 23044
rect 17444 22988 17454 23044
rect 18050 22988 18060 23044
rect 18116 22988 19068 23044
rect 19124 22988 19134 23044
rect 21186 22988 21196 23044
rect 21252 22988 23548 23044
rect 23604 22988 23614 23044
rect 32162 22988 32172 23044
rect 32228 22988 34972 23044
rect 35028 22988 35038 23044
rect 2818 22876 2828 22932
rect 2884 22876 6076 22932
rect 6132 22876 6142 22932
rect 11666 22876 11676 22932
rect 11732 22876 13132 22932
rect 13188 22876 13198 22932
rect 47200 22848 48000 22960
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 6738 22652 6748 22708
rect 6804 22652 12796 22708
rect 12852 22652 12862 22708
rect 4050 22428 4060 22484
rect 4116 22428 12684 22484
rect 12740 22428 12750 22484
rect 40002 22428 40012 22484
rect 40068 22428 44828 22484
rect 44884 22428 44894 22484
rect 12562 22316 12572 22372
rect 12628 22316 13804 22372
rect 13860 22316 17780 22372
rect 21410 22316 21420 22372
rect 21476 22316 24444 22372
rect 24500 22316 25004 22372
rect 25060 22316 25070 22372
rect 33170 22316 33180 22372
rect 33236 22316 34412 22372
rect 34468 22316 36876 22372
rect 36932 22316 36942 22372
rect 40786 22316 40796 22372
rect 40852 22316 42028 22372
rect 42084 22316 42094 22372
rect 3042 22204 3052 22260
rect 3108 22204 13020 22260
rect 13076 22204 13086 22260
rect 15026 22204 15036 22260
rect 15092 22204 16380 22260
rect 16436 22204 16446 22260
rect 6066 22092 6076 22148
rect 6132 22092 8428 22148
rect 8484 22092 8494 22148
rect 9202 22092 9212 22148
rect 9268 22092 9278 22148
rect 11554 22092 11564 22148
rect 11620 22092 14476 22148
rect 14532 22092 16716 22148
rect 16772 22092 16782 22148
rect 9212 22036 9268 22092
rect 17724 22036 17780 22316
rect 19394 22204 19404 22260
rect 19460 22204 21868 22260
rect 21924 22204 21934 22260
rect 36642 22204 36652 22260
rect 36708 22204 37996 22260
rect 38052 22204 38062 22260
rect 47200 22176 48000 22288
rect 24882 22092 24892 22148
rect 24948 22092 31948 22148
rect 43810 22092 43820 22148
rect 43876 22092 44828 22148
rect 44884 22092 44894 22148
rect 7746 21980 7756 22036
rect 7812 21980 9268 22036
rect 17714 21980 17724 22036
rect 17780 21980 18172 22036
rect 18228 21980 18238 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 31892 21924 31948 22092
rect 38546 21980 38556 22036
rect 38612 21980 41020 22036
rect 41076 21980 41086 22036
rect 3826 21868 3836 21924
rect 3892 21868 9884 21924
rect 9940 21868 9950 21924
rect 15092 21868 17164 21924
rect 17220 21868 18508 21924
rect 18564 21868 19628 21924
rect 19684 21868 19694 21924
rect 27346 21868 27356 21924
rect 27412 21868 29036 21924
rect 29092 21868 29102 21924
rect 31892 21868 32340 21924
rect 34850 21868 34860 21924
rect 34916 21868 38108 21924
rect 38164 21868 38174 21924
rect 41346 21868 41356 21924
rect 41412 21868 43652 21924
rect 15092 21812 15148 21868
rect 32284 21812 32340 21868
rect 43596 21812 43652 21868
rect 13346 21756 13356 21812
rect 13412 21756 15148 21812
rect 23436 21756 28644 21812
rect 29810 21756 29820 21812
rect 29876 21756 32228 21812
rect 32284 21756 35028 21812
rect 41458 21756 41468 21812
rect 41524 21756 41534 21812
rect 43596 21756 44716 21812
rect 44772 21756 44782 21812
rect 13906 21644 13916 21700
rect 13972 21644 16380 21700
rect 16436 21644 16446 21700
rect 23436 21588 23492 21756
rect 28588 21700 28644 21756
rect 32172 21700 32228 21756
rect 34972 21700 35028 21756
rect 41468 21700 41524 21756
rect 25330 21644 25340 21700
rect 25396 21644 25788 21700
rect 25844 21644 26908 21700
rect 26964 21644 26974 21700
rect 28588 21644 31948 21700
rect 32162 21644 32172 21700
rect 32228 21644 32238 21700
rect 34962 21644 34972 21700
rect 35028 21644 35038 21700
rect 41468 21644 44044 21700
rect 44100 21644 44110 21700
rect 31892 21588 31948 21644
rect 8372 21532 9548 21588
rect 9604 21532 12124 21588
rect 12180 21532 12190 21588
rect 23426 21532 23436 21588
rect 23492 21532 23502 21588
rect 31892 21532 33964 21588
rect 34020 21532 34030 21588
rect 37874 21532 37884 21588
rect 37940 21532 39004 21588
rect 39060 21532 39070 21588
rect 41458 21532 41468 21588
rect 41524 21532 42588 21588
rect 42644 21532 42654 21588
rect 45042 21532 45052 21588
rect 45108 21532 45612 21588
rect 45668 21532 45678 21588
rect 5394 21420 5404 21476
rect 5460 21420 6636 21476
rect 6692 21420 8316 21476
rect 8372 21420 8428 21532
rect 47200 21504 48000 21616
rect 9874 21420 9884 21476
rect 9940 21420 10556 21476
rect 10612 21420 10622 21476
rect 43810 21308 43820 21364
rect 43876 21308 44716 21364
rect 44772 21308 44782 21364
rect 25666 21196 25676 21252
rect 25732 21196 27132 21252
rect 27188 21196 27198 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 21522 20860 21532 20916
rect 21588 20860 23884 20916
rect 23940 20860 23950 20916
rect 26786 20860 26796 20916
rect 26852 20860 27804 20916
rect 27860 20860 28588 20916
rect 28644 20860 30268 20916
rect 30324 20860 31276 20916
rect 31332 20860 31342 20916
rect 47200 20832 48000 20944
rect 17938 20748 17948 20804
rect 18004 20748 20412 20804
rect 20468 20748 23660 20804
rect 23716 20748 23726 20804
rect 37090 20748 37100 20804
rect 37156 20748 37548 20804
rect 37604 20748 40684 20804
rect 40740 20748 40750 20804
rect 41206 20748 41244 20804
rect 41300 20748 41310 20804
rect 3042 20636 3052 20692
rect 3108 20636 9324 20692
rect 9380 20636 9390 20692
rect 3826 20524 3836 20580
rect 3892 20524 6972 20580
rect 7028 20524 7038 20580
rect 20290 20524 20300 20580
rect 20356 20524 21420 20580
rect 21476 20524 21486 20580
rect 36530 20524 36540 20580
rect 36596 20524 37436 20580
rect 37492 20524 37502 20580
rect 43698 20524 43708 20580
rect 43764 20524 44828 20580
rect 44884 20524 44894 20580
rect 44370 20412 44380 20468
rect 44436 20412 46284 20468
rect 46340 20412 46350 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 44818 20300 44828 20356
rect 44884 20300 45724 20356
rect 45780 20300 45790 20356
rect 1810 20188 1820 20244
rect 1876 20188 1886 20244
rect 43362 20188 43372 20244
rect 43428 20188 44492 20244
rect 44548 20188 44558 20244
rect 1820 19908 1876 20188
rect 47200 20160 48000 20272
rect 28130 20076 28140 20132
rect 28196 20076 32060 20132
rect 32116 20076 32126 20132
rect 33618 20076 33628 20132
rect 33684 20076 34076 20132
rect 34132 20076 34142 20132
rect 35858 20076 35868 20132
rect 35924 20076 38892 20132
rect 38948 20076 38958 20132
rect 40450 20076 40460 20132
rect 40516 20076 42924 20132
rect 42980 20076 42990 20132
rect 45714 20076 45724 20132
rect 45780 20076 45790 20132
rect 45724 20020 45780 20076
rect 7634 19964 7644 20020
rect 7700 19964 8540 20020
rect 8596 19964 8606 20020
rect 10658 19964 10668 20020
rect 10724 19964 12460 20020
rect 12516 19964 12526 20020
rect 17826 19964 17836 20020
rect 17892 19964 20860 20020
rect 20916 19964 20926 20020
rect 28466 19964 28476 20020
rect 28532 19964 33068 20020
rect 33124 19964 33134 20020
rect 33282 19964 33292 20020
rect 33348 19964 33964 20020
rect 34020 19964 34030 20020
rect 37986 19964 37996 20020
rect 38052 19964 45780 20020
rect 1820 19852 10220 19908
rect 10276 19852 10286 19908
rect 23090 19852 23100 19908
rect 23156 19852 25228 19908
rect 25284 19852 25294 19908
rect 26002 19852 26012 19908
rect 26068 19852 31052 19908
rect 31108 19852 31118 19908
rect 31892 19852 33740 19908
rect 33796 19852 33806 19908
rect 36194 19852 36204 19908
rect 36260 19852 39228 19908
rect 39284 19852 39294 19908
rect 41906 19852 41916 19908
rect 41972 19852 41982 19908
rect 31892 19796 31948 19852
rect 41916 19796 41972 19852
rect 28018 19740 28028 19796
rect 28084 19740 31948 19796
rect 34972 19740 41972 19796
rect 6066 19628 6076 19684
rect 6132 19628 6748 19684
rect 6804 19628 6814 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 34972 19572 35028 19740
rect 38322 19628 38332 19684
rect 38388 19628 39788 19684
rect 39844 19628 42924 19684
rect 42980 19628 45052 19684
rect 45108 19628 45118 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 47200 19572 48000 19600
rect 1922 19516 1932 19572
rect 1988 19516 2492 19572
rect 2548 19516 2558 19572
rect 20290 19516 20300 19572
rect 20356 19516 20748 19572
rect 20804 19516 20814 19572
rect 25106 19516 25116 19572
rect 25172 19516 35028 19572
rect 46162 19516 46172 19572
rect 46228 19516 48000 19572
rect 47200 19488 48000 19516
rect 14802 19404 14812 19460
rect 14868 19404 15820 19460
rect 15876 19404 15886 19460
rect 29138 19404 29148 19460
rect 29204 19404 30044 19460
rect 30100 19404 30110 19460
rect 3938 19292 3948 19348
rect 4004 19292 5964 19348
rect 6020 19292 6030 19348
rect 16370 19292 16380 19348
rect 16436 19292 19852 19348
rect 19908 19292 19918 19348
rect 27570 19292 27580 19348
rect 27636 19292 31052 19348
rect 31108 19292 31118 19348
rect 31938 19292 31948 19348
rect 32004 19292 33292 19348
rect 33348 19292 34636 19348
rect 34692 19292 35980 19348
rect 36036 19292 36046 19348
rect 39890 19292 39900 19348
rect 39956 19292 43820 19348
rect 43876 19292 43886 19348
rect 13692 19180 14364 19236
rect 14420 19180 14924 19236
rect 14980 19180 14990 19236
rect 25778 19180 25788 19236
rect 25844 19180 28588 19236
rect 28644 19180 29260 19236
rect 29316 19180 29326 19236
rect 32498 19180 32508 19236
rect 32564 19180 33516 19236
rect 33572 19180 33582 19236
rect 13692 19124 13748 19180
rect 2258 19068 2268 19124
rect 2324 19068 5964 19124
rect 6020 19068 6030 19124
rect 11442 19068 11452 19124
rect 11508 19068 12236 19124
rect 12292 19068 12302 19124
rect 12562 19068 12572 19124
rect 12628 19068 13692 19124
rect 13748 19068 13758 19124
rect 14130 19068 14140 19124
rect 14196 19068 14206 19124
rect 32722 19068 32732 19124
rect 32788 19068 42140 19124
rect 42196 19068 42206 19124
rect 46050 19068 46060 19124
rect 46116 19068 46126 19124
rect 14140 18900 14196 19068
rect 15922 18956 15932 19012
rect 15988 18956 19180 19012
rect 19236 18956 19246 19012
rect 20514 18956 20524 19012
rect 20580 18956 22316 19012
rect 22372 18956 22382 19012
rect 32274 18956 32284 19012
rect 32340 18956 36092 19012
rect 36148 18956 36158 19012
rect 38612 18956 41132 19012
rect 41188 18956 41198 19012
rect 8194 18844 8204 18900
rect 8260 18844 14196 18900
rect 32162 18844 32172 18900
rect 32228 18844 34412 18900
rect 34468 18844 34478 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 38612 18788 38668 18956
rect 46060 18900 46116 19068
rect 47200 18900 48000 18928
rect 46060 18844 48000 18900
rect 47200 18816 48000 18844
rect 29810 18732 29820 18788
rect 29876 18732 38668 18788
rect 9202 18620 9212 18676
rect 9268 18620 11228 18676
rect 11284 18620 11294 18676
rect 18834 18620 18844 18676
rect 18900 18620 20300 18676
rect 20356 18620 20366 18676
rect 28914 18620 28924 18676
rect 28980 18620 31276 18676
rect 31332 18620 31342 18676
rect 37314 18620 37324 18676
rect 37380 18620 40124 18676
rect 40180 18620 40190 18676
rect 44034 18620 44044 18676
rect 44100 18620 44492 18676
rect 44548 18620 44940 18676
rect 44996 18620 45006 18676
rect 1698 18508 1708 18564
rect 1764 18508 3388 18564
rect 3444 18508 3454 18564
rect 7970 18508 7980 18564
rect 8036 18508 9436 18564
rect 9492 18508 9502 18564
rect 12114 18508 12124 18564
rect 12180 18508 13468 18564
rect 13524 18508 13534 18564
rect 29698 18508 29708 18564
rect 29764 18508 30604 18564
rect 30660 18508 30670 18564
rect 33842 18508 33852 18564
rect 33908 18508 35644 18564
rect 35700 18508 35710 18564
rect 37650 18508 37660 18564
rect 37716 18508 38892 18564
rect 38948 18508 38958 18564
rect 41570 18508 41580 18564
rect 41636 18508 45724 18564
rect 45780 18508 45790 18564
rect 16258 18396 16268 18452
rect 16324 18396 17836 18452
rect 17892 18396 17902 18452
rect 18162 18396 18172 18452
rect 18228 18396 18620 18452
rect 18676 18396 19628 18452
rect 19684 18396 19694 18452
rect 20850 18396 20860 18452
rect 20916 18396 20926 18452
rect 22530 18396 22540 18452
rect 22596 18396 23660 18452
rect 23716 18396 24332 18452
rect 24388 18396 25340 18452
rect 25396 18396 25406 18452
rect 26898 18396 26908 18452
rect 26964 18396 31724 18452
rect 31780 18396 31790 18452
rect 36978 18396 36988 18452
rect 37044 18396 39452 18452
rect 39508 18396 40348 18452
rect 40404 18396 40414 18452
rect 15698 18284 15708 18340
rect 15764 18284 16716 18340
rect 16772 18284 16782 18340
rect 18946 18284 18956 18340
rect 19012 18284 19852 18340
rect 19908 18284 19918 18340
rect 20860 18228 20916 18396
rect 31378 18284 31388 18340
rect 31444 18284 31948 18340
rect 32004 18284 32014 18340
rect 37314 18284 37324 18340
rect 37380 18284 38556 18340
rect 38612 18284 41356 18340
rect 41412 18284 41422 18340
rect 42466 18284 42476 18340
rect 42532 18284 44716 18340
rect 44772 18284 44782 18340
rect 47200 18228 48000 18256
rect 3042 18172 3052 18228
rect 3108 18172 5404 18228
rect 5460 18172 5470 18228
rect 20860 18172 25676 18228
rect 25732 18172 28252 18228
rect 28308 18172 32508 18228
rect 32564 18172 32574 18228
rect 40898 18172 40908 18228
rect 40964 18172 42028 18228
rect 42084 18172 42094 18228
rect 46050 18172 46060 18228
rect 46116 18172 48000 18228
rect 47200 18144 48000 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 8642 17948 8652 18004
rect 8708 17948 9884 18004
rect 9940 17948 9950 18004
rect 21858 17724 21868 17780
rect 21924 17724 22540 17780
rect 22596 17724 22606 17780
rect 30258 17724 30268 17780
rect 30324 17724 34076 17780
rect 34132 17724 35308 17780
rect 35364 17724 35374 17780
rect 8082 17612 8092 17668
rect 8148 17612 9212 17668
rect 9268 17612 9278 17668
rect 10210 17612 10220 17668
rect 10276 17612 13468 17668
rect 13524 17612 13534 17668
rect 14914 17612 14924 17668
rect 14980 17612 16940 17668
rect 16996 17612 19180 17668
rect 19236 17612 20188 17668
rect 20244 17612 21084 17668
rect 21140 17612 22764 17668
rect 22820 17612 22830 17668
rect 0 17556 800 17584
rect 47200 17556 48000 17584
rect 0 17500 3500 17556
rect 3556 17500 3566 17556
rect 11442 17500 11452 17556
rect 11508 17500 13580 17556
rect 13636 17500 13646 17556
rect 21522 17500 21532 17556
rect 21588 17500 22428 17556
rect 22484 17500 22494 17556
rect 25330 17500 25340 17556
rect 25396 17500 27020 17556
rect 27076 17500 27580 17556
rect 27636 17500 27646 17556
rect 33618 17500 33628 17556
rect 33684 17500 35084 17556
rect 35140 17500 35150 17556
rect 38612 17500 44268 17556
rect 44324 17500 44940 17556
rect 44996 17500 45006 17556
rect 46050 17500 46060 17556
rect 46116 17500 48000 17556
rect 0 17472 800 17500
rect 38612 17444 38668 17500
rect 47200 17472 48000 17500
rect 6626 17388 6636 17444
rect 6692 17388 9772 17444
rect 9828 17388 9838 17444
rect 13010 17388 13020 17444
rect 13076 17388 14364 17444
rect 14420 17388 14430 17444
rect 31892 17388 38668 17444
rect 40786 17388 40796 17444
rect 40852 17388 42140 17444
rect 42196 17388 42206 17444
rect 31892 17332 31948 17388
rect 31714 17276 31724 17332
rect 31780 17276 31948 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 18274 17164 18284 17220
rect 18340 17164 19068 17220
rect 19124 17164 19134 17220
rect 8978 17052 8988 17108
rect 9044 17052 10108 17108
rect 10164 17052 10174 17108
rect 16370 17052 16380 17108
rect 16436 17052 17724 17108
rect 17780 17052 17790 17108
rect 43810 17052 43820 17108
rect 43876 17052 44940 17108
rect 44996 17052 45006 17108
rect 2034 16940 2044 16996
rect 2100 16940 10220 16996
rect 10276 16940 10286 16996
rect 18050 16940 18060 16996
rect 18116 16940 18956 16996
rect 19012 16940 19022 16996
rect 35746 16940 35756 16996
rect 35812 16940 36204 16996
rect 36260 16940 36270 16996
rect 36614 16940 36652 16996
rect 36708 16940 36718 16996
rect 41122 16940 41132 16996
rect 41188 16940 43708 16996
rect 43764 16940 43774 16996
rect 44482 16940 44492 16996
rect 44548 16940 46508 16996
rect 46564 16940 46574 16996
rect 47200 16884 48000 16912
rect 4946 16828 4956 16884
rect 5012 16828 9436 16884
rect 9492 16828 9502 16884
rect 10658 16828 10668 16884
rect 10724 16828 12460 16884
rect 12516 16828 12526 16884
rect 14130 16828 14140 16884
rect 14196 16828 15148 16884
rect 15204 16828 15214 16884
rect 28914 16828 28924 16884
rect 28980 16828 29596 16884
rect 29652 16828 30492 16884
rect 30548 16828 30558 16884
rect 33170 16828 33180 16884
rect 33236 16828 36764 16884
rect 36820 16828 36830 16884
rect 40562 16828 40572 16884
rect 40628 16828 41020 16884
rect 41076 16828 41356 16884
rect 41412 16828 44380 16884
rect 44436 16828 44446 16884
rect 46050 16828 46060 16884
rect 46116 16828 48000 16884
rect 47200 16800 48000 16828
rect 13682 16716 13692 16772
rect 13748 16716 14812 16772
rect 14868 16716 14878 16772
rect 34178 16716 34188 16772
rect 34244 16716 36316 16772
rect 36372 16716 36382 16772
rect 39442 16716 39452 16772
rect 39508 16716 45500 16772
rect 45556 16716 45566 16772
rect 6962 16604 6972 16660
rect 7028 16604 9100 16660
rect 9156 16604 9166 16660
rect 22866 16604 22876 16660
rect 22932 16604 23660 16660
rect 23716 16604 23726 16660
rect 24770 16604 24780 16660
rect 24836 16604 26236 16660
rect 26292 16604 26302 16660
rect 34738 16604 34748 16660
rect 34804 16604 38332 16660
rect 38388 16604 38398 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16258 16380 16268 16436
rect 16324 16380 17500 16436
rect 17556 16380 17566 16436
rect 4834 16268 4844 16324
rect 4900 16268 10444 16324
rect 10500 16268 10510 16324
rect 15026 16268 15036 16324
rect 15092 16268 16828 16324
rect 16884 16268 16894 16324
rect 47200 16212 48000 16240
rect 14018 16156 14028 16212
rect 14084 16156 15484 16212
rect 15540 16156 15550 16212
rect 45490 16156 45500 16212
rect 45556 16156 48000 16212
rect 47200 16128 48000 16156
rect 8372 16044 8540 16100
rect 8596 16044 9212 16100
rect 9268 16044 9278 16100
rect 14578 16044 14588 16100
rect 14644 16044 15260 16100
rect 15316 16044 15326 16100
rect 23986 16044 23996 16100
rect 24052 16044 24892 16100
rect 24948 16044 25116 16100
rect 25172 16044 28924 16100
rect 28980 16044 28990 16100
rect 34850 16044 34860 16100
rect 34916 16044 35868 16100
rect 35924 16044 35934 16100
rect 36530 16044 36540 16100
rect 36596 16044 37324 16100
rect 37380 16044 37390 16100
rect 8372 15876 8428 16044
rect 17826 15932 17836 15988
rect 17892 15932 18620 15988
rect 18676 15932 18686 15988
rect 21746 15932 21756 15988
rect 21812 15932 22652 15988
rect 22708 15932 22718 15988
rect 6290 15820 6300 15876
rect 6356 15820 8428 15876
rect 12338 15820 12348 15876
rect 12404 15820 12908 15876
rect 12964 15820 13692 15876
rect 13748 15820 14028 15876
rect 14084 15820 14094 15876
rect 23426 15820 23436 15876
rect 23492 15820 25116 15876
rect 25172 15820 25182 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 12674 15596 12684 15652
rect 12740 15596 13580 15652
rect 13636 15596 13646 15652
rect 24658 15596 24668 15652
rect 24724 15596 26012 15652
rect 26068 15596 26078 15652
rect 47200 15540 48000 15568
rect 8306 15484 8316 15540
rect 8372 15428 8428 15540
rect 9202 15484 9212 15540
rect 9268 15484 9996 15540
rect 10052 15484 10332 15540
rect 10388 15484 13020 15540
rect 13076 15484 13086 15540
rect 17154 15484 17164 15540
rect 17220 15484 19740 15540
rect 19796 15484 19806 15540
rect 25890 15484 25900 15540
rect 25956 15484 28140 15540
rect 28196 15484 28206 15540
rect 30146 15484 30156 15540
rect 30212 15484 31612 15540
rect 31668 15484 31678 15540
rect 38770 15484 38780 15540
rect 38836 15484 39676 15540
rect 39732 15484 39742 15540
rect 45490 15484 45500 15540
rect 45556 15484 48000 15540
rect 47200 15456 48000 15484
rect 8372 15372 9548 15428
rect 9604 15372 9614 15428
rect 26450 15372 26460 15428
rect 26516 15372 26908 15428
rect 39218 15372 39228 15428
rect 39284 15372 45388 15428
rect 45444 15372 45454 15428
rect 5058 15260 5068 15316
rect 5124 15260 5740 15316
rect 5796 15260 5806 15316
rect 26852 15204 26908 15372
rect 28914 15260 28924 15316
rect 28980 15260 29708 15316
rect 29764 15260 29774 15316
rect 41122 15260 41132 15316
rect 41188 15260 45612 15316
rect 45668 15260 45678 15316
rect 7970 15148 7980 15204
rect 8036 15148 8876 15204
rect 8932 15148 8942 15204
rect 9874 15148 9884 15204
rect 9940 15148 10780 15204
rect 10836 15148 12348 15204
rect 12404 15148 12414 15204
rect 20290 15148 20300 15204
rect 20356 15148 26236 15204
rect 26292 15148 26302 15204
rect 26852 15148 27916 15204
rect 27972 15148 27982 15204
rect 33506 15148 33516 15204
rect 33572 15148 34748 15204
rect 34804 15148 34814 15204
rect 37650 15148 37660 15204
rect 37716 15148 40236 15204
rect 40292 15148 40302 15204
rect 41206 15148 41244 15204
rect 41300 15148 41310 15204
rect 7858 15036 7868 15092
rect 7924 15036 8988 15092
rect 9044 15036 9054 15092
rect 22866 15036 22876 15092
rect 22932 15036 23884 15092
rect 23940 15036 23950 15092
rect 24882 15036 24892 15092
rect 24948 15036 27244 15092
rect 27300 15036 27310 15092
rect 32386 15036 32396 15092
rect 32452 15036 34300 15092
rect 34356 15036 34366 15092
rect 38434 15036 38444 15092
rect 38500 15036 39788 15092
rect 39844 15036 40908 15092
rect 40964 15036 40974 15092
rect 32722 14924 32732 14980
rect 32788 14924 33964 14980
rect 34020 14924 34030 14980
rect 41906 14924 41916 14980
rect 41972 14924 45388 14980
rect 45444 14924 45454 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 47200 14868 48000 14896
rect 8418 14812 8428 14868
rect 8484 14812 9884 14868
rect 9940 14812 9950 14868
rect 33394 14812 33404 14868
rect 33460 14812 34636 14868
rect 34692 14812 34702 14868
rect 45714 14812 45724 14868
rect 45780 14812 48000 14868
rect 47200 14784 48000 14812
rect 1586 14700 1596 14756
rect 1652 14700 6524 14756
rect 6580 14700 6590 14756
rect 31154 14700 31164 14756
rect 31220 14700 32396 14756
rect 32452 14700 32462 14756
rect 33282 14700 33292 14756
rect 33348 14700 35644 14756
rect 35700 14700 35710 14756
rect 23874 14588 23884 14644
rect 23940 14588 24220 14644
rect 24276 14588 24286 14644
rect 32162 14588 32172 14644
rect 32228 14588 33068 14644
rect 33124 14588 33134 14644
rect 33730 14588 33740 14644
rect 33796 14588 35420 14644
rect 35476 14588 35486 14644
rect 45938 14588 45948 14644
rect 46004 14588 46620 14644
rect 46676 14588 46686 14644
rect 35186 14364 35196 14420
rect 35252 14364 35756 14420
rect 35812 14364 35822 14420
rect 45938 14364 45948 14420
rect 46004 14364 46014 14420
rect 1922 14252 1932 14308
rect 1988 14252 2716 14308
rect 2772 14252 3164 14308
rect 3220 14252 3230 14308
rect 32834 14252 32844 14308
rect 32900 14252 33740 14308
rect 33796 14252 33806 14308
rect 36306 14252 36316 14308
rect 36372 14252 37548 14308
rect 37604 14252 37614 14308
rect 45948 14196 46004 14364
rect 47200 14196 48000 14224
rect 45948 14140 48000 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 47200 14112 48000 14140
rect 2370 13916 2380 13972
rect 2436 13916 4844 13972
rect 4900 13916 4910 13972
rect 16818 13916 16828 13972
rect 16884 13916 18396 13972
rect 18452 13916 18462 13972
rect 26114 13804 26124 13860
rect 26180 13804 28028 13860
rect 28084 13804 28094 13860
rect 32498 13804 32508 13860
rect 32564 13804 33404 13860
rect 33460 13804 34076 13860
rect 34132 13804 34524 13860
rect 34580 13804 34590 13860
rect 37090 13804 37100 13860
rect 37156 13804 42476 13860
rect 42532 13804 42542 13860
rect 43474 13804 43484 13860
rect 43540 13804 44380 13860
rect 44436 13804 44446 13860
rect 34524 13636 34580 13804
rect 3154 13580 3164 13636
rect 3220 13580 5852 13636
rect 5908 13580 8428 13636
rect 8484 13580 8494 13636
rect 20850 13580 20860 13636
rect 20916 13580 22988 13636
rect 23044 13580 23054 13636
rect 29810 13580 29820 13636
rect 29876 13580 33292 13636
rect 33348 13580 33358 13636
rect 34524 13580 34860 13636
rect 34916 13580 34926 13636
rect 43810 13580 43820 13636
rect 43876 13580 44828 13636
rect 44884 13580 44894 13636
rect 47200 13524 48000 13552
rect 1810 13468 1820 13524
rect 1876 13468 5068 13524
rect 5124 13468 5134 13524
rect 35970 13468 35980 13524
rect 36036 13468 37436 13524
rect 37492 13468 37502 13524
rect 40002 13468 40012 13524
rect 40068 13468 41132 13524
rect 41188 13468 41198 13524
rect 43586 13468 43596 13524
rect 43652 13468 48000 13524
rect 47200 13440 48000 13468
rect 7746 13356 7756 13412
rect 7812 13356 8764 13412
rect 8820 13356 8830 13412
rect 9426 13356 9436 13412
rect 9492 13356 11788 13412
rect 11844 13356 11854 13412
rect 24994 13356 25004 13412
rect 25060 13356 27580 13412
rect 27636 13356 27646 13412
rect 32610 13356 32620 13412
rect 32676 13356 34412 13412
rect 34468 13356 34478 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 4386 13132 4396 13188
rect 4452 13132 6972 13188
rect 7028 13132 7038 13188
rect 30370 13132 30380 13188
rect 30436 13132 32732 13188
rect 32788 13132 32798 13188
rect 5618 13020 5628 13076
rect 5684 13020 9324 13076
rect 9380 13020 9390 13076
rect 14354 13020 14364 13076
rect 14420 13020 19292 13076
rect 19348 13020 19358 13076
rect 34850 13020 34860 13076
rect 34916 13020 35868 13076
rect 35924 13020 35934 13076
rect 43708 13020 46452 13076
rect 43708 12852 43764 13020
rect 1474 12796 1484 12852
rect 1540 12796 2380 12852
rect 2436 12796 2446 12852
rect 35970 12796 35980 12852
rect 36036 12796 39116 12852
rect 39172 12796 39182 12852
rect 43250 12796 43260 12852
rect 43316 12796 43764 12852
rect 43820 12908 45052 12964
rect 45108 12908 46172 12964
rect 46228 12908 46238 12964
rect 43820 12740 43876 12908
rect 46396 12852 46452 13020
rect 47200 12852 48000 12880
rect 46396 12796 48000 12852
rect 47200 12768 48000 12796
rect 28466 12684 28476 12740
rect 28532 12684 43876 12740
rect 44258 12684 44268 12740
rect 44324 12684 44334 12740
rect 44268 12628 44324 12684
rect 2594 12572 2604 12628
rect 2660 12572 3500 12628
rect 3556 12572 3566 12628
rect 5506 12572 5516 12628
rect 5572 12572 6748 12628
rect 6804 12572 6814 12628
rect 28578 12572 28588 12628
rect 28644 12572 43036 12628
rect 43092 12572 44324 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 8642 12460 8652 12516
rect 8708 12460 10556 12516
rect 10612 12460 10622 12516
rect 27458 12236 27468 12292
rect 27524 12236 30380 12292
rect 30436 12236 30446 12292
rect 40338 12236 40348 12292
rect 40404 12236 42924 12292
rect 42980 12236 42990 12292
rect 47200 12180 48000 12208
rect 43586 12124 43596 12180
rect 43652 12124 48000 12180
rect 47200 12096 48000 12124
rect 9650 12012 9660 12068
rect 9716 12012 12012 12068
rect 12068 12012 12078 12068
rect 28242 12012 28252 12068
rect 28308 12012 29372 12068
rect 29428 12012 29438 12068
rect 33842 12012 33852 12068
rect 33908 12012 35084 12068
rect 35140 12012 35150 12068
rect 40114 12012 40124 12068
rect 40180 12012 41916 12068
rect 41972 12012 41982 12068
rect 2034 11900 2044 11956
rect 2100 11900 4284 11956
rect 4340 11900 4350 11956
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 29250 11676 29260 11732
rect 29316 11676 31948 11732
rect 36866 11676 36876 11732
rect 36932 11676 39340 11732
rect 39396 11676 39406 11732
rect 41346 11676 41356 11732
rect 41412 11676 42028 11732
rect 42084 11676 42094 11732
rect 31892 11508 31948 11676
rect 32386 11564 32396 11620
rect 32452 11564 38052 11620
rect 37996 11508 38052 11564
rect 47200 11508 48000 11536
rect 29586 11452 29596 11508
rect 29652 11452 30492 11508
rect 30548 11452 30558 11508
rect 31892 11452 33404 11508
rect 33460 11452 33470 11508
rect 37986 11452 37996 11508
rect 38052 11452 38062 11508
rect 41346 11452 41356 11508
rect 41412 11452 42252 11508
rect 42308 11452 42318 11508
rect 45602 11452 45612 11508
rect 45668 11452 48000 11508
rect 47200 11424 48000 11452
rect 1586 11228 1596 11284
rect 1652 11228 2380 11284
rect 2436 11228 2446 11284
rect 39666 11228 39676 11284
rect 39732 11228 43932 11284
rect 43988 11228 43998 11284
rect 37090 11116 37100 11172
rect 37156 11116 44940 11172
rect 44996 11116 45006 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 47200 10836 48000 10864
rect 33842 10780 33852 10836
rect 33908 10780 43708 10836
rect 44034 10780 44044 10836
rect 44100 10780 44828 10836
rect 44884 10780 48000 10836
rect 43652 10724 43708 10780
rect 47200 10752 48000 10780
rect 32946 10668 32956 10724
rect 33012 10668 35420 10724
rect 35476 10668 35486 10724
rect 36530 10668 36540 10724
rect 36596 10668 38668 10724
rect 38724 10668 38734 10724
rect 43652 10668 45724 10724
rect 45780 10668 45790 10724
rect 24434 10444 24444 10500
rect 24500 10444 26572 10500
rect 26628 10444 26638 10500
rect 33730 10444 33740 10500
rect 33796 10444 34412 10500
rect 34468 10444 34478 10500
rect 42130 10332 42140 10388
rect 42196 10332 42476 10388
rect 42532 10332 42542 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 47200 10164 48000 10192
rect 42466 10108 42476 10164
rect 42532 10108 43820 10164
rect 43876 10108 43886 10164
rect 45490 10108 45500 10164
rect 45556 10108 46060 10164
rect 46116 10108 48000 10164
rect 47200 10080 48000 10108
rect 24098 9996 24108 10052
rect 24164 9996 28588 10052
rect 28644 9996 28654 10052
rect 36642 9996 36652 10052
rect 36708 9996 42140 10052
rect 42196 9996 42206 10052
rect 43586 9996 43596 10052
rect 43652 9996 45388 10052
rect 45444 9996 45454 10052
rect 33394 9772 33404 9828
rect 33460 9772 37100 9828
rect 37156 9772 37166 9828
rect 5282 9660 5292 9716
rect 5348 9660 9212 9716
rect 9268 9660 9278 9716
rect 38546 9548 38556 9604
rect 38612 9548 44940 9604
rect 44996 9548 45006 9604
rect 47200 9492 48000 9520
rect 43586 9436 43596 9492
rect 43652 9436 43932 9492
rect 43988 9436 48000 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 47200 9408 48000 9436
rect 33506 9100 33516 9156
rect 33572 9100 35644 9156
rect 35700 9100 35710 9156
rect 33618 8988 33628 9044
rect 33684 8988 43260 9044
rect 43316 8988 43326 9044
rect 44678 8876 44716 8932
rect 44772 8876 44782 8932
rect 47200 8820 48000 8848
rect 44258 8764 44268 8820
rect 44324 8764 48000 8820
rect 47200 8736 48000 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 31714 8316 31724 8372
rect 31780 8316 32844 8372
rect 32900 8316 32910 8372
rect 47200 8148 48000 8176
rect 46050 8092 46060 8148
rect 46116 8092 48000 8148
rect 47200 8064 48000 8092
rect 2818 7980 2828 8036
rect 2884 7980 3388 8036
rect 3444 7980 18396 8036
rect 18452 7980 18462 8036
rect 25218 7980 25228 8036
rect 25284 7980 43932 8036
rect 43988 7980 43998 8036
rect 44930 7980 44940 8036
rect 44996 7980 45006 8036
rect 44940 7924 44996 7980
rect 30258 7868 30268 7924
rect 30324 7868 44996 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 0 7476 800 7504
rect 47200 7476 48000 7504
rect 0 7420 2044 7476
rect 2100 7420 2110 7476
rect 37090 7420 37100 7476
rect 37156 7420 44940 7476
rect 44996 7420 45006 7476
rect 45714 7420 45724 7476
rect 45780 7420 48000 7476
rect 0 7392 800 7420
rect 47200 7392 48000 7420
rect 2930 7308 2940 7364
rect 2996 7308 3500 7364
rect 3556 7308 22204 7364
rect 22260 7308 22270 7364
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 31266 6972 31276 7028
rect 31332 6972 33628 7028
rect 33684 6972 33694 7028
rect 0 6804 800 6832
rect 47200 6804 48000 6832
rect 0 6748 1932 6804
rect 1988 6748 1998 6804
rect 34178 6748 34188 6804
rect 34244 6748 38556 6804
rect 38612 6748 38622 6804
rect 44370 6748 44380 6804
rect 44436 6748 45276 6804
rect 45332 6748 45342 6804
rect 45612 6748 48000 6804
rect 0 6720 800 6748
rect 45612 6692 45668 6748
rect 47200 6720 48000 6748
rect 2930 6636 2940 6692
rect 2996 6636 16604 6692
rect 16660 6636 16670 6692
rect 45602 6636 45612 6692
rect 45668 6636 45678 6692
rect 44034 6524 44044 6580
rect 44100 6524 45836 6580
rect 45892 6524 45902 6580
rect 38546 6412 38556 6468
rect 38612 6412 44940 6468
rect 44996 6412 45006 6468
rect 2146 6300 2156 6356
rect 2212 6300 18620 6356
rect 18676 6300 18686 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 0 6132 800 6160
rect 47200 6132 48000 6160
rect 0 6076 2044 6132
rect 2100 6076 2110 6132
rect 23874 6076 23884 6132
rect 23940 6076 24444 6132
rect 24500 6076 25228 6132
rect 25284 6076 25294 6132
rect 32610 6076 32620 6132
rect 32676 6076 33852 6132
rect 33908 6076 33918 6132
rect 46162 6076 46172 6132
rect 46228 6076 48000 6132
rect 0 6048 800 6076
rect 47200 6048 48000 6076
rect 8372 5964 20748 6020
rect 20804 5964 20814 6020
rect 8372 5908 8428 5964
rect 2930 5852 2940 5908
rect 2996 5852 8428 5908
rect 21634 5852 21644 5908
rect 21700 5852 22428 5908
rect 22484 5852 22494 5908
rect 18274 5740 18284 5796
rect 18340 5740 20412 5796
rect 20468 5740 20972 5796
rect 21028 5740 21038 5796
rect 28242 5740 28252 5796
rect 28308 5740 28812 5796
rect 28868 5740 42364 5796
rect 42420 5740 42430 5796
rect 8866 5628 8876 5684
rect 8932 5628 23660 5684
rect 23716 5628 23726 5684
rect 27010 5628 27020 5684
rect 27076 5628 43820 5684
rect 43876 5628 43886 5684
rect 10546 5516 10556 5572
rect 10612 5516 22204 5572
rect 22260 5516 22270 5572
rect 0 5460 800 5488
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 47200 5460 48000 5488
rect 0 5404 1932 5460
rect 1988 5404 1998 5460
rect 45490 5404 45500 5460
rect 45556 5404 46172 5460
rect 46228 5404 48000 5460
rect 0 5376 800 5404
rect 47200 5376 48000 5404
rect 10098 5292 10108 5348
rect 10164 5292 23100 5348
rect 23156 5292 23166 5348
rect 12562 5180 12572 5236
rect 12628 5180 14700 5236
rect 14756 5180 14766 5236
rect 18498 5180 18508 5236
rect 18564 5180 22988 5236
rect 23044 5180 23054 5236
rect 8372 5068 13692 5124
rect 13748 5068 13758 5124
rect 14802 5068 14812 5124
rect 14868 5068 15596 5124
rect 15652 5068 15662 5124
rect 16370 5068 16380 5124
rect 16436 5068 17500 5124
rect 17556 5068 18060 5124
rect 18116 5068 18126 5124
rect 18396 5068 22764 5124
rect 22820 5068 22830 5124
rect 23426 5068 23436 5124
rect 23492 5068 24444 5124
rect 24500 5068 24510 5124
rect 40338 5068 40348 5124
rect 40404 5068 44940 5124
rect 44996 5068 45006 5124
rect 8372 5012 8428 5068
rect 18396 5012 18452 5068
rect 2146 4956 2156 5012
rect 2212 4956 8428 5012
rect 11778 4956 11788 5012
rect 11844 4956 18452 5012
rect 21746 4956 21756 5012
rect 21812 4956 22652 5012
rect 22708 4956 22718 5012
rect 33394 4956 33404 5012
rect 33460 4956 37100 5012
rect 37156 4956 37166 5012
rect 31490 4844 31500 4900
rect 31556 4844 37212 4900
rect 37268 4844 37278 4900
rect 39330 4844 39340 4900
rect 39396 4844 41356 4900
rect 41412 4844 41422 4900
rect 43586 4844 43596 4900
rect 0 4788 800 4816
rect 43652 4788 43708 4900
rect 47200 4788 48000 4816
rect 0 4732 1708 4788
rect 1764 4732 2492 4788
rect 2548 4732 2558 4788
rect 26450 4732 26460 4788
rect 26516 4732 28588 4788
rect 28644 4732 28654 4788
rect 34066 4732 34076 4788
rect 34132 4732 42252 4788
rect 42308 4732 42318 4788
rect 43652 4732 48000 4788
rect 0 4704 800 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 47200 4704 48000 4732
rect 17714 4508 17724 4564
rect 17780 4508 23212 4564
rect 23268 4508 23278 4564
rect 26226 4508 26236 4564
rect 26292 4508 28028 4564
rect 28084 4508 28094 4564
rect 33842 4508 33852 4564
rect 33908 4508 35420 4564
rect 35476 4508 36428 4564
rect 36484 4508 36494 4564
rect 40114 4508 40124 4564
rect 40180 4508 40908 4564
rect 40964 4508 40974 4564
rect 20066 4396 20076 4452
rect 20132 4396 20412 4452
rect 20468 4396 20478 4452
rect 29362 4396 29372 4452
rect 29428 4396 31164 4452
rect 31220 4396 31230 4452
rect 33058 4396 33068 4452
rect 33124 4396 35868 4452
rect 35924 4396 35934 4452
rect 44146 4396 44156 4452
rect 44212 4396 45836 4452
rect 45892 4396 45902 4452
rect 24210 4284 24220 4340
rect 24276 4284 31948 4340
rect 33170 4284 33180 4340
rect 33236 4284 34748 4340
rect 34804 4284 34814 4340
rect 31892 4228 31948 4284
rect 2034 4172 2044 4228
rect 2100 4172 18284 4228
rect 18340 4172 18350 4228
rect 26226 4172 26236 4228
rect 26292 4172 27188 4228
rect 31892 4172 34356 4228
rect 34850 4172 34860 4228
rect 34916 4172 36652 4228
rect 36708 4172 36718 4228
rect 42354 4172 42364 4228
rect 42420 4172 45612 4228
rect 45668 4172 45678 4228
rect 0 4116 800 4144
rect 27132 4116 27188 4172
rect 34300 4116 34356 4172
rect 47200 4116 48000 4144
rect 0 4060 1708 4116
rect 1764 4060 2492 4116
rect 2548 4060 2558 4116
rect 27122 4060 27132 4116
rect 27188 4060 27198 4116
rect 33282 4060 33292 4116
rect 33348 4060 34076 4116
rect 34132 4060 34142 4116
rect 34300 4060 41916 4116
rect 41972 4060 41982 4116
rect 43586 4060 43596 4116
rect 43652 4060 48000 4116
rect 0 4032 800 4060
rect 47200 4032 48000 4060
rect 37874 3948 37884 4004
rect 37940 3948 39788 4004
rect 39844 3948 39854 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 7186 3724 7196 3780
rect 7252 3724 11900 3780
rect 11956 3724 11966 3780
rect 33506 3724 33516 3780
rect 33572 3724 36540 3780
rect 36596 3724 36606 3780
rect 10994 3612 11004 3668
rect 11060 3612 23548 3668
rect 23604 3612 23614 3668
rect 29586 3612 29596 3668
rect 29652 3612 30492 3668
rect 30548 3612 30558 3668
rect 36306 3612 36316 3668
rect 36372 3612 36988 3668
rect 37044 3612 37054 3668
rect 38994 3612 39004 3668
rect 39060 3612 40236 3668
rect 40292 3612 40302 3668
rect 42690 3612 42700 3668
rect 42756 3612 46060 3668
rect 46116 3612 46126 3668
rect 8754 3500 8764 3556
rect 8820 3500 12068 3556
rect 12226 3500 12236 3556
rect 12292 3500 13468 3556
rect 13524 3500 13534 3556
rect 15092 3500 23324 3556
rect 23380 3500 23390 3556
rect 24434 3500 24444 3556
rect 24500 3500 25116 3556
rect 25172 3500 25182 3556
rect 25666 3500 25676 3556
rect 25732 3500 26460 3556
rect 26516 3500 26908 3556
rect 26964 3500 26974 3556
rect 27122 3500 27132 3556
rect 27188 3500 27692 3556
rect 27748 3500 27758 3556
rect 33618 3500 33628 3556
rect 33684 3500 34972 3556
rect 35028 3500 35038 3556
rect 0 3444 800 3472
rect 12012 3444 12068 3500
rect 15092 3444 15148 3500
rect 47200 3444 48000 3472
rect 0 3388 1708 3444
rect 1764 3388 2940 3444
rect 2996 3388 3006 3444
rect 12012 3388 15148 3444
rect 21186 3388 21196 3444
rect 21252 3388 22092 3444
rect 22148 3388 22158 3444
rect 26226 3388 26236 3444
rect 26292 3388 27244 3444
rect 27300 3388 27310 3444
rect 28242 3388 28252 3444
rect 28308 3388 29260 3444
rect 29316 3388 29326 3444
rect 32946 3388 32956 3444
rect 33012 3388 33852 3444
rect 33908 3388 34300 3444
rect 34356 3388 34366 3444
rect 38546 3388 38556 3444
rect 38612 3388 39116 3444
rect 39172 3388 39182 3444
rect 43026 3388 43036 3444
rect 43092 3388 48000 3444
rect 0 3360 800 3388
rect 47200 3360 48000 3388
rect 34962 3276 34972 3332
rect 35028 3276 35980 3332
rect 36036 3276 36046 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 2772 800 2800
rect 47200 2772 48000 2800
rect 0 2716 2380 2772
rect 2436 2716 2446 2772
rect 45266 2716 45276 2772
rect 45332 2716 48000 2772
rect 0 2688 800 2716
rect 47200 2688 48000 2716
rect 47200 2100 48000 2128
rect 44370 2044 44380 2100
rect 44436 2044 48000 2100
rect 47200 2016 48000 2044
rect 47200 1428 48000 1456
rect 43586 1372 43596 1428
rect 43652 1372 48000 1428
rect 47200 1344 48000 1372
rect 47200 756 48000 784
rect 44818 700 44828 756
rect 44884 700 48000 756
rect 47200 672 48000 700
rect 47200 84 48000 112
rect 45266 28 45276 84
rect 45332 28 48000 84
rect 47200 0 48000 28
<< via3 >>
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 44716 21756 44772 21812
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 41244 20748 41300 20804
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 36652 16940 36708 16996
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 41244 15148 41300 15204
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 36652 9996 36708 10052
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 44716 8876 44772 8932
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 44716 4768 44748
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 43932 20128 44748
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 44716 35488 44748
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 44716 21812 44772 21822
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 41244 20804 41300 20814
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 36652 16996 36708 17006
rect 36652 10052 36708 16940
rect 41244 15204 41300 20748
rect 41244 15138 41300 15148
rect 36652 9986 36708 9996
rect 44716 8932 44772 21756
rect 44716 8866 44772 8876
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32368 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 1 26656
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _180_
timestamp 1698431365
transform 1 0 6048 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14000 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _182_
timestamp 1698431365
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _183_
timestamp 1698431365
transform -1 0 14112 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _184_
timestamp 1698431365
transform -1 0 10080 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _185_
timestamp 1698431365
transform -1 0 14672 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _186_
timestamp 1698431365
transform 1 0 5712 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _187_
timestamp 1698431365
transform -1 0 2240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _188_
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _189_
timestamp 1698431365
transform -1 0 12768 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _190_
timestamp 1698431365
transform -1 0 10192 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _191_
timestamp 1698431365
transform -1 0 9072 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _192_
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _193_
timestamp 1698431365
transform 1 0 1792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _194_
timestamp 1698431365
transform 1 0 1792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _195_
timestamp 1698431365
transform -1 0 2352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _196_
timestamp 1698431365
transform 1 0 1792 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _197_
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _198_
timestamp 1698431365
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _199_
timestamp 1698431365
transform 1 0 3248 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _200_
timestamp 1698431365
transform 1 0 1792 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _201_
timestamp 1698431365
transform 1 0 1792 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _202_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _203_
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _204_
timestamp 1698431365
transform -1 0 16912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _205_
timestamp 1698431365
transform 1 0 11424 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _206_
timestamp 1698431365
transform -1 0 11424 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _207_
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _208_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _209_
timestamp 1698431365
transform -1 0 13104 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _210_
timestamp 1698431365
transform -1 0 14000 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _211_
timestamp 1698431365
transform -1 0 14672 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _212_
timestamp 1698431365
transform -1 0 11760 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _213_
timestamp 1698431365
transform -1 0 8736 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _214_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _215_
timestamp 1698431365
transform -1 0 7280 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _216_
timestamp 1698431365
transform -1 0 8960 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _217_
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _218_
timestamp 1698431365
transform -1 0 6832 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _219_
timestamp 1698431365
transform -1 0 6160 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _220_
timestamp 1698431365
transform 1 0 1792 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _221_
timestamp 1698431365
transform 1 0 1792 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _222_
timestamp 1698431365
transform -1 0 6160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _223_
timestamp 1698431365
transform -1 0 3472 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _224_
timestamp 1698431365
transform -1 0 12768 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _225_
timestamp 1698431365
transform -1 0 17024 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _226_
timestamp 1698431365
transform -1 0 17920 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _227_
timestamp 1698431365
transform -1 0 17920 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _228_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _229_
timestamp 1698431365
transform -1 0 14784 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _230_
timestamp 1698431365
transform 1 0 11312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _231_
timestamp 1698431365
transform -1 0 11312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _232_
timestamp 1698431365
transform -1 0 12544 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _233_
timestamp 1698431365
transform -1 0 15456 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _234_
timestamp 1698431365
transform -1 0 14000 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _235_
timestamp 1698431365
transform -1 0 24080 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _236_
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _237_
timestamp 1698431365
transform -1 0 25760 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _238_
timestamp 1698431365
transform -1 0 25760 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _239_
timestamp 1698431365
transform -1 0 23520 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _240_
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _241_
timestamp 1698431365
transform -1 0 21840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _242_
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _243_
timestamp 1698431365
transform -1 0 24752 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _244_
timestamp 1698431365
transform 1 0 21280 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _245_
timestamp 1698431365
transform -1 0 20720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _246_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _247_
timestamp 1698431365
transform -1 0 19376 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _248_
timestamp 1698431365
transform 1 0 17808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _249_
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _250_
timestamp 1698431365
transform -1 0 19600 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _251_
timestamp 1698431365
transform 1 0 18480 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _252_
timestamp 1698431365
transform -1 0 18256 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _253_
timestamp 1698431365
transform -1 0 19152 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _254_
timestamp 1698431365
transform -1 0 18368 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _255_
timestamp 1698431365
transform -1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _256_
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _257_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _258_
timestamp 1698431365
transform -1 0 25760 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _259_
timestamp 1698431365
transform -1 0 24528 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _260_
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _261_
timestamp 1698431365
transform 1 0 27888 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _262_
timestamp 1698431365
transform -1 0 27216 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _263_
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _264_
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _265_
timestamp 1698431365
transform -1 0 22736 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _266_
timestamp 1698431365
transform -1 0 23856 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _267_
timestamp 1698431365
transform -1 0 22064 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _268_
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _269_
timestamp 1698431365
transform 1 0 35728 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _270_
timestamp 1698431365
transform 1 0 35728 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _271_
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _272_
timestamp 1698431365
transform 1 0 34720 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _273_
timestamp 1698431365
transform -1 0 34272 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _274_
timestamp 1698431365
transform -1 0 33600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _275_
timestamp 1698431365
transform -1 0 30464 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _276_
timestamp 1698431365
transform -1 0 32704 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _277_
timestamp 1698431365
transform 1 0 34384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _278_
timestamp 1698431365
transform -1 0 35616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _279_
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _280_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _281_
timestamp 1698431365
transform -1 0 45584 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _282_
timestamp 1698431365
transform 1 0 45472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _283_
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _284_
timestamp 1698431365
transform 1 0 39648 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _285_
timestamp 1698431365
transform 1 0 38080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _286_
timestamp 1698431365
transform -1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _287_
timestamp 1698431365
transform -1 0 45472 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _288_
timestamp 1698431365
transform 1 0 42784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _289_
timestamp 1698431365
transform 1 0 39648 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _290_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35056 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _291_
timestamp 1698431365
transform 1 0 42112 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _292_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _293_
timestamp 1698431365
transform -1 0 39424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _294_
timestamp 1698431365
transform -1 0 36288 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _295_
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _296_
timestamp 1698431365
transform -1 0 36064 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _297_
timestamp 1698431365
transform -1 0 37520 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _298_
timestamp 1698431365
transform -1 0 40208 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _299_
timestamp 1698431365
transform -1 0 36288 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _300_
timestamp 1698431365
transform -1 0 41440 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _301_
timestamp 1698431365
transform 1 0 38864 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _302_
timestamp 1698431365
transform 1 0 45360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _303_
timestamp 1698431365
transform 1 0 45360 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _304_
timestamp 1698431365
transform 1 0 45360 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _305_
timestamp 1698431365
transform 1 0 43568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _306_
timestamp 1698431365
transform 1 0 45360 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _307_
timestamp 1698431365
transform -1 0 45360 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _308_
timestamp 1698431365
transform -1 0 45248 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _309_
timestamp 1698431365
transform -1 0 45360 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _310_
timestamp 1698431365
transform -1 0 43344 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _311_
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _312_
timestamp 1698431365
transform -1 0 32256 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _313_
timestamp 1698431365
transform 1 0 33040 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _314_
timestamp 1698431365
transform 1 0 35616 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _315_
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _316_
timestamp 1698431365
transform -1 0 33600 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _317_
timestamp 1698431365
transform -1 0 31696 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _318_
timestamp 1698431365
transform 1 0 30688 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _319_
timestamp 1698431365
transform -1 0 31024 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _320_
timestamp 1698431365
transform 1 0 28112 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _321_
timestamp 1698431365
transform -1 0 32256 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _322_
timestamp 1698431365
transform -1 0 27776 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _323_
timestamp 1698431365
transform -1 0 30576 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _324_
timestamp 1698431365
transform -1 0 26208 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _325_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _326_
timestamp 1698431365
transform 1 0 23632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _327_
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _328_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _329_
timestamp 1698431365
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _330_
timestamp 1698431365
transform -1 0 24080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _331_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _332_
timestamp 1698431365
transform -1 0 21952 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _333_
timestamp 1698431365
transform -1 0 19600 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _334_
timestamp 1698431365
transform -1 0 32256 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _335_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _336_
timestamp 1698431365
transform -1 0 31360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _337_
timestamp 1698431365
transform -1 0 33600 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _338_
timestamp 1698431365
transform -1 0 26880 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _339_
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _340_
timestamp 1698431365
transform -1 0 34944 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _341_
timestamp 1698431365
transform -1 0 34272 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _342_
timestamp 1698431365
transform -1 0 32256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _343_
timestamp 1698431365
transform -1 0 33600 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _344_
timestamp 1698431365
transform -1 0 31584 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _345_
timestamp 1698431365
transform 1 0 37968 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _346_
timestamp 1698431365
transform -1 0 44352 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _347_
timestamp 1698431365
transform -1 0 45360 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _348_
timestamp 1698431365
transform -1 0 45920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _349_
timestamp 1698431365
transform -1 0 45248 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _350_
timestamp 1698431365
transform -1 0 45360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _351_
timestamp 1698431365
transform 1 0 43456 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _352_
timestamp 1698431365
transform -1 0 43456 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _353_
timestamp 1698431365
transform -1 0 44464 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _354_
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _355_
timestamp 1698431365
transform -1 0 41440 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _356_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13216 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _357_
timestamp 1698431365
transform 1 0 8960 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _358_
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _359_
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _360_
timestamp 1698431365
transform 1 0 5040 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _361_
timestamp 1698431365
transform -1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _362_
timestamp 1698431365
transform -1 0 13216 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _363_
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _364_
timestamp 1698431365
transform 1 0 8288 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _365_
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _366_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _367_
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _368_
timestamp 1698431365
transform -1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _369_
timestamp 1698431365
transform -1 0 13216 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _370_
timestamp 1698431365
transform 1 0 1904 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _371_
timestamp 1698431365
transform -1 0 5376 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _372_
timestamp 1698431365
transform 1 0 2352 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _373_
timestamp 1698431365
transform -1 0 5488 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _374_
timestamp 1698431365
transform -1 0 5712 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _375_
timestamp 1698431365
transform -1 0 5376 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _376_
timestamp 1698431365
transform -1 0 16912 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _377_
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _378_
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _379_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _380_
timestamp 1698431365
transform 1 0 13216 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _381_
timestamp 1698431365
transform 1 0 11760 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _382_
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _383_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _384_
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _385_
timestamp 1698431365
transform 1 0 7952 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _386_
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _387_
timestamp 1698431365
transform -1 0 7728 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _388_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _389_
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _390_
timestamp 1698431365
transform -1 0 7280 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _391_
timestamp 1698431365
transform 1 0 2352 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _392_
timestamp 1698431365
transform -1 0 9296 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _393_
timestamp 1698431365
transform -1 0 5488 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _394_
timestamp 1698431365
transform 1 0 2016 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _395_
timestamp 1698431365
transform -1 0 5376 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _396_
timestamp 1698431365
transform -1 0 19376 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _397_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _398_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _399_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _400_
timestamp 1698431365
transform 1 0 9296 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _401_
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _402_
timestamp 1698431365
transform -1 0 13216 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _403_
timestamp 1698431365
transform 1 0 8064 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _404_
timestamp 1698431365
transform 1 0 11984 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _405_
timestamp 1698431365
transform 1 0 9296 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _406_
timestamp 1698431365
transform -1 0 25760 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _407_
timestamp 1698431365
transform 1 0 21056 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _408_
timestamp 1698431365
transform 1 0 20608 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _409_
timestamp 1698431365
transform -1 0 24976 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _410_
timestamp 1698431365
transform 1 0 17136 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _411_
timestamp 1698431365
transform -1 0 21056 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _412_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _413_
timestamp 1698431365
transform -1 0 24528 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _414_
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _415_
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _416_
timestamp 1698431365
transform -1 0 20048 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _417_
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _418_
timestamp 1698431365
transform 1 0 13216 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _419_
timestamp 1698431365
transform 1 0 13216 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _420_
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _421_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _422_
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _423_
timestamp 1698431365
transform 1 0 13216 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _424_
timestamp 1698431365
transform -1 0 18928 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _425_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _426_
timestamp 1698431365
transform -1 0 26096 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _427_
timestamp 1698431365
transform 1 0 21056 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _428_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _429_
timestamp 1698431365
transform -1 0 28896 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _430_
timestamp 1698431365
transform 1 0 23744 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _431_
timestamp 1698431365
transform 1 0 22736 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _432_
timestamp 1698431365
transform 1 0 21056 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _433_
timestamp 1698431365
transform -1 0 24976 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _434_
timestamp 1698431365
transform 1 0 20160 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _435_
timestamp 1698431365
transform 1 0 19152 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _436_
timestamp 1698431365
transform -1 0 40656 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _437_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _438_
timestamp 1698431365
transform -1 0 36736 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _439_
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _440_
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _441_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _442_
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _443_
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _444_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _445_
timestamp 1698431365
transform 1 0 30464 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _446_
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _447_
timestamp 1698431365
transform 1 0 40656 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _448_
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _449_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _450_
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _451_
timestamp 1698431365
transform 1 0 36736 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _452_
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _453_
timestamp 1698431365
transform 1 0 40656 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _454_
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _455_
timestamp 1698431365
transform 1 0 37856 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _456_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _457_
timestamp 1698431365
transform 1 0 34160 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _458_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _459_
timestamp 1698431365
transform 1 0 32816 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _460_
timestamp 1698431365
transform 1 0 35056 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _461_
timestamp 1698431365
transform 1 0 33600 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _462_
timestamp 1698431365
transform -1 0 36736 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _463_
timestamp 1698431365
transform -1 0 40544 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _464_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _465_
timestamp 1698431365
transform 1 0 31584 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _466_
timestamp 1698431365
transform 1 0 42000 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _467_
timestamp 1698431365
transform 1 0 41440 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _468_
timestamp 1698431365
transform -1 0 45584 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _469_
timestamp 1698431365
transform 1 0 40880 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _470_
timestamp 1698431365
transform 1 0 40656 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _471_
timestamp 1698431365
transform 1 0 41440 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _472_
timestamp 1698431365
transform 1 0 41776 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _473_
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _474_
timestamp 1698431365
transform 1 0 38864 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _475_
timestamp 1698431365
transform 1 0 37184 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _476_
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _477_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _478_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _479_
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _480_
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _481_
timestamp 1698431365
transform -1 0 32816 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _482_
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _483_
timestamp 1698431365
transform 1 0 25984 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _484_
timestamp 1698431365
transform -1 0 32816 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _485_
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _486_
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _487_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _488_
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _489_
timestamp 1698431365
transform 1 0 19600 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _490_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _491_
timestamp 1698431365
transform -1 0 20048 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _492_
timestamp 1698431365
transform -1 0 24192 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _493_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _494_
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _495_
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _496_
timestamp 1698431365
transform -1 0 32816 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _497_
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _498_
timestamp 1698431365
transform 1 0 25648 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _499_
timestamp 1698431365
transform 1 0 24304 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _500_
timestamp 1698431365
transform 1 0 29120 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _501_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _502_
timestamp 1698431365
transform 1 0 24976 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _503_
timestamp 1698431365
transform -1 0 29904 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _504_
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _505_
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _506_
timestamp 1698431365
transform 1 0 36736 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _507_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _508_
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _509_
timestamp 1698431365
transform 1 0 41328 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _510_
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _511_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _512_
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _513_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _514_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _515_
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _536_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _537_
timestamp 1698431365
transform 1 0 31696 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _538_
timestamp 1698431365
transform 1 0 37408 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _539_
timestamp 1698431365
transform 1 0 38864 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _540_
timestamp 1698431365
transform 1 0 43792 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _541_
timestamp 1698431365
transform -1 0 24192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _542_
timestamp 1698431365
transform -1 0 19376 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _543_
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _544_
timestamp 1698431365
transform -1 0 26768 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _545_
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _546_
timestamp 1698431365
transform 1 0 33040 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _547_
timestamp 1698431365
transform -1 0 22736 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _548_
timestamp 1698431365
transform 1 0 29120 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _549_
timestamp 1698431365
transform 1 0 25872 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _550_
timestamp 1698431365
transform -1 0 45360 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _551_
timestamp 1698431365
transform -1 0 22960 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _552_
timestamp 1698431365
transform 1 0 13664 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _553_
timestamp 1698431365
transform 1 0 25424 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _554_
timestamp 1698431365
transform -1 0 23520 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _555_
timestamp 1698431365
transform 1 0 14560 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _556_
timestamp 1698431365
transform 1 0 12096 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _557_
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _558_
timestamp 1698431365
transform 1 0 23072 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _559_
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _560_
timestamp 1698431365
transform -1 0 28672 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _561_
timestamp 1698431365
transform -1 0 23856 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _562_
timestamp 1698431365
transform 1 0 26656 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _563_
timestamp 1698431365
transform 1 0 15456 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _564_
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _565_
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _566_
timestamp 1698431365
transform -1 0 20944 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _567_
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _568_
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _569_
timestamp 1698431365
transform -1 0 18928 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _570_
timestamp 1698431365
transform 1 0 31024 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _571_
timestamp 1698431365
transform 1 0 27328 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _572_
timestamp 1698431365
transform 1 0 38752 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _573_
timestamp 1698431365
transform -1 0 14000 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _574_
timestamp 1698431365
transform 1 0 40096 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _575_
timestamp 1698431365
transform -1 0 21280 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _576_
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _577_
timestamp 1698431365
transform 1 0 23632 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _578_
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _579_
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _580_
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _581_
timestamp 1698431365
transform 1 0 45696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _582_
timestamp 1698431365
transform 1 0 43792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _583_
timestamp 1698431365
transform 1 0 39872 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _584_
timestamp 1698431365
transform 1 0 36960 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _585_
timestamp 1698431365
transform 1 0 33712 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _586_
timestamp 1698431365
transform -1 0 22736 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _587_
timestamp 1698431365
transform -1 0 17136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _588_
timestamp 1698431365
transform 1 0 38080 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _589_
timestamp 1698431365
transform 1 0 26544 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _590_
timestamp 1698431365
transform 1 0 39424 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _591_
timestamp 1698431365
transform 1 0 44240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _592_
timestamp 1698431365
transform 1 0 29792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _593_
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _594_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _595_
timestamp 1698431365
transform 1 0 38080 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1698431365
transform 1 0 8400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I
timestamp 1698431365
transform 1 0 2688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1698431365
transform 1 0 3136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1698431365
transform 1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I
timestamp 1698431365
transform -1 0 10640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1698431365
transform 1 0 8848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__I
timestamp 1698431365
transform 1 0 8960 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__I
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I
timestamp 1698431365
transform 1 0 17920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__I
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__I
timestamp 1698431365
transform 1 0 12320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I
timestamp 1698431365
transform 1 0 11312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__I
timestamp 1698431365
transform -1 0 9968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I
timestamp 1698431365
transform 1 0 10416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__I
timestamp 1698431365
transform 1 0 24976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__I
timestamp 1698431365
transform 1 0 20832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I
timestamp 1698431365
transform 1 0 33600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I
timestamp 1698431365
transform 1 0 43792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__I
timestamp 1698431365
transform 1 0 46032 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__I
timestamp 1698431365
transform 1 0 46144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__I
timestamp 1698431365
transform 1 0 46144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I
timestamp 1698431365
transform 1 0 42448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__I
timestamp 1698431365
transform 1 0 45584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1698431365
transform -1 0 38864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__I
timestamp 1698431365
transform 1 0 41664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__CLK
timestamp 1698431365
transform 1 0 5824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__CLK
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__CLK
timestamp 1698431365
transform 1 0 6272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__CLK
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__CLK
timestamp 1698431365
transform 1 0 9968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__CLK
timestamp 1698431365
transform -1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__CLK
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__CLK
timestamp 1698431365
transform 1 0 8064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__CLK
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__CLK
timestamp 1698431365
transform 1 0 7168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__CLK
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__CLK
timestamp 1698431365
transform 1 0 6160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__CLK
timestamp 1698431365
transform -1 0 5936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__CLK
timestamp 1698431365
transform 1 0 6048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__D
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__CLK
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__CLK
timestamp 1698431365
transform 1 0 13552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__CLK
timestamp 1698431365
transform -1 0 12432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__CLK
timestamp 1698431365
transform -1 0 12208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__CLK
timestamp 1698431365
transform 1 0 14896 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__CLK
timestamp 1698431365
transform 1 0 9968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__CLK
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__CLK
timestamp 1698431365
transform 1 0 14336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__CLK
timestamp 1698431365
transform 1 0 41216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__CLK
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__CLK
timestamp 1698431365
transform -1 0 41776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__CLK
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__CLK
timestamp 1698431365
transform 1 0 41216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__CLK
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__CLK
timestamp 1698431365
transform 1 0 40432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__CLK
timestamp 1698431365
transform 1 0 36960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__CLK
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__D
timestamp 1698431365
transform 1 0 30016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__CLK
timestamp 1698431365
transform 1 0 44912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__CLK
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__I
timestamp 1698431365
transform -1 0 28896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__I
timestamp 1698431365
transform -1 0 35504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__I
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__I
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__I
timestamp 1698431365
transform 1 0 33824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform -1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_prog_clk_I
timestamp 1698431365
transform 1 0 7616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_prog_clk_I
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_prog_clk_I
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_prog_clk_I
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_prog_clk_I
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_prog_clk_I
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_prog_clk_I
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_prog_clk_I
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_prog_clk_I
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_prog_clk_I
timestamp 1698431365
transform 1 0 27776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_prog_clk_I
timestamp 1698431365
transform 1 0 36960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_prog_clk_I
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_prog_clk_I
timestamp 1698431365
transform 1 0 29232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_prog_clk_I
timestamp 1698431365
transform -1 0 27104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_prog_clk_I
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_prog_clk_I
timestamp 1698431365
transform 1 0 37072 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 41776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 13552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 25088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 13552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 11984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 14224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 11424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 33376 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 29904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 23856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 46368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 19824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 24640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 45696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 39760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 37968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 31696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 23184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 26544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 31024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 20496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 33936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 9520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 25424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 34384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 18032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 22288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 35056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 40992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 46368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 44800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 35728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 34832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 30352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 46144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 42672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 26320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 7504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 31696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 44016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 43232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform -1 0 42784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform -1 0 18256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 20944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 45584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 44688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 37968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform -1 0 39760 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform -1 0 45696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output99_I
timestamp 1698431365
transform 1 0 43792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1698431365
transform 1 0 46144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output105_I
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1698431365
transform -1 0 3584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output123_I
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1698431365
transform -1 0 9184 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1698431365
transform -1 0 24080 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1698431365
transform 1 0 9968 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1698431365
transform 1 0 17808 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1698431365
transform -1 0 20496 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1698431365
transform -1 0 32032 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1698431365
transform -1 0 30912 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1698431365
transform -1 0 39984 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1698431365
transform -1 0 40096 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1698431365
transform 1 0 28896 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1698431365
transform -1 0 40208 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_16 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32
timestamp 1698431365
transform 1 0 4928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_44 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_54
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_114
timestamp 1698431365
transform 1 0 14112 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_122
timestamp 1698431365
transform 1 0 15008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_156
timestamp 1698431365
transform 1 0 18816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_191
timestamp 1698431365
transform 1 0 22736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_221
timestamp 1698431365
transform 1 0 26096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_251
timestamp 1698431365
transform 1 0 29456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_265
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_276
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_287
timestamp 1698431365
transform 1 0 33488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_312
timestamp 1698431365
transform 1 0 36288 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_323
timestamp 1698431365
transform 1 0 37520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_352
timestamp 1698431365
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_366
timestamp 1698431365
transform 1 0 42336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_394
timestamp 1698431365
transform 1 0 45472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_44
timestamp 1698431365
transform 1 0 6272 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_52
timestamp 1698431365
transform 1 0 7168 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_56
timestamp 1698431365
transform 1 0 7616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_83
timestamp 1698431365
transform 1 0 10640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_87
timestamp 1698431365
transform 1 0 11088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_89
timestamp 1698431365
transform 1 0 11312 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_92
timestamp 1698431365
transform 1 0 11648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_94
timestamp 1698431365
transform 1 0 11872 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_107
timestamp 1698431365
transform 1 0 13328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_111
timestamp 1698431365
transform 1 0 13776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_131
timestamp 1698431365
transform 1 0 16016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_135
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_137
timestamp 1698431365
transform 1 0 16688 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_155
timestamp 1698431365
transform 1 0 18704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_169
timestamp 1698431365
transform 1 0 20272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_173
timestamp 1698431365
transform 1 0 20720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_185
timestamp 1698431365
transform 1 0 22064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_201
timestamp 1698431365
transform 1 0 23856 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_233
timestamp 1698431365
transform 1 0 27440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_243
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_251
timestamp 1698431365
transform 1 0 29456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_255
timestamp 1698431365
transform 1 0 29904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_294
timestamp 1698431365
transform 1 0 34272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_301
timestamp 1698431365
transform 1 0 35056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_305
timestamp 1698431365
transform 1 0 35504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_313
timestamp 1698431365
transform 1 0 36400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_317
timestamp 1698431365
transform 1 0 36848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_329
timestamp 1698431365
transform 1 0 38192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_333
timestamp 1698431365
transform 1 0 38640 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_358
timestamp 1698431365
transform 1 0 41440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_360
timestamp 1698431365
transform 1 0 41664 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_367
timestamp 1698431365
transform 1 0 42448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_389
timestamp 1698431365
transform 1 0 44912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_69
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_73
timestamp 1698431365
transform 1 0 9520 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_89
timestamp 1698431365
transform 1 0 11312 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_93
timestamp 1698431365
transform 1 0 11760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_95
timestamp 1698431365
transform 1 0 11984 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_113
timestamp 1698431365
transform 1 0 14000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_117
timestamp 1698431365
transform 1 0 14448 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_124
timestamp 1698431365
transform 1 0 15232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_132
timestamp 1698431365
transform 1 0 16128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_134
timestamp 1698431365
transform 1 0 16352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_147
timestamp 1698431365
transform 1 0 17808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_157
timestamp 1698431365
transform 1 0 18928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_215
timestamp 1698431365
transform 1 0 25424 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_231
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_235
timestamp 1698431365
transform 1 0 27664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_237
timestamp 1698431365
transform 1 0 27888 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_260
timestamp 1698431365
transform 1 0 30464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_262
timestamp 1698431365
transform 1 0 30688 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_295
timestamp 1698431365
transform 1 0 34384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_299
timestamp 1698431365
transform 1 0 34832 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_303
timestamp 1698431365
transform 1 0 35280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_307
timestamp 1698431365
transform 1 0 35728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_334
timestamp 1698431365
transform 1 0 38752 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_341
timestamp 1698431365
transform 1 0 39536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_343
timestamp 1698431365
transform 1 0 39760 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_350
timestamp 1698431365
transform 1 0 40544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_354
timestamp 1698431365
transform 1 0 40992 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_358
timestamp 1698431365
transform 1 0 41440 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_361
timestamp 1698431365
transform 1 0 41776 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_369
timestamp 1698431365
transform 1 0 42672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_373
timestamp 1698431365
transform 1 0 43120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_398
timestamp 1698431365
transform 1 0 45920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_16
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_48
timestamp 1698431365
transform 1 0 6720 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_64
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_158
timestamp 1698431365
transform 1 0 19040 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_166
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_178
timestamp 1698431365
transform 1 0 21280 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_182
timestamp 1698431365
transform 1 0 21728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_184
timestamp 1698431365
transform 1 0 21952 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_191
timestamp 1698431365
transform 1 0 22736 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_204
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_242
timestamp 1698431365
transform 1 0 28448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_246
timestamp 1698431365
transform 1 0 28896 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_288
timestamp 1698431365
transform 1 0 33600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_292
timestamp 1698431365
transform 1 0 34048 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_324
timestamp 1698431365
transform 1 0 37632 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_340
timestamp 1698431365
transform 1 0 39424 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_384
timestamp 1698431365
transform 1 0 44352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_16
timestamp 1698431365
transform 1 0 3136 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_349
timestamp 1698431365
transform 1 0 40432 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_357
timestamp 1698431365
transform 1 0 41328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_359
timestamp 1698431365
transform 1 0 41552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_376
timestamp 1698431365
transform 1 0 43456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_398
timestamp 1698431365
transform 1 0 45920 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_16
timestamp 1698431365
transform 1 0 3136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_20
timestamp 1698431365
transform 1 0 3584 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_52
timestamp 1698431365
transform 1 0 7168 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_354
timestamp 1698431365
transform 1 0 40992 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_371
timestamp 1698431365
transform 1 0 42896 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_379
timestamp 1698431365
transform 1 0 43792 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_383
timestamp 1698431365
transform 1 0 44240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_387
timestamp 1698431365
transform 1 0 44688 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_16
timestamp 1698431365
transform 1 0 3136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_20
timestamp 1698431365
transform 1 0 3584 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_333
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_341
timestamp 1698431365
transform 1 0 39536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_345
timestamp 1698431365
transform 1 0 39984 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_362
timestamp 1698431365
transform 1 0 41888 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_378
timestamp 1698431365
transform 1 0 43680 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_398
timestamp 1698431365
transform 1 0 45920 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_294
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_312
timestamp 1698431365
transform 1 0 36288 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_344
timestamp 1698431365
transform 1 0 39872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_368
timestamp 1698431365
transform 1 0 42560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_376
timestamp 1698431365
transform 1 0 43456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_378
timestamp 1698431365
transform 1 0 43680 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_381
timestamp 1698431365
transform 1 0 44016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_385
timestamp 1698431365
transform 1 0 44464 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_57
timestamp 1698431365
transform 1 0 7728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_65
timestamp 1698431365
transform 1 0 8624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_67
timestamp 1698431365
transform 1 0 8848 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_84
timestamp 1698431365
transform 1 0 10752 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_100
timestamp 1698431365
transform 1 0 12544 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_295
timestamp 1698431365
transform 1 0 34384 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_345
timestamp 1698431365
transform 1 0 39984 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_353
timestamp 1698431365
transform 1 0 40880 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_370
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_372
timestamp 1698431365
transform 1 0 43008 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_398
timestamp 1698431365
transform 1 0 45920 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_36
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_54
timestamp 1698431365
transform 1 0 7392 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_97
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_129
timestamp 1698431365
transform 1 0 15792 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_240
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_272
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_310
timestamp 1698431365
transform 1 0 36064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_318
timestamp 1698431365
transform 1 0 36960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_320
timestamp 1698431365
transform 1 0 37184 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_337
timestamp 1698431365
transform 1 0 39088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_345
timestamp 1698431365
transform 1 0 39984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_368
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_386
timestamp 1698431365
transform 1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_390
timestamp 1698431365
transform 1 0 45024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_392
timestamp 1698431365
transform 1 0 45248 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_401
timestamp 1698431365
transform 1 0 46256 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_6
timestamp 1698431365
transform 1 0 2016 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_23
timestamp 1698431365
transform 1 0 3920 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_43
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_60
timestamp 1698431365
transform 1 0 8064 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_68
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_85
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_194
timestamp 1698431365
transform 1 0 23072 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_210
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_228
timestamp 1698431365
transform 1 0 26880 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_264
timestamp 1698431365
transform 1 0 30912 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_280
timestamp 1698431365
transform 1 0 32704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_284
timestamp 1698431365
transform 1 0 33152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_342
timestamp 1698431365
transform 1 0 39648 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_358
timestamp 1698431365
transform 1 0 41440 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_362
timestamp 1698431365
transform 1 0 41888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_380
timestamp 1698431365
transform 1 0 43904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_398
timestamp 1698431365
transform 1 0 45920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_36
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_48
timestamp 1698431365
transform 1 0 6720 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_65
timestamp 1698431365
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_92
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_110
timestamp 1698431365
transform 1 0 13664 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_126
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_134
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_240
timestamp 1698431365
transform 1 0 28224 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_248
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_265
timestamp 1698431365
transform 1 0 31024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_298
timestamp 1698431365
transform 1 0 34720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_316
timestamp 1698431365
transform 1 0 36736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_318
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_335
timestamp 1698431365
transform 1 0 38864 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_343
timestamp 1698431365
transform 1 0 39760 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_377
timestamp 1698431365
transform 1 0 43568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_385
timestamp 1698431365
transform 1 0 44464 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_6
timestamp 1698431365
transform 1 0 2016 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_23
timestamp 1698431365
transform 1 0 3920 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_31
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_43
timestamp 1698431365
transform 1 0 6160 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_60
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_76
timestamp 1698431365
transform 1 0 9856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_141
timestamp 1698431365
transform 1 0 17136 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_203
timestamp 1698431365
transform 1 0 24080 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_219
timestamp 1698431365
transform 1 0 25872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_237
timestamp 1698431365
transform 1 0 27888 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_273
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_281
timestamp 1698431365
transform 1 0 32816 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_304
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_306
timestamp 1698431365
transform 1 0 35616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_343
timestamp 1698431365
transform 1 0 39760 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_351
timestamp 1698431365
transform 1 0 40656 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_368
timestamp 1698431365
transform 1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_370
timestamp 1698431365
transform 1 0 42784 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_398
timestamp 1698431365
transform 1 0 45920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_4
timestamp 1698431365
transform 1 0 1792 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_61
timestamp 1698431365
transform 1 0 8176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_65
timestamp 1698431365
transform 1 0 8624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_98
timestamp 1698431365
transform 1 0 12320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_115
timestamp 1698431365
transform 1 0 14224 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_123
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_192
timestamp 1698431365
transform 1 0 22848 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_200
timestamp 1698431365
transform 1 0 23744 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_248
timestamp 1698431365
transform 1 0 29120 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_265
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_301
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_309
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_326
timestamp 1698431365
transform 1 0 37856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_336
timestamp 1698431365
transform 1 0 38976 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_344
timestamp 1698431365
transform 1 0 39872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_360
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_364
timestamp 1698431365
transform 1 0 42112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_372
timestamp 1698431365
transform 1 0 43008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_376
timestamp 1698431365
transform 1 0 43456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_378
timestamp 1698431365
transform 1 0 43680 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_397
timestamp 1698431365
transform 1 0 45808 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_401
timestamp 1698431365
transform 1 0 46256 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_14
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_71
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_75
timestamp 1698431365
transform 1 0 9744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_79
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_96
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_135
timestamp 1698431365
transform 1 0 16464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_199
timestamp 1698431365
transform 1 0 23632 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_287
timestamp 1698431365
transform 1 0 33488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_295
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_350
timestamp 1698431365
transform 1 0 40544 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_366
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_24
timestamp 1698431365
transform 1 0 4032 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_32
timestamp 1698431365
transform 1 0 4928 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_78
timestamp 1698431365
transform 1 0 10080 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_82
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_86
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_106
timestamp 1698431365
transform 1 0 13216 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_114
timestamp 1698431365
transform 1 0 14112 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_131
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_166
timestamp 1698431365
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_202
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_243
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_316
timestamp 1698431365
transform 1 0 36736 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_324
timestamp 1698431365
transform 1 0 37632 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_328
timestamp 1698431365
transform 1 0 38080 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_43
timestamp 1698431365
transform 1 0 6160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_96
timestamp 1698431365
transform 1 0 12096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_100
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_159
timestamp 1698431365
transform 1 0 19152 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_106
timestamp 1698431365
transform 1 0 13216 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_113
timestamp 1698431365
transform 1 0 14000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_131
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_167
timestamp 1698431365
transform 1 0 20048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_175
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_386
timestamp 1698431365
transform 1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_39
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_114
timestamp 1698431365
transform 1 0 14112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_118
timestamp 1698431365
transform 1 0 14560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_122
timestamp 1698431365
transform 1 0 15008 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_231
timestamp 1698431365
transform 1 0 27216 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_253
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_353
timestamp 1698431365
transform 1 0 40880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_361
timestamp 1698431365
transform 1 0 41776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_363
timestamp 1698431365
transform 1 0 42000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_380
timestamp 1698431365
transform 1 0 43904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_382
timestamp 1698431365
transform 1 0 44128 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_152
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_193
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_316
timestamp 1698431365
transform 1 0 36736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_386
timestamp 1698431365
transform 1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_55
timestamp 1698431365
transform 1 0 7504 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_58
timestamp 1698431365
transform 1 0 7840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_119
timestamp 1698431365
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_169
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_184
timestamp 1698431365
transform 1 0 21952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_186
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_221
timestamp 1698431365
transform 1 0 26096 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_229
timestamp 1698431365
transform 1 0 26992 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_233
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_235
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_345
timestamp 1698431365
transform 1 0 39984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_4
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_43
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_168
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_172
timestamp 1698431365
transform 1 0 20608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_255
timestamp 1698431365
transform 1 0 29904 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_263
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_294
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_340
timestamp 1698431365
transform 1 0 39424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_360
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_377
timestamp 1698431365
transform 1 0 43568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_381
timestamp 1698431365
transform 1 0 44016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_383
timestamp 1698431365
transform 1 0 44240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_203
timestamp 1698431365
transform 1 0 24080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_205
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_281
timestamp 1698431365
transform 1 0 32816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_285
timestamp 1698431365
transform 1 0 33264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_287
timestamp 1698431365
transform 1 0 33488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_37
timestamp 1698431365
transform 1 0 5488 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_79
timestamp 1698431365
transform 1 0 10192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_83
timestamp 1698431365
transform 1 0 10640 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_130
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_132
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_168
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_395
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_399
timestamp 1698431365
transform 1 0 46032 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_102
timestamp 1698431365
transform 1 0 12768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_104
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_152
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_156
timestamp 1698431365
transform 1 0 18816 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_288
timestamp 1698431365
transform 1 0 33600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_292
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_347
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_358
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_362
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_397
timestamp 1698431365
transform 1 0 45808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_401
timestamp 1698431365
transform 1 0 46256 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_60
timestamp 1698431365
transform 1 0 8064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_62
timestamp 1698431365
transform 1 0 8288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_65
timestamp 1698431365
transform 1 0 8624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_124
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_132
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698431365
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_272
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_280
timestamp 1698431365
transform 1 0 32704 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_297
timestamp 1698431365
transform 1 0 34608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_323
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_360
timestamp 1698431365
transform 1 0 41664 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_364
timestamp 1698431365
transform 1 0 42112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_366
timestamp 1698431365
transform 1 0 42336 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_393
timestamp 1698431365
transform 1 0 45360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_397
timestamp 1698431365
transform 1 0 45808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_401
timestamp 1698431365
transform 1 0 46256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_16
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_57
timestamp 1698431365
transform 1 0 7728 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_65
timestamp 1698431365
transform 1 0 8624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_316
timestamp 1698431365
transform 1 0 36736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_318
timestamp 1698431365
transform 1 0 36960 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_356
timestamp 1698431365
transform 1 0 41216 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_391
timestamp 1698431365
transform 1 0 45136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_399
timestamp 1698431365
transform 1 0 46032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_401
timestamp 1698431365
transform 1 0 46256 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_39
timestamp 1698431365
transform 1 0 5712 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_66
timestamp 1698431365
transform 1 0 8736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_70
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_119
timestamp 1698431365
transform 1 0 14672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_144
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_179
timestamp 1698431365
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_196
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_204
timestamp 1698431365
transform 1 0 24192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_261
timestamp 1698431365
transform 1 0 30576 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_268
timestamp 1698431365
transform 1 0 31360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_329
timestamp 1698431365
transform 1 0 38192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_399
timestamp 1698431365
transform 1 0 46032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_401
timestamp 1698431365
transform 1 0 46256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_78
timestamp 1698431365
transform 1 0 10080 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_86
timestamp 1698431365
transform 1 0 10976 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_127
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_153
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_161
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_198
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_272
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_398
timestamp 1698431365
transform 1 0 45920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_43
timestamp 1698431365
transform 1 0 6160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_57
timestamp 1698431365
transform 1 0 7728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_93
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_97
timestamp 1698431365
transform 1 0 12208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_286
timestamp 1698431365
transform 1 0 33376 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_294
timestamp 1698431365
transform 1 0 34272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_398
timestamp 1698431365
transform 1 0 45920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_10
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_53
timestamp 1698431365
transform 1 0 7280 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_61
timestamp 1698431365
transform 1 0 8176 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_74
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_103
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_105
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_218
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_226
timestamp 1698431365
transform 1 0 26656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_286
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_348
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_392
timestamp 1698431365
transform 1 0 45248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_26
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_49
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_51
timestamp 1698431365
transform 1 0 7056 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_58
timestamp 1698431365
transform 1 0 7840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_100
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_111
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_119
timestamp 1698431365
transform 1 0 14672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_163
timestamp 1698431365
transform 1 0 19600 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_209
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_213
timestamp 1698431365
transform 1 0 25200 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_217
timestamp 1698431365
transform 1 0 25648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_395
timestamp 1698431365
transform 1 0 45584 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_399
timestamp 1698431365
transform 1 0 46032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_401
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_19
timestamp 1698431365
transform 1 0 3472 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_27
timestamp 1698431365
transform 1 0 4368 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_148
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_289
timestamp 1698431365
transform 1 0 33712 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_297
timestamp 1698431365
transform 1 0 34608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_392
timestamp 1698431365
transform 1 0 45248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_399
timestamp 1698431365
transform 1 0 46032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_401
timestamp 1698431365
transform 1 0 46256 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_26
timestamp 1698431365
transform 1 0 4256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_113
timestamp 1698431365
transform 1 0 14000 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_126
timestamp 1698431365
transform 1 0 15456 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_161
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_218
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_226
timestamp 1698431365
transform 1 0 26656 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_319
timestamp 1698431365
transform 1 0 37072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_354
timestamp 1698431365
transform 1 0 40992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_358
timestamp 1698431365
transform 1 0 41440 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_362
timestamp 1698431365
transform 1 0 41888 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_399
timestamp 1698431365
transform 1 0 46032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_401
timestamp 1698431365
transform 1 0 46256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_40
timestamp 1698431365
transform 1 0 5824 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_44
timestamp 1698431365
transform 1 0 6272 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_79
timestamp 1698431365
transform 1 0 10192 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_129
timestamp 1698431365
transform 1 0 15792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_131
timestamp 1698431365
transform 1 0 16016 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_218
timestamp 1698431365
transform 1 0 25760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_254
timestamp 1698431365
transform 1 0 29792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_258
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_262
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_316
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_320
timestamp 1698431365
transform 1 0 37184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_324
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_393
timestamp 1698431365
transform 1 0 45360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_397
timestamp 1698431365
transform 1 0 45808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_6
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_23
timestamp 1698431365
transform 1 0 3920 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_31
timestamp 1698431365
transform 1 0 4816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_281
timestamp 1698431365
transform 1 0 32816 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_289
timestamp 1698431365
transform 1 0 33712 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_329
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_375
timestamp 1698431365
transform 1 0 43344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_399
timestamp 1698431365
transform 1 0 46032 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_401
timestamp 1698431365
transform 1 0 46256 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_8
timestamp 1698431365
transform 1 0 2240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_43
timestamp 1698431365
transform 1 0 6160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_65
timestamp 1698431365
transform 1 0 8624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_146
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_163
timestamp 1698431365
transform 1 0 19600 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_171
timestamp 1698431365
transform 1 0 20496 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_277
timestamp 1698431365
transform 1 0 32368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_304
timestamp 1698431365
transform 1 0 35392 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_320
timestamp 1698431365
transform 1 0 37184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_338
timestamp 1698431365
transform 1 0 39200 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_356
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_392
timestamp 1698431365
transform 1 0 45248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_400
timestamp 1698431365
transform 1 0 46144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_18
timestamp 1698431365
transform 1 0 3360 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_41
timestamp 1698431365
transform 1 0 5936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_61
timestamp 1698431365
transform 1 0 8176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_63
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_96
timestamp 1698431365
transform 1 0 12096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_100
timestamp 1698431365
transform 1 0 12544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_141
timestamp 1698431365
transform 1 0 17136 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_164
timestamp 1698431365
transform 1 0 19712 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_183
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_198
timestamp 1698431365
transform 1 0 23520 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_223
timestamp 1698431365
transform 1 0 26320 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_272
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_280
timestamp 1698431365
transform 1 0 32704 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_297
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_342
timestamp 1698431365
transform 1 0 39648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_344
timestamp 1698431365
transform 1 0 39872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_347
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_399
timestamp 1698431365
transform 1 0 46032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_401
timestamp 1698431365
transform 1 0 46256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_37
timestamp 1698431365
transform 1 0 5488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_41
timestamp 1698431365
transform 1 0 5936 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_49
timestamp 1698431365
transform 1 0 6832 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_53
timestamp 1698431365
transform 1 0 7280 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_91
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_95
timestamp 1698431365
transform 1 0 11984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_131
timestamp 1698431365
transform 1 0 16016 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_167
timestamp 1698431365
transform 1 0 20048 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_175
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_177
timestamp 1698431365
transform 1 0 21168 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_194
timestamp 1698431365
transform 1 0 23072 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_237
timestamp 1698431365
transform 1 0 27888 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_245
timestamp 1698431365
transform 1 0 28784 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_268
timestamp 1698431365
transform 1 0 31360 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_300
timestamp 1698431365
transform 1 0 34944 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_316
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_318
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_335
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_343
timestamp 1698431365
transform 1 0 39760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_347
timestamp 1698431365
transform 1 0 40208 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_358
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_395
timestamp 1698431365
transform 1 0 45584 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_399
timestamp 1698431365
transform 1 0 46032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_401
timestamp 1698431365
transform 1 0 46256 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_49
timestamp 1698431365
transform 1 0 6832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_67
timestamp 1698431365
transform 1 0 8848 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_83
timestamp 1698431365
transform 1 0 10640 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_87
timestamp 1698431365
transform 1 0 11088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_117
timestamp 1698431365
transform 1 0 14448 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_134
timestamp 1698431365
transform 1 0 16352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_138
timestamp 1698431365
transform 1 0 16800 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_142
timestamp 1698431365
transform 1 0 17248 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_159
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_202
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_210
timestamp 1698431365
transform 1 0 24864 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_227
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_283
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_342
timestamp 1698431365
transform 1 0 39648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_350
timestamp 1698431365
transform 1 0 40544 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_367
timestamp 1698431365
transform 1 0 42448 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_399
timestamp 1698431365
transform 1 0 46032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_401
timestamp 1698431365
transform 1 0 46256 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_26
timestamp 1698431365
transform 1 0 4256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_30
timestamp 1698431365
transform 1 0 4704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_32
timestamp 1698431365
transform 1 0 4928 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_49
timestamp 1698431365
transform 1 0 6832 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_65
timestamp 1698431365
transform 1 0 8624 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_112
timestamp 1698431365
transform 1 0 13888 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_116
timestamp 1698431365
transform 1 0 14336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_176
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_184
timestamp 1698431365
transform 1 0 21952 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_356
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_358
timestamp 1698431365
transform 1 0 41440 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_395
timestamp 1698431365
transform 1 0 45584 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_399
timestamp 1698431365
transform 1 0 46032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_401
timestamp 1698431365
transform 1 0 46256 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_135
timestamp 1698431365
transform 1 0 16464 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_151
timestamp 1698431365
transform 1 0 18256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_153
timestamp 1698431365
transform 1 0 18480 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_203
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_235
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_334
timestamp 1698431365
transform 1 0 38752 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_350
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_368
timestamp 1698431365
transform 1 0 42560 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_395
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_399
timestamp 1698431365
transform 1 0 46032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_401
timestamp 1698431365
transform 1 0 46256 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_104
timestamp 1698431365
transform 1 0 12992 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_108
timestamp 1698431365
transform 1 0 13440 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_125
timestamp 1698431365
transform 1 0 15344 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_190
timestamp 1698431365
transform 1 0 22624 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_314
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_322
timestamp 1698431365
transform 1 0 37408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_324
timestamp 1698431365
transform 1 0 37632 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_341
timestamp 1698431365
transform 1 0 39536 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_364
timestamp 1698431365
transform 1 0 42112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_382
timestamp 1698431365
transform 1 0 44128 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_398
timestamp 1698431365
transform 1 0 45920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_139
timestamp 1698431365
transform 1 0 16912 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_143
timestamp 1698431365
transform 1 0 17360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_145
timestamp 1698431365
transform 1 0 17584 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_162
timestamp 1698431365
transform 1 0 19488 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_170
timestamp 1698431365
transform 1 0 20384 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_353
timestamp 1698431365
transform 1 0 40880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_355
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_372
timestamp 1698431365
transform 1 0 43008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_380
timestamp 1698431365
transform 1 0 43904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_395
timestamp 1698431365
transform 1 0 45584 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_399
timestamp 1698431365
transform 1 0 46032 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_401
timestamp 1698431365
transform 1 0 46256 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_360
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_377
timestamp 1698431365
transform 1 0 43568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_385
timestamp 1698431365
transform 1 0 44464 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_349
timestamp 1698431365
transform 1 0 40432 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_357
timestamp 1698431365
transform 1 0 41328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_359
timestamp 1698431365
transform 1 0 41552 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_376
timestamp 1698431365
transform 1 0 43456 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_397
timestamp 1698431365
transform 1 0 45808 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_368
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_376
timestamp 1698431365
transform 1 0 43456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_380
timestamp 1698431365
transform 1 0 43904 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_401
timestamp 1698431365
transform 1 0 46256 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_393
timestamp 1698431365
transform 1 0 45360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_395
timestamp 1698431365
transform 1 0 45584 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_220
timestamp 1698431365
transform 1 0 25984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_224
timestamp 1698431365
transform 1 0 26432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_244
timestamp 1698431365
transform 1 0 28672 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_252
timestamp 1698431365
transform 1 0 29568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_262
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_278
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_314
timestamp 1698431365
transform 1 0 36512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_324
timestamp 1698431365
transform 1 0 37632 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_328
timestamp 1698431365
transform 1 0 38080 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_336
timestamp 1698431365
transform 1 0 38976 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_368
timestamp 1698431365
transform 1 0 42560 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_376
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_393
timestamp 1698431365
transform 1 0 45360 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_397
timestamp 1698431365
transform 1 0 45808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_399
timestamp 1698431365
transform 1 0 46032 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_6
timestamp 1698431365
transform 1 0 2016 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_22
timestamp 1698431365
transform 1 0 3808 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_30
timestamp 1698431365
transform 1 0 4704 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_59
timestamp 1698431365
transform 1 0 7952 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_91
timestamp 1698431365
transform 1 0 11536 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_99
timestamp 1698431365
transform 1 0 12432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_116
timestamp 1698431365
transform 1 0 14336 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_148
timestamp 1698431365
transform 1 0 17920 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_151
timestamp 1698431365
transform 1 0 18256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_161
timestamp 1698431365
transform 1 0 19376 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_191
timestamp 1698431365
transform 1 0 22736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_193
timestamp 1698431365
transform 1 0 22960 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_200
timestamp 1698431365
transform 1 0 23744 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_208
timestamp 1698431365
transform 1 0 24640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_212
timestamp 1698431365
transform 1 0 25088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_214
timestamp 1698431365
transform 1 0 25312 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_227
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_327
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_352
timestamp 1698431365
transform 1 0 40768 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_368
timestamp 1698431365
transform 1 0 42560 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_376
timestamp 1698431365
transform 1 0 43456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_378
timestamp 1698431365
transform 1 0 43680 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_398
timestamp 1698431365
transform 1 0 45920 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_144
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_149
timestamp 1698431365
transform 1 0 18032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_163
timestamp 1698431365
transform 1 0 19600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_167
timestamp 1698431365
transform 1 0 20048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_171
timestamp 1698431365
transform 1 0 20496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_197
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_218
timestamp 1698431365
transform 1 0 25760 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_222
timestamp 1698431365
transform 1 0 26208 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_233
timestamp 1698431365
transform 1 0 27440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_237
timestamp 1698431365
transform 1 0 27888 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_251
timestamp 1698431365
transform 1 0 29456 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_265
timestamp 1698431365
transform 1 0 31024 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_290
timestamp 1698431365
transform 1 0 33824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_292
timestamp 1698431365
transform 1 0 34048 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_295
timestamp 1698431365
transform 1 0 34384 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_307
timestamp 1698431365
transform 1 0 35728 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_323
timestamp 1698431365
transform 1 0 37520 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_327
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_339
timestamp 1698431365
transform 1 0 39312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_354
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_365
timestamp 1698431365
transform 1 0 42224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_375
timestamp 1698431365
transform 1 0 43344 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_383
timestamp 1698431365
transform 1 0 44240 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_387
timestamp 1698431365
transform 1 0 44688 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_36
timestamp 1698431365
transform 1 0 5376 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_52
timestamp 1698431365
transform 1 0 7168 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_61
timestamp 1698431365
transform 1 0 8176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_65
timestamp 1698431365
transform 1 0 8624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_67
timestamp 1698431365
transform 1 0 8848 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_80
timestamp 1698431365
transform 1 0 10304 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_96
timestamp 1698431365
transform 1 0 12096 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_106
timestamp 1698431365
transform 1 0 13216 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_125
timestamp 1698431365
transform 1 0 15344 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_133
timestamp 1698431365
transform 1 0 16240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_135
timestamp 1698431365
transform 1 0 16464 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_138
timestamp 1698431365
transform 1 0 16800 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_153
timestamp 1698431365
transform 1 0 18480 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_155
timestamp 1698431365
transform 1 0 18704 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_186
timestamp 1698431365
transform 1 0 22176 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_206
timestamp 1698431365
transform 1 0 24416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_210
timestamp 1698431365
transform 1 0 24864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_212
timestamp 1698431365
transform 1 0 25088 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_237
timestamp 1698431365
transform 1 0 27888 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_250
timestamp 1698431365
transform 1 0 29344 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_264
timestamp 1698431365
transform 1 0 30912 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_284
timestamp 1698431365
transform 1 0 33152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_294
timestamp 1698431365
transform 1 0 34272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_301
timestamp 1698431365
transform 1 0 35056 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_305
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_339
timestamp 1698431365
transform 1 0 39312 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_352
timestamp 1698431365
transform 1 0 40768 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_366
timestamp 1698431365
transform 1 0 42336 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_386
timestamp 1698431365
transform 1 0 44576 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform 1 0 33152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 16464 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 17136 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 44128 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform 1 0 1680 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 39200 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 34608 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform 1 0 2128 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 44464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform 1 0 22064 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 36736 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 35616 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 36288 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform 1 0 13440 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 27888 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 42784 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform 1 0 21280 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 36176 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 24080 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 22064 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 28560 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform -1 0 42560 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 26320 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 36288 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform 1 0 21504 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform -1 0 12096 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 16352 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform 1 0 37072 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 27888 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 28224 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 46368 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform -1 0 44240 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform 1 0 14784 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 31808 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 39648 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform -1 0 7392 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform -1 0 14224 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold50
timestamp 1698431365
transform 1 0 6384 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform -1 0 43568 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform -1 0 43456 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform -1 0 39984 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 14224 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform -1 0 28224 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 39088 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform -1 0 43904 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform -1 0 43904 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform -1 0 20384 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform -1 0 42896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform -1 0 43568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform -1 0 39648 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 21056 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform 1 0 29120 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform -1 0 31808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold69
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold70
timestamp 1698431365
transform -1 0 34720 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold71
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold72
timestamp 1698431365
transform -1 0 11872 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold73
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold74
timestamp 1698431365
transform -1 0 31920 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold75
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold76
timestamp 1698431365
transform -1 0 19152 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold77
timestamp 1698431365
transform -1 0 10304 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold78
timestamp 1698431365
transform -1 0 36064 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold79
timestamp 1698431365
transform -1 0 46368 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold80
timestamp 1698431365
transform -1 0 46368 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold81
timestamp 1698431365
transform -1 0 8288 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold82
timestamp 1698431365
transform -1 0 26880 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold83
timestamp 1698431365
transform -1 0 35616 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold84
timestamp 1698431365
transform -1 0 39760 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold85
timestamp 1698431365
transform -1 0 16352 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold86
timestamp 1698431365
transform -1 0 46368 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold87
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold88
timestamp 1698431365
transform -1 0 35056 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold89
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold90
timestamp 1698431365
transform 1 0 2128 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold91
timestamp 1698431365
transform 1 0 2128 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold92
timestamp 1698431365
transform 1 0 37744 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold93
timestamp 1698431365
transform -1 0 45808 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold94
timestamp 1698431365
transform 1 0 31248 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold95
timestamp 1698431365
transform 1 0 13552 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold96
timestamp 1698431365
transform -1 0 34608 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold97
timestamp 1698431365
transform -1 0 19488 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold98
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold99
timestamp 1698431365
transform -1 0 32592 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold100
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold101
timestamp 1698431365
transform 1 0 2464 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold102
timestamp 1698431365
transform -1 0 4032 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold103
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold104
timestamp 1698431365
transform -1 0 28672 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold105
timestamp 1698431365
transform -1 0 43008 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold106
timestamp 1698431365
transform 1 0 6272 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold107
timestamp 1698431365
transform -1 0 31024 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold108
timestamp 1698431365
transform -1 0 16912 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold109
timestamp 1698431365
transform -1 0 5264 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold110
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold111
timestamp 1698431365
transform -1 0 43792 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold112
timestamp 1698431365
transform -1 0 12208 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold113
timestamp 1698431365
transform -1 0 16016 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold114
timestamp 1698431365
transform -1 0 30688 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold115
timestamp 1698431365
transform -1 0 41888 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold116
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold117
timestamp 1698431365
transform 1 0 17808 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold118
timestamp 1698431365
transform 1 0 6384 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold119
timestamp 1698431365
transform 1 0 41664 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold120
timestamp 1698431365
transform -1 0 37856 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold121
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold122
timestamp 1698431365
transform -1 0 27888 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold123
timestamp 1698431365
transform -1 0 34384 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold124
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold125
timestamp 1698431365
transform -1 0 13664 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold126
timestamp 1698431365
transform -1 0 42784 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold127
timestamp 1698431365
transform -1 0 42560 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold128
timestamp 1698431365
transform -1 0 39648 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold129
timestamp 1698431365
transform -1 0 26768 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold130
timestamp 1698431365
transform -1 0 20272 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold131
timestamp 1698431365
transform -1 0 39536 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold132
timestamp 1698431365
transform -1 0 8064 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold133
timestamp 1698431365
transform 1 0 11424 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold134
timestamp 1698431365
transform 1 0 14224 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold135
timestamp 1698431365
transform -1 0 42448 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold136
timestamp 1698431365
transform 1 0 6272 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold137
timestamp 1698431365
transform -1 0 46368 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold138
timestamp 1698431365
transform 1 0 10304 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold139
timestamp 1698431365
transform -1 0 23968 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold140
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold141
timestamp 1698431365
transform -1 0 24640 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold142
timestamp 1698431365
transform -1 0 16016 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold143
timestamp 1698431365
transform -1 0 45808 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold144
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold145
timestamp 1698431365
transform 1 0 7056 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold146
timestamp 1698431365
transform -1 0 6832 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold147
timestamp 1698431365
transform -1 0 43568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold148
timestamp 1698431365
transform 1 0 36960 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold149
timestamp 1698431365
transform 1 0 43568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold150
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold151
timestamp 1698431365
transform -1 0 39648 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold152
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold153
timestamp 1698431365
transform -1 0 8624 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold154
timestamp 1698431365
transform -1 0 39984 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold155
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold156
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold157
timestamp 1698431365
transform 1 0 8960 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold158
timestamp 1698431365
transform -1 0 20048 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 42448 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 6720 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 18928 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 14224 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 27888 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 10752 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 34272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 31024 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 24528 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 46368 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 19600 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 46368 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 40432 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 31696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 23184 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 27216 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 31696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 20944 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 34608 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 9520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 27216 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 19600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 34384 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 17808 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 35056 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 35056 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform -1 0 46368 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 43792 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform -1 0 36400 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 35280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform -1 0 31024 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform -1 0 45696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform -1 0 43344 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform -1 0 27888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform -1 0 39312 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform -1 0 8176 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 38640 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform -1 0 32368 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 43792 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform -1 0 43008 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform -1 0 46368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform -1 0 22288 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform -1 0 46256 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 39760 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input62 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46368 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output63 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44800 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output64
timestamp 1698431365
transform 1 0 20944 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform -1 0 18480 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform -1 0 9072 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform 1 0 44800 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 41216 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output69
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output70
timestamp 1698431365
transform 1 0 32368 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output71
timestamp 1698431365
transform -1 0 22736 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44800 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output73
timestamp 1698431365
transform 1 0 26320 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output74
timestamp 1698431365
transform 1 0 29904 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output75 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output76
timestamp 1698431365
transform 1 0 36400 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output77
timestamp 1698431365
transform 1 0 24304 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output78
timestamp 1698431365
transform 1 0 26320 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output79
timestamp 1698431365
transform -1 0 24192 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output80
timestamp 1698431365
transform 1 0 28336 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output81
timestamp 1698431365
transform -1 0 13328 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output82
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output83
timestamp 1698431365
transform -1 0 18816 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output84
timestamp 1698431365
transform -1 0 26544 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output85
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output86
timestamp 1698431365
transform -1 0 10752 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output87
timestamp 1698431365
transform 1 0 24976 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output88
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output89
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output90
timestamp 1698431365
transform 1 0 29792 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output91
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output92
timestamp 1698431365
transform 1 0 28224 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output93
timestamp 1698431365
transform 1 0 32032 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output94
timestamp 1698431365
transform -1 0 14112 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output95
timestamp 1698431365
transform 1 0 39648 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output96
timestamp 1698431365
transform 1 0 28336 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output97
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output98
timestamp 1698431365
transform -1 0 3136 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output99
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output100
timestamp 1698431365
transform 1 0 44800 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output101
timestamp 1698431365
transform -1 0 20384 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output102
timestamp 1698431365
transform 1 0 9184 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output103
timestamp 1698431365
transform 1 0 22288 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output104
timestamp 1698431365
transform 1 0 44800 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output105
timestamp 1698431365
transform 1 0 42896 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output106
timestamp 1698431365
transform 1 0 43456 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output107
timestamp 1698431365
transform -1 0 3136 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output108
timestamp 1698431365
transform 1 0 41216 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output109
timestamp 1698431365
transform 1 0 44800 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output110
timestamp 1698431365
transform -1 0 3136 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output111
timestamp 1698431365
transform -1 0 3136 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output112
timestamp 1698431365
transform 1 0 44800 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output113
timestamp 1698431365
transform -1 0 37968 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output114
timestamp 1698431365
transform 1 0 44800 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output115
timestamp 1698431365
transform 1 0 44800 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output116
timestamp 1698431365
transform -1 0 46368 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output117
timestamp 1698431365
transform -1 0 39312 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output118
timestamp 1698431365
transform 1 0 44800 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output119
timestamp 1698431365
transform 1 0 44800 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output120
timestamp 1698431365
transform 1 0 44800 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output121
timestamp 1698431365
transform 1 0 44800 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output122
timestamp 1698431365
transform 1 0 41104 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output123
timestamp 1698431365
transform 1 0 44800 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_53 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 46592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 46592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 46592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 46592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 46592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 46592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 46592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 46592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 46592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 46592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 46592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 46592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 46592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 46592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 46592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 46592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 46592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 46592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 46592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 46592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 46592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 46592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 46592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 46592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 46592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 46592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 46592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 46592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 46592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 46592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 46592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 46592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 46592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 46592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 46592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 46592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 46592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 46592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 46592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 46592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 46592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 46592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 46592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 46592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 46592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 46592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 46592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 46592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__124 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__125
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__126
timestamp 1698431365
transform -1 0 36288 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__127
timestamp 1698431365
transform 1 0 44128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__128
timestamp 1698431365
transform -1 0 18032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__129
timestamp 1698431365
transform 1 0 43792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__130
timestamp 1698431365
transform 1 0 43344 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__131
timestamp 1698431365
transform 1 0 45920 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__132
timestamp 1698431365
transform 1 0 44576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__133
timestamp 1698431365
transform -1 0 36288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__134
timestamp 1698431365
transform 1 0 43344 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__135
timestamp 1698431365
transform -1 0 30352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__136
timestamp 1698431365
transform -1 0 2688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__137
timestamp 1698431365
transform -1 0 29456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__138
timestamp 1698431365
transform 1 0 45808 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__139
timestamp 1698431365
transform -1 0 16240 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__140
timestamp 1698431365
transform -1 0 18704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__141
timestamp 1698431365
transform -1 0 2016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__142
timestamp 1698431365
transform 1 0 45024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__1__143
timestamp 1698431365
transform -1 0 10640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_117
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_118
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_119
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_120
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_121
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_122
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_123
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_124
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_125
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_126
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_128
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_129
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_130
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_131
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_133
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_134
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_135
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_136
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_137
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_139
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_140
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_141
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_142
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_143
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_144
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_145
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_146
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_147
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_148
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_150
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_151
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_152
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_153
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_154
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_155
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_156
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_157
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_158
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_159
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_161
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_162
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_163
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_164
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_165
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_166
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_167
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_168
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_169
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_170
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_172
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_173
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_174
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_175
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_176
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_177
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_178
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_179
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_180
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_181
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_183
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_184
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_191
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_192
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_194
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_195
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_196
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_197
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_198
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_199
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_200
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_201
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_202
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_203
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_205
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_206
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_207
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_208
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_209
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_210
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_211
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_212
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_213
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_214
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_216
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_217
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_218
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_219
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_220
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_221
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_222
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_223
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_224
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_225
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_227
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_228
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_229
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_230
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_231
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_232
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_233
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_234
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_235
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_236
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_238
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_239
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_240
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_241
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_242
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_243
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_244
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_245
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_246
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_247
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_249
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_250
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_251
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_252
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_253
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_254
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_255
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_256
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_257
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_258
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_260
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_261
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_262
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_263
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_264
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_265
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_266
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_267
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_268
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_269
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_271
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_272
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_273
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_274
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_275
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_276
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_277
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_278
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_279
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_280
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_282
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_283
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_284
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_285
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_286
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_287
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_288
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_289
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_290
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_291
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_293
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_294
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_295
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_296
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_297
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_298
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_299
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_300
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_301
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_302
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_304
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_305
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_306
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_307
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_308
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_309
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_310
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_311
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_312
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_313
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_315
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_316
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_317
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_318
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_319
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_320
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_321
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_322
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_323
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_324
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_326
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_327
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_328
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_329
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_330
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_331
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_332
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_333
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_334
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_335
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_337
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_338
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_339
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_340
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_341
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_342
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_343
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_344
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_345
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_346
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_348
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_349
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_350
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_351
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_352
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_353
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_354
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_355
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_356
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_357
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_359
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_360
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_361
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_362
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_363
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_364
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_365
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_366
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_367
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_368
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_370
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_371
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_372
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_373
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_374
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_375
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_376
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_377
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_378
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_379
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_381
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_382
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_383
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_384
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_385
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_386
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_387
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_388
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_389
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_390
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_392
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_393
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_394
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_395
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_396
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_397
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_398
timestamp 1698431365
transform 1 0 8960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_399
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_400
timestamp 1698431365
transform 1 0 16576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_401
timestamp 1698431365
transform 1 0 20384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 24192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 31808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 39424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 43232 0 1 43904
box -86 -86 310 870
<< labels >>
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 2 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 3 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 47200 26208 48000 26320 0 FreeSans 448 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 24192 47200 24304 48000 0 FreeSans 448 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal2 s 13440 47200 13552 48000 0 FreeSans 448 90 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chanx_left_in[2]
port 18 nsew signal input
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 chanx_left_in[3]
port 19 nsew signal input
flabel metal2 s 26880 47200 26992 48000 0 FreeSans 448 90 0 0 chanx_left_in[4]
port 20 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chanx_left_in[5]
port 21 nsew signal input
flabel metal2 s 32256 47200 32368 48000 0 FreeSans 448 90 0 0 chanx_left_in[6]
port 22 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 chanx_left_in[7]
port 23 nsew signal input
flabel metal2 s 30240 47200 30352 48000 0 FreeSans 448 90 0 0 chanx_left_in[8]
port 24 nsew signal input
flabel metal2 s 22848 47200 22960 48000 0 FreeSans 448 90 0 0 chanx_left_in[9]
port 25 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chanx_left_out[0]
port 26 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 chanx_left_out[10]
port 27 nsew signal tristate
flabel metal2 s 16800 47200 16912 48000 0 FreeSans 448 90 0 0 chanx_left_out[11]
port 28 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chanx_left_out[12]
port 29 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 chanx_left_out[13]
port 30 nsew signal tristate
flabel metal3 s 47200 44352 48000 44464 0 FreeSans 448 0 0 0 chanx_left_out[14]
port 31 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 chanx_left_out[15]
port 32 nsew signal tristate
flabel metal2 s 14784 47200 14896 48000 0 FreeSans 448 90 0 0 chanx_left_out[16]
port 33 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 chanx_left_out[17]
port 34 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 chanx_left_out[18]
port 35 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 chanx_left_out[19]
port 36 nsew signal tristate
flabel metal3 s 47200 43008 48000 43120 0 FreeSans 448 0 0 0 chanx_left_out[1]
port 37 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 chanx_left_out[2]
port 38 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 chanx_left_out[3]
port 39 nsew signal tristate
flabel metal3 s 47200 2688 48000 2800 0 FreeSans 448 0 0 0 chanx_left_out[4]
port 40 nsew signal tristate
flabel metal2 s 20160 47200 20272 48000 0 FreeSans 448 90 0 0 chanx_left_out[5]
port 41 nsew signal tristate
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 chanx_left_out[6]
port 42 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 chanx_left_out[7]
port 43 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 chanx_left_out[8]
port 44 nsew signal tristate
flabel metal2 s 26208 47200 26320 48000 0 FreeSans 448 90 0 0 chanx_left_out[9]
port 45 nsew signal tristate
flabel metal3 s 47200 40992 48000 41104 0 FreeSans 448 0 0 0 chanx_right_in[0]
port 46 nsew signal input
flabel metal2 s 18816 47200 18928 48000 0 FreeSans 448 90 0 0 chanx_right_in[10]
port 47 nsew signal input
flabel metal2 s 46368 0 46480 800 0 FreeSans 448 90 0 0 chanx_right_in[11]
port 48 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 chanx_right_in[12]
port 49 nsew signal input
flabel metal3 s 47200 43680 48000 43792 0 FreeSans 448 0 0 0 chanx_right_in[13]
port 50 nsew signal input
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 chanx_right_in[14]
port 51 nsew signal input
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 chanx_right_in[15]
port 52 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 chanx_right_in[16]
port 53 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 chanx_right_in[17]
port 54 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 chanx_right_in[18]
port 55 nsew signal input
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 chanx_right_in[19]
port 56 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 chanx_right_in[1]
port 57 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 chanx_right_in[2]
port 58 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 chanx_right_in[3]
port 59 nsew signal input
flabel metal2 s 20832 47200 20944 48000 0 FreeSans 448 90 0 0 chanx_right_in[4]
port 60 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 chanx_right_in[5]
port 61 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 chanx_right_in[6]
port 62 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 chanx_right_in[7]
port 63 nsew signal input
flabel metal2 s 25536 47200 25648 48000 0 FreeSans 448 90 0 0 chanx_right_in[8]
port 64 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 chanx_right_in[9]
port 65 nsew signal input
flabel metal3 s 47200 42336 48000 42448 0 FreeSans 448 0 0 0 chanx_right_out[0]
port 66 nsew signal tristate
flabel metal2 s 23520 47200 23632 48000 0 FreeSans 448 90 0 0 chanx_right_out[10]
port 67 nsew signal tristate
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 chanx_right_out[11]
port 68 nsew signal tristate
flabel metal2 s 28896 47200 29008 48000 0 FreeSans 448 90 0 0 chanx_right_out[12]
port 69 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chanx_right_out[13]
port 70 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chanx_right_out[14]
port 71 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chanx_right_out[15]
port 72 nsew signal tristate
flabel metal3 s 47200 4032 48000 4144 0 FreeSans 448 0 0 0 chanx_right_out[16]
port 73 nsew signal tristate
flabel metal2 s 24864 47200 24976 48000 0 FreeSans 448 90 0 0 chanx_right_out[17]
port 74 nsew signal tristate
flabel metal2 s 14112 47200 14224 48000 0 FreeSans 448 90 0 0 chanx_right_out[18]
port 75 nsew signal tristate
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chanx_right_out[19]
port 76 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 chanx_right_out[1]
port 77 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chanx_right_out[2]
port 78 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 chanx_right_out[3]
port 79 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 chanx_right_out[4]
port 80 nsew signal tristate
flabel metal2 s 29568 47200 29680 48000 0 FreeSans 448 90 0 0 chanx_right_out[5]
port 81 nsew signal tristate
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chanx_right_out[6]
port 82 nsew signal tristate
flabel metal2 s 27552 47200 27664 48000 0 FreeSans 448 90 0 0 chanx_right_out[7]
port 83 nsew signal tristate
flabel metal3 s 0 2688 800 2800 0 FreeSans 448 0 0 0 chanx_right_out[8]
port 84 nsew signal tristate
flabel metal2 s 30912 47200 31024 48000 0 FreeSans 448 90 0 0 chanx_right_out[9]
port 85 nsew signal tristate
flabel metal2 s 34272 47200 34384 48000 0 FreeSans 448 90 0 0 chany_bottom_in[0]
port 86 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chany_bottom_in[10]
port 87 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 chany_bottom_in[11]
port 88 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 chany_bottom_in[12]
port 89 nsew signal input
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 chany_bottom_in[13]
port 90 nsew signal input
flabel metal2 s 34944 47200 35056 48000 0 FreeSans 448 90 0 0 chany_bottom_in[14]
port 91 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 chany_bottom_in[15]
port 92 nsew signal input
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 chany_bottom_in[16]
port 93 nsew signal input
flabel metal3 s 47200 19488 48000 19600 0 FreeSans 448 0 0 0 chany_bottom_in[17]
port 94 nsew signal input
flabel metal3 s 47200 10752 48000 10864 0 FreeSans 448 0 0 0 chany_bottom_in[18]
port 95 nsew signal input
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 chany_bottom_in[19]
port 96 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 chany_bottom_in[1]
port 97 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 chany_bottom_in[2]
port 98 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 chany_bottom_in[3]
port 99 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 chany_bottom_in[4]
port 100 nsew signal input
flabel metal3 s 47200 5376 48000 5488 0 FreeSans 448 0 0 0 chany_bottom_in[5]
port 101 nsew signal input
flabel metal2 s 41664 47200 41776 48000 0 FreeSans 448 90 0 0 chany_bottom_in[6]
port 102 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 chany_bottom_in[7]
port 103 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 chany_bottom_in[8]
port 104 nsew signal input
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 chany_bottom_in[9]
port 105 nsew signal input
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 chany_bottom_out[0]
port 106 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 chany_bottom_out[10]
port 107 nsew signal tristate
flabel metal2 s 38976 47200 39088 48000 0 FreeSans 448 90 0 0 chany_bottom_out[11]
port 108 nsew signal tristate
flabel metal3 s 47200 4704 48000 4816 0 FreeSans 448 0 0 0 chany_bottom_out[12]
port 109 nsew signal tristate
flabel metal2 s 28224 47200 28336 48000 0 FreeSans 448 90 0 0 chany_bottom_out[13]
port 110 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 chany_bottom_out[14]
port 111 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 chany_bottom_out[15]
port 112 nsew signal tristate
flabel metal3 s 47200 1344 48000 1456 0 FreeSans 448 0 0 0 chany_bottom_out[16]
port 113 nsew signal tristate
flabel metal3 s 47200 14112 48000 14224 0 FreeSans 448 0 0 0 chany_bottom_out[17]
port 114 nsew signal tristate
flabel metal3 s 47200 15456 48000 15568 0 FreeSans 448 0 0 0 chany_bottom_out[18]
port 115 nsew signal tristate
flabel metal2 s 19488 47200 19600 48000 0 FreeSans 448 90 0 0 chany_bottom_out[19]
port 116 nsew signal tristate
flabel metal2 s 8064 47200 8176 48000 0 FreeSans 448 90 0 0 chany_bottom_out[1]
port 117 nsew signal tristate
flabel metal2 s 22176 47200 22288 48000 0 FreeSans 448 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal3 s 47200 18144 48000 18256 0 FreeSans 448 0 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal3 s 47200 672 48000 784 0 FreeSans 448 0 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal3 s 47200 13440 48000 13552 0 FreeSans 448 0 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 42336 47200 42448 48000 0 FreeSans 448 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal3 s 47200 41664 48000 41776 0 FreeSans 448 0 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 40320 47200 40432 48000 0 FreeSans 448 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 7392 47200 7504 48000 0 FreeSans 448 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 38304 47200 38416 48000 0 FreeSans 448 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal3 s 47200 24192 48000 24304 0 FreeSans 448 0 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 31584 47200 31696 48000 0 FreeSans 448 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal3 s 47200 9408 48000 9520 0 FreeSans 448 0 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal3 s 47200 32256 48000 32368 0 FreeSans 448 0 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal3 s 47200 12768 48000 12880 0 FreeSans 448 0 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal3 s 47200 6048 48000 6160 0 FreeSans 448 0 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 18144 47200 18256 48000 0 FreeSans 448 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal3 s 47200 25536 48000 25648 0 FreeSans 448 0 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 21504 47200 21616 48000 0 FreeSans 448 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal3 s 47200 10080 48000 10192 0 FreeSans 448 0 0 0 chany_top_in[2]
port 138 nsew signal input
flabel metal3 s 47200 22848 48000 22960 0 FreeSans 448 0 0 0 chany_top_in[3]
port 139 nsew signal input
flabel metal3 s 47200 8736 48000 8848 0 FreeSans 448 0 0 0 chany_top_in[4]
port 140 nsew signal input
flabel metal2 s 36960 47200 37072 48000 0 FreeSans 448 90 0 0 chany_top_in[5]
port 141 nsew signal input
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 chany_top_in[6]
port 142 nsew signal input
flabel metal3 s 47200 28224 48000 28336 0 FreeSans 448 0 0 0 chany_top_in[7]
port 143 nsew signal input
flabel metal2 s 39648 47200 39760 48000 0 FreeSans 448 90 0 0 chany_top_in[8]
port 144 nsew signal input
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 chany_top_in[9]
port 145 nsew signal input
flabel metal2 s 17472 47200 17584 48000 0 FreeSans 448 90 0 0 chany_top_out[0]
port 146 nsew signal tristate
flabel metal3 s 47200 7392 48000 7504 0 FreeSans 448 0 0 0 chany_top_out[10]
port 147 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 chany_top_out[11]
port 148 nsew signal tristate
flabel metal3 s 47200 3360 48000 3472 0 FreeSans 448 0 0 0 chany_top_out[12]
port 149 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 chany_top_out[13]
port 150 nsew signal tristate
flabel metal3 s 47200 12096 48000 12208 0 FreeSans 448 0 0 0 chany_top_out[14]
port 151 nsew signal tristate
flabel metal2 s 36288 47200 36400 48000 0 FreeSans 448 90 0 0 chany_top_out[15]
port 152 nsew signal tristate
flabel metal3 s 47200 0 48000 112 0 FreeSans 448 0 0 0 chany_top_out[16]
port 153 nsew signal tristate
flabel metal3 s 47200 6720 48000 6832 0 FreeSans 448 0 0 0 chany_top_out[17]
port 154 nsew signal tristate
flabel metal3 s 47200 17472 48000 17584 0 FreeSans 448 0 0 0 chany_top_out[18]
port 155 nsew signal tristate
flabel metal3 s 47200 16128 48000 16240 0 FreeSans 448 0 0 0 chany_top_out[19]
port 156 nsew signal tristate
flabel metal2 s 37632 47200 37744 48000 0 FreeSans 448 90 0 0 chany_top_out[1]
port 157 nsew signal tristate
flabel metal3 s 47200 14784 48000 14896 0 FreeSans 448 0 0 0 chany_top_out[2]
port 158 nsew signal tristate
flabel metal3 s 47200 8064 48000 8176 0 FreeSans 448 0 0 0 chany_top_out[3]
port 159 nsew signal tristate
flabel metal3 s 47200 2016 48000 2128 0 FreeSans 448 0 0 0 chany_top_out[4]
port 160 nsew signal tristate
flabel metal3 s 47200 11424 48000 11536 0 FreeSans 448 0 0 0 chany_top_out[5]
port 161 nsew signal tristate
flabel metal3 s 47200 16800 48000 16912 0 FreeSans 448 0 0 0 chany_top_out[6]
port 162 nsew signal tristate
flabel metal2 s 40992 47200 41104 48000 0 FreeSans 448 90 0 0 chany_top_out[7]
port 163 nsew signal tristate
flabel metal2 s 35616 47200 35728 48000 0 FreeSans 448 90 0 0 chany_top_out[8]
port 164 nsew signal tristate
flabel metal3 s 47200 18816 48000 18928 0 FreeSans 448 0 0 0 chany_top_out[9]
port 165 nsew signal tristate
flabel metal3 s 47200 21504 48000 21616 0 FreeSans 448 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 166 nsew signal input
flabel metal3 s 47200 30912 48000 31024 0 FreeSans 448 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 167 nsew signal input
flabel metal3 s 47200 30240 48000 30352 0 FreeSans 448 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 168 nsew signal input
flabel metal3 s 47200 28896 48000 29008 0 FreeSans 448 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 169 nsew signal input
flabel metal3 s 47200 26880 48000 26992 0 FreeSans 448 0 0 0 pReset
port 170 nsew signal input
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 prog_clk
port 171 nsew signal input
flabel metal3 s 47200 31584 48000 31696 0 FreeSans 448 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 172 nsew signal input
flabel metal3 s 47200 27552 48000 27664 0 FreeSans 448 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 173 nsew signal input
flabel metal3 s 47200 29568 48000 29680 0 FreeSans 448 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 174 nsew signal input
flabel metal3 s 47200 20832 48000 20944 0 FreeSans 448 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 175 nsew signal input
flabel metal3 s 47200 22176 48000 22288 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 176 nsew signal input
flabel metal3 s 47200 23520 48000 23632 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 177 nsew signal input
flabel metal3 s 47200 20160 48000 20272 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 178 nsew signal input
flabel metal3 s 47200 24864 48000 24976 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 179 nsew signal input
flabel metal4 s 4448 3076 4768 44748 0 FreeSans 1280 90 0 0 vdd
port 180 nsew power bidirectional
flabel metal4 s 35168 3076 35488 44748 0 FreeSans 1280 90 0 0 vdd
port 180 nsew power bidirectional
flabel metal4 s 19808 3076 20128 44748 0 FreeSans 1280 90 0 0 vss
port 181 nsew ground bidirectional
rlabel metal1 23968 44688 23968 44688 0 vdd
rlabel metal1 23968 43904 23968 43904 0 vss
rlabel metal2 13496 17304 13496 17304 0 _000_
rlabel metal2 12152 17976 12152 17976 0 _001_
rlabel metal2 11480 16688 11480 16688 0 _002_
rlabel metal2 8344 16240 8344 16240 0 _003_
rlabel metal2 8232 17192 8232 17192 0 _004_
rlabel metal2 6216 14056 6216 14056 0 _005_
rlabel metal2 2016 15512 2016 15512 0 _006_
rlabel metal2 4536 11200 4536 11200 0 _007_
rlabel metal2 11480 19040 11480 19040 0 _008_
rlabel metal2 8680 20832 8680 20832 0 _009_
rlabel metal2 6104 21896 6104 21896 0 _010_
rlabel metal2 5992 18872 5992 18872 0 _011_
rlabel metal2 2184 17752 2184 17752 0 _012_
rlabel metal2 10248 19992 10248 19992 0 _013_
rlabel metal3 3640 13944 3640 13944 0 _014_
rlabel metal2 2296 14168 2296 14168 0 _015_
rlabel metal2 5544 23576 5544 23576 0 _016_
rlabel metal2 3640 24080 3640 24080 0 _017_
rlabel metal2 2464 20216 2464 20216 0 _018_
rlabel metal2 2184 20552 2184 20552 0 _019_
rlabel metal2 13944 22456 13944 22456 0 _020_
rlabel metal2 15064 22008 15064 22008 0 _021_
rlabel metal2 11928 21896 11928 21896 0 _022_
rlabel metal2 10136 20888 10136 20888 0 _023_
rlabel metal2 16128 24920 16128 24920 0 _024_
rlabel metal2 14952 25480 14952 25480 0 _025_
rlabel metal2 12488 26068 12488 26068 0 _026_
rlabel metal2 12600 25144 12600 25144 0 _027_
rlabel metal2 12264 24472 12264 24472 0 _028_
rlabel metal2 11256 26600 11256 26600 0 _029_
rlabel metal3 9128 26488 9128 26488 0 _030_
rlabel metal2 4760 25312 4760 25312 0 _031_
rlabel metal2 8680 29792 8680 29792 0 _032_
rlabel metal2 7560 29176 7560 29176 0 _033_
rlabel metal2 4312 28336 4312 28336 0 _034_
rlabel metal2 5600 27160 5600 27160 0 _035_
rlabel metal2 2072 30744 2072 30744 0 _036_
rlabel metal2 2240 34328 2240 34328 0 _037_
rlabel metal3 5320 28728 5320 28728 0 _038_
rlabel metal2 2688 27720 2688 27720 0 _039_
rlabel metal2 16408 30464 16408 30464 0 _040_
rlabel metal2 16520 31920 16520 31920 0 _041_
rlabel metal2 17416 30072 17416 30072 0 _042_
rlabel metal2 16520 34328 16520 34328 0 _043_
rlabel metal3 13328 30184 13328 30184 0 _044_
rlabel metal3 12040 29624 12040 29624 0 _045_
rlabel metal2 10808 31864 10808 31864 0 _046_
rlabel metal2 11256 28504 11256 28504 0 _047_
rlabel metal2 14952 30688 14952 30688 0 _048_
rlabel metal2 12488 30016 12488 30016 0 _049_
rlabel metal2 26040 29792 26040 29792 0 _050_
rlabel metal2 24248 31136 24248 31136 0 _051_
rlabel metal2 25256 30184 25256 30184 0 _052_
rlabel metal2 23016 32424 23016 32424 0 _053_
rlabel metal2 20440 30856 20440 30856 0 _054_
rlabel metal2 18088 31640 18088 31640 0 _055_
rlabel metal2 24136 27328 24136 27328 0 _056_
rlabel metal2 21560 28392 21560 28392 0 _057_
rlabel metal2 22456 26684 22456 26684 0 _058_
rlabel metal2 20328 28336 20328 28336 0 _059_
rlabel metal2 18872 26432 18872 26432 0 _060_
rlabel metal2 18088 27440 18088 27440 0 _061_
rlabel metal2 16520 26628 16520 26628 0 _062_
rlabel metal2 19096 29176 19096 29176 0 _063_
rlabel metal2 19880 17920 19880 17920 0 _064_
rlabel metal2 17752 17024 17752 17024 0 _065_
rlabel metal2 17864 15904 17864 15904 0 _066_
rlabel metal3 17080 18424 17080 18424 0 _067_
rlabel metal2 19208 19152 19208 19152 0 _068_
rlabel metal2 19880 19152 19880 19152 0 _069_
rlabel metal2 23128 19488 23128 19488 0 _070_
rlabel metal2 24024 19320 24024 19320 0 _071_
rlabel metal2 27888 17528 27888 17528 0 _072_
rlabel metal2 25928 16240 25928 16240 0 _073_
rlabel metal2 26712 15960 26712 15960 0 _074_
rlabel metal2 24696 15512 24696 15512 0 _075_
rlabel metal2 24248 13832 24248 13832 0 _076_
rlabel metal2 22232 16744 22232 16744 0 _077_
rlabel metal2 23240 16912 23240 16912 0 _078_
rlabel metal2 21672 18144 21672 18144 0 _079_
rlabel metal2 36288 13048 36288 13048 0 _080_
rlabel metal2 36232 12040 36232 12040 0 _081_
rlabel metal2 35560 13048 35560 13048 0 _082_
rlabel metal2 35112 13720 35112 13720 0 _083_
rlabel metal2 33768 14056 33768 14056 0 _084_
rlabel metal2 33096 14224 33096 14224 0 _085_
rlabel metal3 30912 15512 30912 15512 0 _086_
rlabel metal2 31864 16128 31864 16128 0 _087_
rlabel metal2 34888 14952 34888 14952 0 _088_
rlabel metal2 33656 17472 33656 17472 0 _089_
rlabel metal2 44856 17920 44856 17920 0 _090_
rlabel metal2 43624 18256 43624 18256 0 _091_
rlabel metal3 43680 18536 43680 18536 0 _092_
rlabel metal2 41048 15736 41048 15736 0 _093_
rlabel metal2 40040 16016 40040 16016 0 _094_
rlabel metal2 38584 14560 38584 14560 0 _095_
rlabel metal3 44352 22120 44352 22120 0 _096_
rlabel metal2 43848 20944 43848 20944 0 _097_
rlabel metal2 43512 20552 43512 20552 0 _098_
rlabel metal2 40376 21952 40376 21952 0 _099_
rlabel metal2 39928 22904 39928 22904 0 _100_
rlabel metal2 37128 23520 37128 23520 0 _101_
rlabel metal2 35896 20888 35896 20888 0 _102_
rlabel metal2 35784 19936 35784 19936 0 _103_
rlabel metal2 38024 27552 38024 27552 0 _104_
rlabel metal2 35784 26600 35784 26600 0 _105_
rlabel metal2 37240 25816 37240 25816 0 _106_
rlabel metal2 37576 25536 37576 25536 0 _107_
rlabel metal2 36008 22736 36008 22736 0 _108_
rlabel metal2 34776 24304 34776 24304 0 _109_
rlabel metal2 45248 23352 45248 23352 0 _110_
rlabel metal2 45752 25144 45752 25144 0 _111_
rlabel metal2 45864 30688 45864 30688 0 _112_
rlabel metal2 43848 31360 43848 31360 0 _113_
rlabel metal2 45752 30464 45752 30464 0 _114_
rlabel metal2 44688 30744 44688 30744 0 _115_
rlabel metal2 45024 31304 45024 31304 0 _116_
rlabel metal2 41608 29848 41608 29848 0 _117_
rlabel metal2 42056 31584 42056 31584 0 _118_
rlabel metal2 40264 31192 40264 31192 0 _119_
rlabel metal2 33544 29736 33544 29736 0 _120_
rlabel metal2 35896 31360 35896 31360 0 _121_
rlabel metal2 32200 31192 32200 31192 0 _122_
rlabel metal2 30968 30128 30968 30128 0 _123_
rlabel metal3 29680 32424 29680 32424 0 _124_
rlabel metal3 30464 32984 30464 32984 0 _125_
rlabel metal2 29736 32704 29736 32704 0 _126_
rlabel metal2 28672 31192 28672 31192 0 _127_
rlabel metal3 30800 29288 30800 29288 0 _128_
rlabel metal3 28616 28056 28616 28056 0 _129_
rlabel metal2 25816 24920 25816 24920 0 _130_
rlabel metal2 28280 26040 28280 26040 0 _131_
rlabel metal2 24024 25536 24024 25536 0 _132_
rlabel metal2 22568 23520 22568 23520 0 _133_
rlabel metal2 20440 24472 20440 24472 0 _134_
rlabel metal2 21336 23744 21336 23744 0 _135_
rlabel metal2 21224 22400 21224 22400 0 _136_
rlabel metal2 24360 21896 24360 21896 0 _137_
rlabel metal2 21448 19936 21448 19936 0 _138_
rlabel metal2 18032 20552 18032 20552 0 _139_
rlabel metal2 29848 21952 29848 21952 0 _140_
rlabel metal2 30072 23800 30072 23800 0 _141_
rlabel metal2 28616 24024 28616 24024 0 _142_
rlabel metal2 27272 24696 27272 24696 0 _143_
rlabel metal3 34216 18984 34216 18984 0 _144_
rlabel metal2 34440 18312 34440 18312 0 _145_
rlabel metal2 28056 20944 28056 20944 0 _146_
rlabel metal2 26936 19264 26936 19264 0 _147_
rlabel metal2 28504 20888 28504 20888 0 _148_
rlabel metal3 29344 19320 29344 19320 0 _149_
rlabel metal3 41888 19320 41888 19320 0 _150_
rlabel metal2 40040 21504 40040 21504 0 _151_
rlabel metal2 43624 27636 43624 27636 0 _152_
rlabel metal2 44576 24920 44576 24920 0 _153_
rlabel metal2 44856 26208 44856 26208 0 _154_
rlabel metal2 43848 26040 43848 26040 0 _155_
rlabel metal2 41496 25312 41496 25312 0 _156_
rlabel metal2 43960 29400 43960 29400 0 _157_
rlabel metal2 39928 29624 39928 29624 0 _158_
rlabel metal2 40936 28168 40936 28168 0 _159_
rlabel metal2 31080 24248 31080 24248 0 _160_
rlabel metal2 31864 27328 31864 27328 0 _161_
rlabel metal2 3192 13944 3192 13944 0 _162_
rlabel metal2 5992 23464 5992 23464 0 _163_
rlabel metal2 11424 21672 11424 21672 0 _164_
rlabel metal2 1960 29400 1960 29400 0 _165_
rlabel metal2 17640 28728 17640 28728 0 _166_
rlabel metal2 21672 28784 21672 28784 0 _167_
rlabel metal3 17416 26152 17416 26152 0 _168_
rlabel metal2 27608 16520 27608 16520 0 _169_
rlabel metal2 34104 18368 34104 18368 0 _170_
rlabel metal2 38360 19712 38360 19712 0 _171_
rlabel metal2 37800 25312 37800 25312 0 _172_
rlabel metal3 45304 29288 45304 29288 0 _173_
rlabel metal2 31584 28056 31584 28056 0 _174_
rlabel metal3 29120 25368 29120 25368 0 _175_
rlabel metal2 31080 23072 31080 23072 0 _176_
rlabel metal2 44184 30184 44184 30184 0 _177_
rlabel metal2 3528 20440 3528 20440 0 ccff_head
rlabel metal2 45752 26908 45752 26908 0 ccff_tail
rlabel metal2 42168 3864 42168 3864 0 chanx_left_in[0]
rlabel metal2 27664 4200 27664 4200 0 chanx_left_in[10]
rlabel metal2 6832 3416 6832 3416 0 chanx_left_in[12]
rlabel metal2 13552 4200 13552 4200 0 chanx_left_in[13]
rlabel metal2 17416 4256 17416 4256 0 chanx_left_in[14]
rlabel metal3 24752 43624 24752 43624 0 chanx_left_in[16]
rlabel metal2 13496 45850 13496 45850 0 chanx_left_in[17]
rlabel metal2 11536 3416 11536 3416 0 chanx_left_in[18]
rlabel metal2 18872 2058 18872 2058 0 chanx_left_in[1]
rlabel metal2 14168 2478 14168 2478 0 chanx_left_in[2]
rlabel metal2 27608 44576 27608 44576 0 chanx_left_in[4]
rlabel metal2 10864 3416 10864 3416 0 chanx_left_in[5]
rlabel metal2 33432 44800 33432 44800 0 chanx_left_in[6]
rlabel metal2 30240 43736 30240 43736 0 chanx_left_in[8]
rlabel metal2 22904 45486 22904 45486 0 chanx_left_in[9]
rlabel metal2 20888 1246 20888 1246 0 chanx_left_out[10]
rlabel metal2 17528 44688 17528 44688 0 chanx_left_out[11]
rlabel metal2 7448 1414 7448 1414 0 chanx_left_out[13]
rlabel metal3 46522 44408 46522 44408 0 chanx_left_out[14]
rlabel metal2 41048 1246 41048 1246 0 chanx_left_out[15]
rlabel metal2 39032 2198 39032 2198 0 chanx_left_out[17]
rlabel metal2 32816 3640 32816 3640 0 chanx_left_out[18]
rlabel metal2 21672 3304 21672 3304 0 chanx_left_out[19]
rlabel metal2 46088 43232 46088 43232 0 chanx_left_out[1]
rlabel metal2 27272 3752 27272 3752 0 chanx_left_out[2]
rlabel metal3 30072 3640 30072 3640 0 chanx_left_out[3]
rlabel metal2 21000 44632 21000 44632 0 chanx_left_out[5]
rlabel metal3 36680 3640 36680 3640 0 chanx_left_out[6]
rlabel metal2 24248 1246 24248 1246 0 chanx_left_out[7]
rlabel metal2 26544 45528 26544 45528 0 chanx_left_out[9]
rlabel metal3 46746 41048 46746 41048 0 chanx_right_in[0]
rlabel metal2 19096 45528 19096 45528 0 chanx_right_in[10]
rlabel metal2 24024 3192 24024 3192 0 chanx_right_in[12]
rlabel metal2 46200 43960 46200 43960 0 chanx_right_in[13]
rlabel metal2 39704 2478 39704 2478 0 chanx_right_in[14]
rlabel metal2 37800 3416 37800 3416 0 chanx_right_in[16]
rlabel metal2 31864 3864 31864 3864 0 chanx_right_in[17]
rlabel metal2 23072 3640 23072 3640 0 chanx_right_in[18]
rlabel metal2 25592 2058 25592 2058 0 chanx_right_in[1]
rlabel metal2 31416 4144 31416 4144 0 chanx_right_in[2]
rlabel metal2 20888 45486 20888 45486 0 chanx_right_in[4]
rlabel metal3 33432 3416 33432 3416 0 chanx_right_in[5]
rlabel metal2 9688 3696 9688 3696 0 chanx_right_in[6]
rlabel metal2 25368 44744 25368 44744 0 chanx_right_in[8]
rlabel metal2 19656 4424 19656 4424 0 chanx_right_in[9]
rlabel metal2 23520 44408 23520 44408 0 chanx_right_out[10]
rlabel metal3 28784 3416 28784 3416 0 chanx_right_out[11]
rlabel metal2 12152 2422 12152 2422 0 chanx_right_out[13]
rlabel metal2 14840 2478 14840 2478 0 chanx_right_out[14]
rlabel metal2 17696 3304 17696 3304 0 chanx_right_out[15]
rlabel metal3 25256 44520 25256 44520 0 chanx_right_out[17]
rlabel metal2 14952 44632 14952 44632 0 chanx_right_out[18]
rlabel metal2 8792 854 8792 854 0 chanx_right_out[19]
rlabel metal2 24920 2058 24920 2058 0 chanx_right_out[1]
rlabel metal2 20216 2058 20216 2058 0 chanx_right_out[2]
rlabel metal2 15568 3304 15568 3304 0 chanx_right_out[3]
rlabel metal2 30408 44464 30408 44464 0 chanx_right_out[5]
rlabel metal2 8120 2030 8120 2030 0 chanx_right_out[6]
rlabel metal2 28840 44856 28840 44856 0 chanx_right_out[7]
rlabel metal2 30968 45906 30968 45906 0 chanx_right_out[9]
rlabel metal2 34552 44688 34552 44688 0 chany_bottom_in[0]
rlabel metal2 16184 2058 16184 2058 0 chany_bottom_in[10]
rlabel metal2 22232 2058 22232 2058 0 chany_bottom_in[12]
rlabel metal3 35784 4200 35784 4200 0 chany_bottom_in[13]
rlabel metal2 35112 43624 35112 43624 0 chany_bottom_in[14]
rlabel metal2 41160 3696 41160 3696 0 chany_bottom_in[16]
rlabel metal2 46200 20104 46200 20104 0 chany_bottom_in[17]
rlabel metal3 46074 10808 46074 10808 0 chany_bottom_in[18]
rlabel metal2 35896 3080 35896 3080 0 chany_bottom_in[1]
rlabel metal3 34328 3528 34328 3528 0 chany_bottom_in[2]
rlabel metal2 30744 4256 30744 4256 0 chany_bottom_in[4]
rlabel metal2 46200 5320 46200 5320 0 chany_bottom_in[5]
rlabel metal2 41776 45528 41776 45528 0 chany_bottom_in[6]
rlabel metal3 27440 3528 27440 3528 0 chany_bottom_in[8]
rlabel metal3 38864 3416 38864 3416 0 chany_bottom_in[9]
rlabel metal2 12824 2030 12824 2030 0 chany_bottom_out[10]
rlabel metal2 40320 44408 40320 44408 0 chany_bottom_out[11]
rlabel metal2 28392 44296 28392 44296 0 chany_bottom_out[13]
rlabel metal2 37576 4200 37576 4200 0 chany_bottom_out[14]
rlabel metal3 1414 7448 1414 7448 0 chany_bottom_out[15]
rlabel metal3 46634 14168 46634 14168 0 chany_bottom_out[17]
rlabel metal3 46410 15512 46410 15512 0 chany_bottom_out[18]
rlabel metal2 19544 45850 19544 45850 0 chany_bottom_out[19]
rlabel metal2 8120 45906 8120 45906 0 chany_bottom_out[1]
rlabel metal2 22232 45486 22232 45486 0 chany_bottom_out[2]
rlabel metal2 46088 18256 46088 18256 0 chany_bottom_out[3]
rlabel metal2 43624 13272 43624 13272 0 chany_bottom_out[5]
rlabel metal2 44072 44464 44072 44464 0 chany_bottom_out[6]
rlabel metal3 1358 5432 1358 5432 0 chany_bottom_out[7]
rlabel metal2 41944 44632 41944 44632 0 chany_bottom_out[9]
rlabel metal2 7448 45850 7448 45850 0 chany_top_in[0]
rlabel metal2 38808 44744 38808 44744 0 chany_top_in[10]
rlabel metal2 31640 45458 31640 45458 0 chany_top_in[12]
rlabel metal2 43960 9352 43960 9352 0 chany_top_in[13]
rlabel metal2 1736 4928 1736 4928 0 chany_top_in[14]
rlabel metal3 43736 12936 43736 12936 0 chany_top_in[16]
rlabel metal2 46088 4816 46088 4816 0 chany_top_in[17]
rlabel metal2 18312 43512 18312 43512 0 chany_top_in[18]
rlabel metal3 21224 43512 21224 43512 0 chany_top_in[1]
rlabel metal2 46088 10360 46088 10360 0 chany_top_in[2]
rlabel metal2 44296 7896 44296 7896 0 chany_top_in[4]
rlabel metal2 38136 44576 38136 44576 0 chany_top_in[5]
rlabel metal3 1246 3416 1246 3416 0 chany_top_in[6]
rlabel metal2 39816 45528 39816 45528 0 chany_top_in[8]
rlabel metal2 1736 4200 1736 4200 0 chany_top_in[9]
rlabel metal2 45752 7056 45752 7056 0 chany_top_out[10]
rlabel metal3 1414 6104 1414 6104 0 chany_top_out[11]
rlabel metal3 1358 6776 1358 6776 0 chany_top_out[13]
rlabel metal2 45416 9968 45416 9968 0 chany_top_out[14]
rlabel metal2 37128 44464 37128 44464 0 chany_top_out[15]
rlabel metal2 45640 5936 45640 5936 0 chany_top_out[17]
rlabel metal3 46690 17528 46690 17528 0 chany_top_out[18]
rlabel metal3 46410 16184 46410 16184 0 chany_top_out[19]
rlabel metal2 38024 45528 38024 45528 0 chany_top_out[1]
rlabel metal2 45752 13216 45752 13216 0 chany_top_out[2]
rlabel metal2 46088 7840 46088 7840 0 chany_top_out[3]
rlabel metal3 46466 11480 46466 11480 0 chany_top_out[5]
rlabel metal3 46690 16856 46690 16856 0 chany_top_out[6]
rlabel metal2 41272 45528 41272 45528 0 chany_top_out[7]
rlabel metal3 46690 18872 46690 18872 0 chany_top_out[9]
rlabel metal2 27048 28952 27048 28952 0 clknet_0_prog_clk
rlabel metal2 1904 13720 1904 13720 0 clknet_4_0_0_prog_clk
rlabel metal2 38584 18816 38584 18816 0 clknet_4_10_0_prog_clk
rlabel metal2 37128 21560 37128 21560 0 clknet_4_11_0_prog_clk
rlabel metal2 31416 25816 31416 25816 0 clknet_4_12_0_prog_clk
rlabel metal2 28168 29456 28168 29456 0 clknet_4_13_0_prog_clk
rlabel metal2 32928 24696 32928 24696 0 clknet_4_14_0_prog_clk
rlabel metal2 44408 30464 44408 30464 0 clknet_4_15_0_prog_clk
rlabel metal2 5544 22736 5544 22736 0 clknet_4_1_0_prog_clk
rlabel metal2 14952 16856 14952 16856 0 clknet_4_2_0_prog_clk
rlabel metal2 13216 20776 13216 20776 0 clknet_4_3_0_prog_clk
rlabel metal3 6832 26264 6832 26264 0 clknet_4_4_0_prog_clk
rlabel metal2 2296 30632 2296 30632 0 clknet_4_5_0_prog_clk
rlabel metal2 19992 24304 19992 24304 0 clknet_4_6_0_prog_clk
rlabel via2 17192 30184 17192 30184 0 clknet_4_7_0_prog_clk
rlabel metal2 29344 21448 29344 21448 0 clknet_4_8_0_prog_clk
rlabel metal2 26936 22400 26936 22400 0 clknet_4_9_0_prog_clk
rlabel metal2 20888 17976 20888 17976 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 27272 13944 27272 13944 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal3 21448 18984 21448 18984 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 17080 17836 17080 17836 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 15400 17080 15400 17080 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 15736 16856 15736 16856 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal2 16744 13384 16744 13384 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal2 15064 15344 15064 15344 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal2 20664 15624 20664 15624 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal2 29400 11312 29400 11312 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal2 34440 12320 34440 12320 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal2 34328 13944 34328 13944 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 33992 12320 33992 12320 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal3 34608 9128 34608 9128 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal3 37632 10696 37632 10696 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal3 34216 10696 34216 10696 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal2 42168 9856 42168 9856 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal2 39368 10696 39368 10696 0 mem_bottom_track_17.DFFR_7_.Q
rlabel metal2 41272 8260 41272 8260 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 42392 7980 42392 7980 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal2 46088 8904 46088 8904 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal2 41048 10976 41048 10976 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal2 42840 7476 42840 7476 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal3 42336 15400 42336 15400 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal2 36456 14504 36456 14504 0 mem_bottom_track_25.DFFR_6_.Q
rlabel metal2 37352 14168 37352 14168 0 mem_bottom_track_25.DFFR_7_.Q
rlabel metal3 41664 12264 41664 12264 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal3 41720 20104 41720 20104 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal2 28168 20328 28168 20328 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal2 29008 20776 29008 20776 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal2 26152 16800 26152 16800 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal2 29064 17192 29064 17192 0 mem_bottom_track_33.DFFR_5_.Q
rlabel metal2 32760 19824 32760 19824 0 mem_bottom_track_33.DFFR_6_.Q
rlabel metal2 35672 14560 35672 14560 0 mem_bottom_track_33.DFFR_7_.Q
rlabel metal3 23296 16632 23296 16632 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal3 23408 15064 23408 15064 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal2 21224 15484 21224 15484 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal2 26320 16632 26320 16632 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal2 27944 12936 27944 12936 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal3 28952 12264 28952 12264 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal2 27608 12824 27608 12824 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal3 37016 20552 37016 20552 0 mem_left_track_1.DFFR_0_.Q
rlabel metal2 36680 20748 36680 20748 0 mem_left_track_1.DFFR_1_.Q
rlabel metal2 37912 22232 37912 22232 0 mem_left_track_1.DFFR_2_.Q
rlabel metal3 41496 18200 41496 18200 0 mem_left_track_1.DFFR_3_.Q
rlabel metal2 43960 10976 43960 10976 0 mem_left_track_1.DFFR_4_.Q
rlabel metal2 43344 11256 43344 11256 0 mem_left_track_1.DFFR_5_.Q
rlabel metal2 46088 9520 46088 9520 0 mem_left_track_1.DFFR_6_.Q
rlabel metal2 44184 22120 44184 22120 0 mem_left_track_1.DFFR_7_.Q
rlabel metal2 38808 30072 38808 30072 0 mem_left_track_17.DFFR_0_.D
rlabel metal3 41048 32760 41048 32760 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 42280 37800 42280 37800 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 40824 30408 40824 30408 0 mem_left_track_17.DFFR_2_.Q
rlabel metal2 45528 35280 45528 35280 0 mem_left_track_17.DFFR_3_.Q
rlabel metal2 45192 33264 45192 33264 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 44408 35280 44408 35280 0 mem_left_track_17.DFFR_5_.Q
rlabel metal2 44408 42056 44408 42056 0 mem_left_track_17.DFFR_6_.Q
rlabel metal2 30072 31472 30072 31472 0 mem_left_track_17.DFFR_7_.Q
rlabel metal3 30856 31080 30856 31080 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 30352 32760 30352 32760 0 mem_left_track_25.DFFR_1_.Q
rlabel metal3 29680 33096 29680 33096 0 mem_left_track_25.DFFR_2_.Q
rlabel metal3 29960 33208 29960 33208 0 mem_left_track_25.DFFR_3_.Q
rlabel metal2 31528 30408 31528 30408 0 mem_left_track_25.DFFR_4_.Q
rlabel metal2 33096 34216 33096 34216 0 mem_left_track_25.DFFR_5_.Q
rlabel metal3 37856 33544 37856 33544 0 mem_left_track_25.DFFR_6_.Q
rlabel metal2 32872 30464 32872 30464 0 mem_left_track_25.DFFR_7_.Q
rlabel metal2 36512 28840 36512 28840 0 mem_left_track_33.DFFR_0_.Q
rlabel metal2 40600 29736 40600 29736 0 mem_left_track_33.DFFR_1_.Q
rlabel metal2 40656 27272 40656 27272 0 mem_left_track_33.DFFR_2_.Q
rlabel metal2 45416 14392 45416 14392 0 mem_left_track_33.DFFR_3_.Q
rlabel metal2 43288 19656 43288 19656 0 mem_left_track_33.DFFR_4_.Q
rlabel metal2 44352 27272 44352 27272 0 mem_left_track_33.DFFR_5_.Q
rlabel metal2 45136 28168 45136 28168 0 mem_left_track_33.DFFR_6_.Q
rlabel metal3 45584 27048 45584 27048 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 39480 16072 39480 16072 0 mem_left_track_9.DFFR_1_.Q
rlabel metal2 35448 25704 35448 25704 0 mem_left_track_9.DFFR_2_.Q
rlabel metal3 37352 22232 37352 22232 0 mem_left_track_9.DFFR_3_.Q
rlabel metal2 36848 26488 36848 26488 0 mem_left_track_9.DFFR_4_.Q
rlabel metal3 33432 32648 33432 32648 0 mem_left_track_9.DFFR_5_.Q
rlabel metal2 37408 28056 37408 28056 0 mem_left_track_9.DFFR_6_.Q
rlabel metal2 29064 30128 29064 30128 0 mem_right_track_0.DFFR_0_.D
rlabel metal3 2016 30408 2016 30408 0 mem_right_track_0.DFFR_0_.Q
rlabel metal2 5768 32200 5768 32200 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 1736 34552 1736 34552 0 mem_right_track_0.DFFR_2_.Q
rlabel metal2 5264 31864 5264 31864 0 mem_right_track_0.DFFR_3_.Q
rlabel metal2 6104 33488 6104 33488 0 mem_right_track_0.DFFR_4_.Q
rlabel metal2 2296 28784 2296 28784 0 mem_right_track_0.DFFR_5_.Q
rlabel metal2 3080 29848 3080 29848 0 mem_right_track_0.DFFR_6_.Q
rlabel metal2 9296 30184 9296 30184 0 mem_right_track_0.DFFR_7_.Q
rlabel metal2 15624 31976 15624 31976 0 mem_right_track_16.DFFR_0_.D
rlabel metal2 17304 32368 17304 32368 0 mem_right_track_16.DFFR_0_.Q
rlabel metal2 20888 31920 20888 31920 0 mem_right_track_16.DFFR_1_.Q
rlabel metal2 21224 34104 21224 34104 0 mem_right_track_16.DFFR_2_.Q
rlabel metal2 24360 33768 24360 33768 0 mem_right_track_16.DFFR_3_.Q
rlabel metal2 27272 33656 27272 33656 0 mem_right_track_16.DFFR_4_.Q
rlabel metal3 18984 29960 18984 29960 0 mem_right_track_16.DFFR_5_.Q
rlabel metal2 13048 30464 13048 30464 0 mem_right_track_16.DFFR_6_.Q
rlabel metal2 15736 32704 15736 32704 0 mem_right_track_16.DFFR_7_.Q
rlabel metal2 16968 30632 16968 30632 0 mem_right_track_24.DFFR_0_.Q
rlabel metal2 16968 28728 16968 28728 0 mem_right_track_24.DFFR_1_.Q
rlabel metal2 18816 28840 18816 28840 0 mem_right_track_24.DFFR_2_.Q
rlabel metal2 16296 28504 16296 28504 0 mem_right_track_24.DFFR_3_.Q
rlabel metal2 22064 29624 22064 29624 0 mem_right_track_24.DFFR_4_.Q
rlabel metal3 24472 33208 24472 33208 0 mem_right_track_24.DFFR_5_.Q
rlabel metal2 20776 28224 20776 28224 0 mem_right_track_24.DFFR_6_.Q
rlabel metal2 24920 28672 24920 28672 0 mem_right_track_24.DFFR_7_.Q
rlabel metal2 28056 24864 28056 24864 0 mem_right_track_32.DFFR_0_.Q
rlabel metal2 29400 25928 29400 25928 0 mem_right_track_32.DFFR_1_.Q
rlabel metal2 30632 23464 30632 23464 0 mem_right_track_32.DFFR_2_.Q
rlabel metal3 28224 21896 28224 21896 0 mem_right_track_32.DFFR_3_.Q
rlabel metal2 19768 14952 19768 14952 0 mem_right_track_32.DFFR_4_.Q
rlabel metal2 18872 17808 18872 17808 0 mem_right_track_32.DFFR_5_.Q
rlabel metal3 31920 22008 31920 22008 0 mem_right_track_32.DFFR_6_.Q
rlabel metal2 11816 29792 11816 29792 0 mem_right_track_8.DFFR_0_.Q
rlabel metal3 8232 32648 8232 32648 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 13160 29792 13160 29792 0 mem_right_track_8.DFFR_2_.Q
rlabel metal2 12936 31864 12936 31864 0 mem_right_track_8.DFFR_3_.Q
rlabel metal2 17080 35728 17080 35728 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 15848 35336 15848 35336 0 mem_right_track_8.DFFR_5_.Q
rlabel metal2 17136 31976 17136 31976 0 mem_right_track_8.DFFR_6_.Q
rlabel metal2 5320 10024 5320 10024 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 11816 12040 11816 12040 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 6776 11648 6776 11648 0 mem_top_track_0.DFFR_2_.Q
rlabel metal2 7784 12320 7784 12320 0 mem_top_track_0.DFFR_3_.Q
rlabel metal2 7000 15232 7000 15232 0 mem_top_track_0.DFFR_4_.Q
rlabel metal2 12544 12264 12544 12264 0 mem_top_track_0.DFFR_5_.Q
rlabel metal2 13608 14728 13608 14728 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 4984 15624 4984 15624 0 mem_top_track_0.DFFR_7_.Q
rlabel metal2 11928 16296 11928 16296 0 mem_top_track_16.DFFR_0_.D
rlabel metal3 6216 20664 6216 20664 0 mem_top_track_16.DFFR_0_.Q
rlabel metal3 8064 22232 8064 22232 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 14728 18200 14728 18200 0 mem_top_track_16.DFFR_2_.Q
rlabel metal3 12432 22904 12432 22904 0 mem_top_track_16.DFFR_3_.Q
rlabel metal3 1960 12824 1960 12824 0 mem_top_track_16.DFFR_4_.Q
rlabel metal2 2744 17752 2744 17752 0 mem_top_track_16.DFFR_5_.Q
rlabel metal2 3416 16968 3416 16968 0 mem_top_track_16.DFFR_6_.Q
rlabel metal2 2856 21000 2856 21000 0 mem_top_track_16.DFFR_7_.Q
rlabel metal2 3976 25704 3976 25704 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 9128 26684 9128 26684 0 mem_top_track_24.DFFR_1_.Q
rlabel metal3 7392 26936 7392 26936 0 mem_top_track_24.DFFR_2_.Q
rlabel metal2 6104 19376 6104 19376 0 mem_top_track_24.DFFR_3_.Q
rlabel metal2 13160 24136 13160 24136 0 mem_top_track_24.DFFR_4_.Q
rlabel metal2 13048 26040 13048 26040 0 mem_top_track_24.DFFR_5_.Q
rlabel metal2 16520 20440 16520 20440 0 mem_top_track_24.DFFR_6_.Q
rlabel metal2 17416 15400 17416 15400 0 mem_top_track_24.DFFR_7_.Q
rlabel metal2 6664 23744 6664 23744 0 mem_top_track_32.DFFR_0_.Q
rlabel metal3 18200 24920 18200 24920 0 mem_top_track_32.DFFR_1_.Q
rlabel metal2 14056 23856 14056 23856 0 mem_top_track_32.DFFR_2_.Q
rlabel metal3 23464 24920 23464 24920 0 mem_top_track_32.DFFR_3_.Q
rlabel metal3 30016 23800 30016 23800 0 mem_top_track_32.DFFR_4_.Q
rlabel metal3 23856 27272 23856 27272 0 mem_top_track_32.DFFR_5_.Q
rlabel metal2 30632 28896 30632 28896 0 mem_top_track_32.DFFR_6_.Q
rlabel metal3 2016 11256 2016 11256 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 5656 13272 5656 13272 0 mem_top_track_8.DFFR_1_.Q
rlabel metal2 8120 13832 8120 13832 0 mem_top_track_8.DFFR_2_.Q
rlabel metal2 6552 13776 6552 13776 0 mem_top_track_8.DFFR_3_.Q
rlabel metal2 3080 17864 3080 17864 0 mem_top_track_8.DFFR_4_.Q
rlabel metal2 7784 18984 7784 18984 0 mem_top_track_8.DFFR_5_.Q
rlabel metal3 10248 18648 10248 18648 0 mem_top_track_8.DFFR_6_.Q
rlabel metal2 2632 10584 2632 10584 0 net1
rlabel metal2 19432 4816 19432 4816 0 net10
rlabel metal2 28504 8848 28504 8848 0 net100
rlabel metal2 20216 43988 20216 43988 0 net101
rlabel metal2 7784 43344 7784 43344 0 net102
rlabel metal2 21896 42448 21896 42448 0 net103
rlabel metal2 31752 12824 31752 12824 0 net104
rlabel metal2 28616 11312 28616 11312 0 net105
rlabel metal3 41328 44296 41328 44296 0 net106
rlabel metal3 5684 5880 5684 5880 0 net107
rlabel metal2 41384 43876 41384 43876 0 net108
rlabel metal2 38584 5712 38584 5712 0 net109
rlabel metal2 14784 4536 14784 4536 0 net11
rlabel metal2 16632 5824 16632 5824 0 net110
rlabel metal2 2968 7392 2968 7392 0 net111
rlabel metal2 34216 5824 34216 5824 0 net112
rlabel metal2 37576 44296 37576 44296 0 net113
rlabel metal2 40376 5040 40376 5040 0 net114
rlabel metal2 44296 5880 44296 5880 0 net115
rlabel metal2 46256 4536 46256 4536 0 net116
rlabel metal2 38584 43064 38584 43064 0 net117
rlabel metal3 35280 9800 35280 9800 0 net118
rlabel metal2 33432 4760 33432 4760 0 net119
rlabel metal2 27384 43876 27384 43876 0 net12
rlabel metal2 30296 6440 30296 6440 0 net120
rlabel metal2 44744 6468 44744 6468 0 net121
rlabel metal3 40600 42616 40600 42616 0 net122
rlabel metal2 27048 5320 27048 5320 0 net123
rlabel metal2 43960 2856 43960 2856 0 net124
rlabel metal2 43064 3360 43064 3360 0 net125
rlabel metal2 36008 44912 36008 44912 0 net126
rlabel metal2 44408 2688 44408 2688 0 net127
rlabel metal2 17752 44632 17752 44632 0 net128
rlabel metal2 43848 3976 43848 3976 0 net129
rlabel metal2 11256 3472 11256 3472 0 net13
rlabel metal3 45486 4760 45486 4760 0 net130
rlabel metal2 46200 39872 46200 39872 0 net131
rlabel metal2 44856 2016 44856 2016 0 net132
rlabel metal2 35000 2030 35000 2030 0 net133
rlabel metal2 43624 4256 43624 4256 0 net134
rlabel metal2 30072 44296 30072 44296 0 net135
rlabel metal3 1582 2744 1582 2744 0 net136
rlabel metal2 29064 4424 29064 4424 0 net137
rlabel metal2 46088 41496 46088 41496 0 net138
rlabel metal3 15400 44184 15400 44184 0 net139
rlabel metal2 28504 42504 28504 42504 0 net14
rlabel metal2 18200 2058 18200 2058 0 net140
rlabel metal3 1246 42392 1246 42392 0 net141
rlabel metal2 45304 3024 45304 3024 0 net142
rlabel metal2 10136 2590 10136 2590 0 net143
rlabel metal3 38136 30296 38136 30296 0 net144
rlabel metal2 34104 33992 34104 33992 0 net145
rlabel metal2 13944 34160 13944 34160 0 net146
rlabel metal2 3864 21392 3864 21392 0 net147
rlabel metal2 13944 19320 13944 19320 0 net148
rlabel metal3 34944 29848 34944 29848 0 net149
rlabel metal2 30296 42784 30296 42784 0 net15
rlabel metal3 18704 17192 18704 17192 0 net150
rlabel metal2 14000 18424 14000 18424 0 net151
rlabel metal2 41384 30268 41384 30268 0 net152
rlabel metal2 3528 29344 3528 29344 0 net153
rlabel metal2 19600 16744 19600 16744 0 net154
rlabel metal3 35616 28728 35616 28728 0 net155
rlabel metal2 29848 30744 29848 30744 0 net156
rlabel metal2 2744 31416 2744 31416 0 net157
rlabel metal2 32200 22680 32200 22680 0 net158
rlabel metal2 23688 28560 23688 28560 0 net159
rlabel metal2 23352 43176 23352 43176 0 net16
rlabel metal2 33656 18088 33656 18088 0 net160
rlabel metal3 28616 21728 28616 21728 0 net161
rlabel metal2 33544 15624 33544 15624 0 net162
rlabel metal3 18424 24024 18424 24024 0 net163
rlabel metal2 25144 31024 25144 31024 0 net164
rlabel metal2 23912 13832 23912 13832 0 net165
rlabel metal2 29848 18984 29848 18984 0 net166
rlabel metal3 22232 15960 22232 15960 0 net167
rlabel metal2 27608 25144 27608 25144 0 net168
rlabel metal2 21896 30520 21896 30520 0 net169
rlabel metal3 45528 41048 45528 41048 0 net17
rlabel metal2 21336 33544 21336 33544 0 net170
rlabel metal2 23968 35560 23968 35560 0 net171
rlabel metal3 25928 26936 25928 26936 0 net172
rlabel metal2 38584 22960 38584 22960 0 net173
rlabel metal2 23912 29232 23912 29232 0 net174
rlabel metal2 33488 22344 33488 22344 0 net175
rlabel metal2 23128 25928 23128 25928 0 net176
rlabel metal3 5432 20552 5432 20552 0 net177
rlabel metal2 4872 17360 4872 17360 0 net178
rlabel metal2 9912 32592 9912 32592 0 net179
rlabel metal2 19096 43176 19096 43176 0 net18
rlabel metal2 37576 21000 37576 21000 0 net180
rlabel metal2 25704 17192 25704 17192 0 net181
rlabel metal2 24472 12488 24472 12488 0 net182
rlabel metal2 42784 12040 42784 12040 0 net183
rlabel metal3 43624 18312 43624 18312 0 net184
rlabel metal2 18760 19544 18760 19544 0 net185
rlabel metal2 42840 14868 42840 14868 0 net186
rlabel metal2 16408 24976 16408 24976 0 net187
rlabel metal2 19488 27048 19488 27048 0 net188
rlabel metal3 29344 30632 29344 30632 0 net189
rlabel metal2 24024 4648 24024 4648 0 net19
rlabel metal2 36680 27720 36680 27720 0 net190
rlabel metal2 5656 15176 5656 15176 0 net191
rlabel metal2 12600 16016 12600 16016 0 net192
rlabel metal2 8008 14392 8008 14392 0 net193
rlabel metal2 41384 34944 41384 34944 0 net194
rlabel metal2 12712 22008 12712 22008 0 net195
rlabel metal2 42112 8680 42112 8680 0 net196
rlabel metal2 37296 16856 37296 16856 0 net197
rlabel metal2 12600 32480 12600 32480 0 net198
rlabel metal2 26152 12040 26152 12040 0 net199
rlabel metal3 31920 4256 31920 4256 0 net2
rlabel metal3 44968 44072 44968 44072 0 net20
rlabel metal2 36008 14392 36008 14392 0 net200
rlabel metal2 41384 26964 41384 26964 0 net201
rlabel metal2 7560 30352 7560 30352 0 net202
rlabel metal2 41328 11480 41328 11480 0 net203
rlabel metal2 17864 31808 17864 31808 0 net204
rlabel metal2 41496 11228 41496 11228 0 net205
rlabel metal2 12376 25928 12376 25928 0 net206
rlabel metal3 41048 12040 41048 12040 0 net207
rlabel metal3 37072 30968 37072 30968 0 net208
rlabel metal2 19656 14784 19656 14784 0 net209
rlabel metal2 39928 4816 39928 4816 0 net21
rlabel metal2 29512 15512 29512 15512 0 net210
rlabel metal2 28168 26320 28168 26320 0 net211
rlabel metal2 6888 21728 6888 21728 0 net212
rlabel metal2 29848 14840 29848 14840 0 net213
rlabel metal3 38360 35560 38360 35560 0 net214
rlabel metal2 9016 18144 9016 18144 0 net215
rlabel metal2 20272 30968 20272 30968 0 net216
rlabel metal2 29176 19712 29176 19712 0 net217
rlabel metal3 16912 16408 16912 16408 0 net218
rlabel metal2 15848 30184 15848 30184 0 net219
rlabel metal2 38136 4256 38136 4256 0 net22
rlabel metal2 8848 28616 8848 28616 0 net220
rlabel metal2 33656 13664 33656 13664 0 net221
rlabel metal2 44968 5824 44968 5824 0 net222
rlabel metal3 44184 21784 44184 21784 0 net223
rlabel metal2 6440 16184 6440 16184 0 net224
rlabel metal3 24304 15848 24304 15848 0 net225
rlabel metal2 32256 28616 32256 28616 0 net226
rlabel metal3 36512 21896 36512 21896 0 net227
rlabel metal2 13944 28504 13944 28504 0 net228
rlabel metal3 41328 33544 41328 33544 0 net229
rlabel metal2 31976 4816 31976 4816 0 net23
rlabel metal2 26040 20720 26040 20720 0 net230
rlabel metal2 29288 13496 29288 13496 0 net231
rlabel metal2 4424 21560 4424 21560 0 net232
rlabel metal2 3752 14504 3752 14504 0 net233
rlabel metal2 2632 13160 2632 13160 0 net234
rlabel metal2 39256 34832 39256 34832 0 net235
rlabel metal2 44296 14364 44296 14364 0 net236
rlabel metal2 32368 35000 32368 35000 0 net237
rlabel metal2 15176 36176 15176 36176 0 net238
rlabel metal2 26376 24360 26376 24360 0 net239
rlabel metal2 22680 4760 22680 4760 0 net24
rlabel metal2 16408 33880 16408 33880 0 net240
rlabel metal3 30184 18536 30184 18536 0 net241
rlabel metal3 29120 30856 29120 30856 0 net242
rlabel metal3 41720 11704 41720 11704 0 net243
rlabel metal2 4088 30184 4088 30184 0 net244
rlabel metal2 2632 15456 2632 15456 0 net245
rlabel metal3 22008 17528 22008 17528 0 net246
rlabel metal2 27160 17416 27160 17416 0 net247
rlabel metal3 40432 38136 40432 38136 0 net248
rlabel metal2 7896 23968 7896 23968 0 net249
rlabel metal2 26712 3696 26712 3696 0 net25
rlabel metal2 28280 14448 28280 14448 0 net250
rlabel metal2 13944 24080 13944 24080 0 net251
rlabel metal2 3640 32984 3640 32984 0 net252
rlabel metal2 4088 28280 4088 28280 0 net253
rlabel metal2 35784 29904 35784 29904 0 net254
rlabel metal2 8680 13496 8680 13496 0 net255
rlabel metal2 14056 29400 14056 29400 0 net256
rlabel metal2 29064 33656 29064 33656 0 net257
rlabel metal2 37688 16408 37688 16408 0 net258
rlabel metal2 18648 33656 18648 33656 0 net259
rlabel metal3 30296 4424 30296 4424 0 net26
rlabel metal2 18872 30912 18872 30912 0 net260
rlabel metal2 8008 31640 8008 31640 0 net261
rlabel metal2 43848 30128 43848 30128 0 net262
rlabel metal2 33768 21560 33768 21560 0 net263
rlabel metal2 9744 23912 9744 23912 0 net264
rlabel metal2 20216 19376 20216 19376 0 net265
rlabel metal2 30408 13832 30408 13832 0 net266
rlabel metal2 4088 24640 4088 24640 0 net267
rlabel metal2 9688 16240 9688 16240 0 net268
rlabel metal2 39984 13496 39984 13496 0 net269
rlabel metal3 21952 42728 21952 42728 0 net27
rlabel metal2 40544 31920 40544 31920 0 net270
rlabel metal2 37688 22344 37688 22344 0 net271
rlabel metal2 21784 31976 21784 31976 0 net272
rlabel metal2 18592 16744 18592 16744 0 net273
rlabel metal2 33432 29736 33432 29736 0 net274
rlabel metal2 6104 16464 6104 16464 0 net275
rlabel metal2 12488 20468 12488 20468 0 net276
rlabel metal2 15848 17976 15848 17976 0 net277
rlabel metal2 37352 27048 37352 27048 0 net278
rlabel metal2 7896 14056 7896 14056 0 net279
rlabel metal2 34104 3752 34104 3752 0 net28
rlabel metal2 39928 25200 39928 25200 0 net280
rlabel metal2 11928 33376 11928 33376 0 net281
rlabel metal2 20384 29960 20384 29960 0 net282
rlabel metal2 6552 30912 6552 30912 0 net283
rlabel metal3 21952 13608 21952 13608 0 net284
rlabel metal2 14616 15624 14616 15624 0 net285
rlabel metal2 44072 31444 44072 31444 0 net286
rlabel metal2 10024 32536 10024 32536 0 net287
rlabel metal2 8680 33376 8680 33376 0 net288
rlabel metal2 4872 34832 4872 34832 0 net289
rlabel metal2 10080 4536 10080 4536 0 net29
rlabel metal3 35000 19656 35000 19656 0 net290
rlabel metal2 38640 36568 38640 36568 0 net291
rlabel metal2 44968 38752 44968 38752 0 net292
rlabel metal2 6048 22344 6048 22344 0 net293
rlabel metal2 31192 16184 31192 16184 0 net294
rlabel metal2 14056 20468 14056 20468 0 net295
rlabel metal2 4480 16856 4480 16856 0 net296
rlabel metal3 33320 25480 33320 25480 0 net297
rlabel metal2 3864 13384 3864 13384 0 net298
rlabel metal2 10472 12936 10472 12936 0 net299
rlabel metal2 26264 5208 26264 5208 0 net3
rlabel metal2 26656 42728 26656 42728 0 net30
rlabel metal2 10640 9912 10640 9912 0 net300
rlabel metal2 4760 26544 4760 26544 0 net301
rlabel metal3 20272 4424 20272 4424 0 net31
rlabel metal3 36568 42728 36568 42728 0 net32
rlabel metal2 17304 5040 17304 5040 0 net33
rlabel metal2 21560 3416 21560 3416 0 net34
rlabel metal2 34552 4368 34552 4368 0 net35
rlabel metal2 35560 42784 35560 42784 0 net36
rlabel metal3 40544 4536 40544 4536 0 net37
rlabel metal2 44072 5824 44072 5824 0 net38
rlabel metal3 45024 4424 45024 4424 0 net39
rlabel metal2 7224 3584 7224 3584 0 net4
rlabel metal3 34496 4424 34496 4424 0 net40
rlabel metal2 34776 3864 34776 3864 0 net41
rlabel metal2 30520 4592 30520 4592 0 net42
rlabel metal2 44520 4256 44520 4256 0 net43
rlabel metal3 41272 42728 41272 42728 0 net44
rlabel metal2 27384 3864 27384 3864 0 net45
rlabel metal2 38808 3920 38808 3920 0 net46
rlabel metal2 7616 42728 7616 42728 0 net47
rlabel metal2 39088 42728 39088 42728 0 net48
rlabel metal2 27608 42000 27608 42000 0 net49
rlabel metal2 12544 3416 12544 3416 0 net5
rlabel metal2 31304 6048 31304 6048 0 net50
rlabel metal2 2072 5264 2072 5264 0 net51
rlabel metal3 35952 4536 35952 4536 0 net52
rlabel metal2 28280 5432 28280 5432 0 net53
rlabel metal2 18760 43176 18760 43176 0 net54
rlabel metal2 21728 42728 21728 42728 0 net55
rlabel metal2 32648 5600 32648 5600 0 net56
rlabel metal3 24864 6104 24864 6104 0 net57
rlabel metal2 38472 43064 38472 43064 0 net58
rlabel metal2 2072 3808 2072 3808 0 net59
rlabel metal3 20496 4536 20496 4536 0 net6
rlabel metal2 40264 43176 40264 43176 0 net60
rlabel metal2 2128 4536 2128 4536 0 net61
rlabel metal2 32200 25480 32200 25480 0 net62
rlabel metal2 44968 27720 44968 27720 0 net63
rlabel metal2 20776 4704 20776 4704 0 net64
rlabel metal2 18592 44072 18592 44072 0 net65
rlabel metal2 8904 5096 8904 5096 0 net66
rlabel metal2 44632 42504 44632 42504 0 net67
rlabel metal2 41384 4200 41384 4200 0 net68
rlabel metal2 39816 3752 39816 3752 0 net69
rlabel metal2 25592 43176 25592 43176 0 net7
rlabel metal2 32480 3528 32480 3528 0 net70
rlabel metal2 22456 3976 22456 3976 0 net71
rlabel metal2 44856 41608 44856 41608 0 net72
rlabel metal2 26376 4704 26376 4704 0 net73
rlabel metal2 30072 3808 30072 3808 0 net74
rlabel metal2 22120 42616 22120 42616 0 net75
rlabel metal2 36568 3640 36568 3640 0 net76
rlabel metal2 23464 5040 23464 5040 0 net77
rlabel metal2 26264 43064 26264 43064 0 net78
rlabel metal2 23800 44296 23800 44296 0 net79
rlabel metal2 14000 42728 14000 42728 0 net8
rlabel metal2 28616 4144 28616 4144 0 net80
rlabel metal2 13048 4592 13048 4592 0 net81
rlabel metal2 15064 4704 15064 4704 0 net82
rlabel metal2 18536 4368 18536 4368 0 net83
rlabel metal2 26096 44296 26096 44296 0 net84
rlabel metal2 14392 43876 14392 43876 0 net85
rlabel metal2 10584 4536 10584 4536 0 net86
rlabel metal3 24808 3528 24808 3528 0 net87
rlabel metal2 20216 4200 20216 4200 0 net88
rlabel metal2 16296 4200 16296 4200 0 net89
rlabel metal2 11928 3360 11928 3360 0 net9
rlabel metal3 28560 42168 28560 42168 0 net90
rlabel metal3 12040 3472 12040 3472 0 net91
rlabel metal2 28392 43876 28392 43876 0 net92
rlabel metal3 31360 42168 31360 42168 0 net93
rlabel metal2 13832 4200 13832 4200 0 net94
rlabel metal2 39536 44072 39536 44072 0 net95
rlabel metal2 27832 42840 27832 42840 0 net96
rlabel metal2 37240 4704 37240 4704 0 net97
rlabel metal2 2856 8120 2856 8120 0 net98
rlabel metal2 43848 11872 43848 11872 0 net99
rlabel metal2 46088 27384 46088 27384 0 pReset
rlabel metal2 22232 25144 22232 25144 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 48000 48000
<< end >>
