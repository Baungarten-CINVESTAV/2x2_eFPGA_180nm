magic
tech gf180mcuD
magscale 1 10
timestamp 1702149479
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 15598 42194 15650 42206
rect 15598 42130 15650 42142
rect 19406 42194 19458 42206
rect 19406 42130 19458 42142
rect 31166 42194 31218 42206
rect 31166 42130 31218 42142
rect 33182 42194 33234 42206
rect 33182 42130 33234 42142
rect 34750 42194 34802 42206
rect 34750 42130 34802 42142
rect 36654 42194 36706 42206
rect 36654 42130 36706 42142
rect 38446 42194 38498 42206
rect 38446 42130 38498 42142
rect 41358 42194 41410 42206
rect 41358 42130 41410 42142
rect 14142 42082 14194 42094
rect 14142 42018 14194 42030
rect 14814 42082 14866 42094
rect 14814 42018 14866 42030
rect 28366 42082 28418 42094
rect 28366 42018 28418 42030
rect 32846 42082 32898 42094
rect 32846 42018 32898 42030
rect 36318 42082 36370 42094
rect 36318 42018 36370 42030
rect 37550 42082 37602 42094
rect 37550 42018 37602 42030
rect 43822 42082 43874 42094
rect 43822 42018 43874 42030
rect 15262 41970 15314 41982
rect 16942 41970 16994 41982
rect 20862 41970 20914 41982
rect 13906 41918 13918 41970
rect 13970 41918 13982 41970
rect 14578 41918 14590 41970
rect 14642 41918 14654 41970
rect 16258 41918 16270 41970
rect 16322 41918 16334 41970
rect 20066 41918 20078 41970
rect 20130 41918 20142 41970
rect 15262 41906 15314 41918
rect 16942 41906 16994 41918
rect 20862 41906 20914 41918
rect 22430 41970 22482 41982
rect 22430 41906 22482 41918
rect 24558 41970 24610 41982
rect 24558 41906 24610 41918
rect 26462 41970 26514 41982
rect 26462 41906 26514 41918
rect 27918 41970 27970 41982
rect 32510 41970 32562 41982
rect 35534 41970 35586 41982
rect 28578 41918 28590 41970
rect 28642 41918 28654 41970
rect 33842 41918 33854 41970
rect 33906 41918 33918 41970
rect 27918 41906 27970 41918
rect 32510 41906 32562 41918
rect 35534 41906 35586 41918
rect 35982 41970 36034 41982
rect 35982 41906 36034 41918
rect 37214 41970 37266 41982
rect 37214 41906 37266 41918
rect 39230 41970 39282 41982
rect 39230 41906 39282 41918
rect 39790 41970 39842 41982
rect 39790 41906 39842 41918
rect 41806 41970 41858 41982
rect 41806 41906 41858 41918
rect 44158 41970 44210 41982
rect 44158 41906 44210 41918
rect 43150 41858 43202 41870
rect 17378 41806 17390 41858
rect 17442 41806 17454 41858
rect 21298 41806 21310 41858
rect 21362 41806 21374 41858
rect 22866 41806 22878 41858
rect 22930 41806 22942 41858
rect 24994 41806 25006 41858
rect 25058 41806 25070 41858
rect 26898 41806 26910 41858
rect 26962 41806 26974 41858
rect 40338 41806 40350 41858
rect 40402 41806 40414 41858
rect 42354 41806 42366 41858
rect 42418 41806 42430 41858
rect 43150 41794 43202 41806
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 14366 41298 14418 41310
rect 20190 41298 20242 41310
rect 19282 41246 19294 41298
rect 19346 41246 19358 41298
rect 14366 41234 14418 41246
rect 20190 41234 20242 41246
rect 21534 41298 21586 41310
rect 21534 41234 21586 41246
rect 23550 41298 23602 41310
rect 23550 41234 23602 41246
rect 24894 41298 24946 41310
rect 32510 41298 32562 41310
rect 27570 41246 27582 41298
rect 27634 41246 27646 41298
rect 24894 41234 24946 41246
rect 32510 41234 32562 41246
rect 37214 41298 37266 41310
rect 37214 41234 37266 41246
rect 37662 41298 37714 41310
rect 40338 41246 40350 41298
rect 40402 41246 40414 41298
rect 42018 41246 42030 41298
rect 42082 41246 42094 41298
rect 44034 41246 44046 41298
rect 44098 41246 44110 41298
rect 37662 41234 37714 41246
rect 17726 41186 17778 41198
rect 17726 41122 17778 41134
rect 20414 41186 20466 41198
rect 23774 41186 23826 41198
rect 37886 41186 37938 41198
rect 21970 41134 21982 41186
rect 22034 41134 22046 41186
rect 26002 41134 26014 41186
rect 26066 41134 26078 41186
rect 42466 41134 42478 41186
rect 42530 41134 42542 41186
rect 42914 41134 42926 41186
rect 42978 41134 42990 41186
rect 20414 41122 20466 41134
rect 23774 41122 23826 41134
rect 37886 41122 37938 41134
rect 17054 41074 17106 41086
rect 17054 41010 17106 41022
rect 25118 41074 25170 41086
rect 25118 41010 25170 41022
rect 31838 41074 31890 41086
rect 31838 41010 31890 41022
rect 16830 40962 16882 40974
rect 16830 40898 16882 40910
rect 18062 40962 18114 40974
rect 18062 40898 18114 40910
rect 18846 40962 18898 40974
rect 18846 40898 18898 40910
rect 20750 40962 20802 40974
rect 20750 40898 20802 40910
rect 21758 40962 21810 40974
rect 21758 40898 21810 40910
rect 24110 40962 24162 40974
rect 24110 40898 24162 40910
rect 25790 40962 25842 40974
rect 25790 40898 25842 40910
rect 27134 40962 27186 40974
rect 27134 40898 27186 40910
rect 38222 40962 38274 40974
rect 38222 40898 38274 40910
rect 39566 40962 39618 40974
rect 39566 40898 39618 40910
rect 39902 40962 39954 40974
rect 39902 40898 39954 40910
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 15150 40626 15202 40638
rect 15150 40562 15202 40574
rect 15822 40626 15874 40638
rect 15822 40562 15874 40574
rect 18846 40626 18898 40638
rect 18846 40562 18898 40574
rect 19742 40626 19794 40638
rect 19742 40562 19794 40574
rect 33406 40626 33458 40638
rect 33406 40562 33458 40574
rect 39454 40626 39506 40638
rect 39454 40562 39506 40574
rect 42590 40626 42642 40638
rect 42590 40562 42642 40574
rect 43710 40626 43762 40638
rect 43710 40562 43762 40574
rect 44158 40626 44210 40638
rect 44158 40562 44210 40574
rect 14814 40514 14866 40526
rect 14814 40450 14866 40462
rect 15486 40514 15538 40526
rect 15486 40450 15538 40462
rect 18510 40514 18562 40526
rect 18510 40450 18562 40462
rect 20078 40514 20130 40526
rect 20078 40450 20130 40462
rect 33070 40514 33122 40526
rect 33070 40450 33122 40462
rect 38782 40514 38834 40526
rect 38782 40450 38834 40462
rect 39118 40514 39170 40526
rect 39118 40450 39170 40462
rect 39790 40514 39842 40526
rect 39790 40450 39842 40462
rect 40350 40514 40402 40526
rect 40350 40450 40402 40462
rect 40910 40514 40962 40526
rect 40910 40450 40962 40462
rect 41918 40514 41970 40526
rect 41918 40450 41970 40462
rect 42926 40514 42978 40526
rect 42926 40450 42978 40462
rect 19506 40350 19518 40402
rect 19570 40350 19582 40402
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 41122 40350 41134 40402
rect 41186 40350 41198 40402
rect 41682 40350 41694 40402
rect 41746 40350 41758 40402
rect 42354 40350 42366 40402
rect 42418 40350 42430 40402
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 44158 39842 44210 39854
rect 44158 39778 44210 39790
rect 19854 39730 19906 39742
rect 19854 39666 19906 39678
rect 40686 39730 40738 39742
rect 40686 39666 40738 39678
rect 39118 39618 39170 39630
rect 41806 39618 41858 39630
rect 39890 39566 39902 39618
rect 39954 39566 39966 39618
rect 39118 39554 39170 39566
rect 41806 39554 41858 39566
rect 39454 39506 39506 39518
rect 39454 39442 39506 39454
rect 40126 39506 40178 39518
rect 40126 39442 40178 39454
rect 41470 39506 41522 39518
rect 41470 39442 41522 39454
rect 42142 39506 42194 39518
rect 42142 39442 42194 39454
rect 42478 39506 42530 39518
rect 42478 39442 42530 39454
rect 42814 39506 42866 39518
rect 42814 39442 42866 39454
rect 43374 39394 43426 39406
rect 43374 39330 43426 39342
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 42366 39058 42418 39070
rect 42366 38994 42418 39006
rect 43150 39058 43202 39070
rect 43150 38994 43202 39006
rect 43822 39058 43874 39070
rect 43822 38994 43874 39006
rect 42814 38946 42866 38958
rect 42814 38882 42866 38894
rect 43486 38946 43538 38958
rect 43486 38882 43538 38894
rect 44034 38782 44046 38834
rect 44098 38782 44110 38834
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 43150 38162 43202 38174
rect 43150 38098 43202 38110
rect 44034 37998 44046 38050
rect 44098 37998 44110 38050
rect 43822 37938 43874 37950
rect 43822 37874 43874 37886
rect 43486 37826 43538 37838
rect 43486 37762 43538 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 43822 37490 43874 37502
rect 43822 37426 43874 37438
rect 44158 37378 44210 37390
rect 44158 37314 44210 37326
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 43710 36370 43762 36382
rect 43710 36306 43762 36318
rect 44158 36258 44210 36270
rect 44158 36194 44210 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 20750 35922 20802 35934
rect 20750 35858 20802 35870
rect 21646 35922 21698 35934
rect 21646 35858 21698 35870
rect 24446 35922 24498 35934
rect 24446 35858 24498 35870
rect 25790 35922 25842 35934
rect 25790 35858 25842 35870
rect 26462 35922 26514 35934
rect 26462 35858 26514 35870
rect 24110 35810 24162 35822
rect 24110 35746 24162 35758
rect 44158 35810 44210 35822
rect 44158 35746 44210 35758
rect 20514 35646 20526 35698
rect 20578 35646 20590 35698
rect 21410 35646 21422 35698
rect 21474 35646 21486 35698
rect 25554 35646 25566 35698
rect 25618 35646 25630 35698
rect 26226 35646 26238 35698
rect 26290 35646 26302 35698
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 11442 31838 11454 31890
rect 11506 31838 11518 31890
rect 18498 31838 18510 31890
rect 18562 31838 18574 31890
rect 22306 31838 22318 31890
rect 22370 31838 22382 31890
rect 42914 31726 42926 31778
rect 42978 31726 42990 31778
rect 12450 31614 12462 31666
rect 12514 31614 12526 31666
rect 17378 31614 17390 31666
rect 17442 31614 17454 31666
rect 23538 31614 23550 31666
rect 23602 31614 23614 31666
rect 44034 31614 44046 31666
rect 44098 31614 44110 31666
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 42702 31218 42754 31230
rect 42702 31154 42754 31166
rect 22542 31106 22594 31118
rect 43822 31106 43874 31118
rect 14130 31054 14142 31106
rect 14194 31054 14206 31106
rect 28690 31054 28702 31106
rect 28754 31054 28766 31106
rect 31490 31054 31502 31106
rect 31554 31054 31566 31106
rect 34626 31054 34638 31106
rect 34690 31054 34702 31106
rect 22542 31042 22594 31054
rect 43822 31042 43874 31054
rect 19630 30994 19682 31006
rect 43598 30994 43650 31006
rect 20290 30942 20302 30994
rect 20354 30942 20366 30994
rect 42466 30942 42478 30994
rect 42530 30942 42542 30994
rect 19630 30930 19682 30942
rect 43598 30930 43650 30942
rect 44158 30994 44210 31006
rect 44158 30930 44210 30942
rect 12898 30830 12910 30882
rect 12962 30830 12974 30882
rect 27794 30830 27806 30882
rect 27858 30830 27870 30882
rect 30482 30830 30494 30882
rect 30546 30830 30558 30882
rect 35970 30830 35982 30882
rect 36034 30830 36046 30882
rect 23326 30770 23378 30782
rect 23326 30706 23378 30718
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 6626 30270 6638 30322
rect 6690 30270 6702 30322
rect 11218 30270 11230 30322
rect 11282 30270 11294 30322
rect 19170 30270 19182 30322
rect 19234 30270 19246 30322
rect 23090 30270 23102 30322
rect 23154 30270 23166 30322
rect 25890 30270 25902 30322
rect 25954 30270 25966 30322
rect 31042 30270 31054 30322
rect 31106 30270 31118 30322
rect 33842 30270 33854 30322
rect 33906 30270 33918 30322
rect 37986 30270 37998 30322
rect 38050 30270 38062 30322
rect 14478 30210 14530 30222
rect 14914 30158 14926 30210
rect 14978 30158 14990 30210
rect 14478 30146 14530 30158
rect 17950 30098 18002 30110
rect 21646 30098 21698 30110
rect 28030 30098 28082 30110
rect 7634 30046 7646 30098
rect 7698 30046 7710 30098
rect 9874 30046 9886 30098
rect 9938 30046 9950 30098
rect 20178 30046 20190 30098
rect 20242 30046 20254 30098
rect 21298 30046 21310 30098
rect 21362 30046 21374 30098
rect 24098 30046 24110 30098
rect 24162 30046 24174 30098
rect 26898 30046 26910 30098
rect 26962 30046 26974 30098
rect 27682 30046 27694 30098
rect 27746 30046 27758 30098
rect 17950 30034 18002 30046
rect 21646 30034 21698 30046
rect 28030 30034 28082 30046
rect 29486 30098 29538 30110
rect 35646 30098 35698 30110
rect 32050 30046 32062 30098
rect 32114 30046 32126 30098
rect 34850 30046 34862 30098
rect 34914 30046 34926 30098
rect 38994 30046 39006 30098
rect 39058 30046 39070 30098
rect 29486 30034 29538 30046
rect 35646 30034 35698 30046
rect 29374 29986 29426 29998
rect 17154 29934 17166 29986
rect 17218 29934 17230 29986
rect 29374 29922 29426 29934
rect 35758 29986 35810 29998
rect 35758 29922 35810 29934
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 5294 29650 5346 29662
rect 20974 29650 21026 29662
rect 24782 29650 24834 29662
rect 20402 29598 20414 29650
rect 20466 29598 20478 29650
rect 24210 29598 24222 29650
rect 24274 29598 24286 29650
rect 5294 29586 5346 29598
rect 20974 29586 21026 29598
rect 24782 29586 24834 29598
rect 25342 29650 25394 29662
rect 29362 29598 29374 29650
rect 29426 29598 29438 29650
rect 25342 29586 25394 29598
rect 4510 29538 4562 29550
rect 25230 29538 25282 29550
rect 8530 29486 8542 29538
rect 8594 29486 8606 29538
rect 13570 29486 13582 29538
rect 13634 29486 13646 29538
rect 16370 29486 16382 29538
rect 16434 29486 16446 29538
rect 35298 29486 35310 29538
rect 35362 29486 35374 29538
rect 37874 29486 37886 29538
rect 37938 29486 37950 29538
rect 4510 29474 4562 29486
rect 25230 29474 25282 29486
rect 1822 29426 1874 29438
rect 17502 29426 17554 29438
rect 21310 29426 21362 29438
rect 26238 29426 26290 29438
rect 2146 29374 2158 29426
rect 2210 29374 2222 29426
rect 17938 29374 17950 29426
rect 18002 29374 18014 29426
rect 21746 29374 21758 29426
rect 21810 29374 21822 29426
rect 26898 29374 26910 29426
rect 26962 29374 26974 29426
rect 1822 29362 1874 29374
rect 17502 29362 17554 29374
rect 21310 29362 21362 29374
rect 26238 29362 26290 29374
rect 31502 29314 31554 29326
rect 7522 29262 7534 29314
rect 7586 29262 7598 29314
rect 12562 29262 12574 29314
rect 12626 29262 12638 29314
rect 15362 29262 15374 29314
rect 15426 29262 15438 29314
rect 31826 29262 31838 29314
rect 31890 29262 31902 29314
rect 34066 29262 34078 29314
rect 34130 29262 34142 29314
rect 36866 29262 36878 29314
rect 36930 29262 36942 29314
rect 31502 29250 31554 29262
rect 29934 29202 29986 29214
rect 29934 29138 29986 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 11566 28866 11618 28878
rect 11566 28802 11618 28814
rect 16270 28866 16322 28878
rect 16270 28802 16322 28814
rect 27694 28866 27746 28878
rect 27694 28802 27746 28814
rect 32734 28866 32786 28878
rect 32734 28802 32786 28814
rect 36542 28866 36594 28878
rect 36542 28802 36594 28814
rect 4946 28702 4958 28754
rect 5010 28702 5022 28754
rect 15026 28702 15038 28754
rect 15090 28702 15102 28754
rect 20626 28702 20638 28754
rect 20690 28702 20702 28754
rect 22306 28702 22318 28754
rect 22370 28702 22382 28754
rect 41794 28702 41806 28754
rect 41858 28702 41870 28754
rect 5742 28642 5794 28654
rect 7422 28642 7474 28654
rect 4834 28590 4846 28642
rect 4898 28590 4910 28642
rect 6738 28590 6750 28642
rect 6802 28590 6814 28642
rect 5742 28578 5794 28590
rect 7422 28578 7474 28590
rect 7870 28642 7922 28654
rect 19742 28642 19794 28654
rect 23998 28642 24050 28654
rect 29038 28642 29090 28654
rect 33070 28642 33122 28654
rect 8418 28590 8430 28642
rect 8482 28590 8494 28642
rect 19394 28590 19406 28642
rect 19458 28590 19470 28642
rect 20514 28590 20526 28642
rect 20578 28590 20590 28642
rect 24658 28590 24670 28642
rect 24722 28590 24734 28642
rect 29698 28590 29710 28642
rect 29762 28590 29774 28642
rect 33506 28590 33518 28642
rect 33570 28590 33582 28642
rect 36978 28590 36990 28642
rect 37042 28590 37054 28642
rect 37538 28590 37550 28642
rect 37602 28590 37614 28642
rect 7870 28578 7922 28590
rect 19742 28578 19794 28590
rect 23998 28578 24050 28590
rect 29038 28578 29090 28590
rect 33070 28578 33122 28590
rect 27918 28530 27970 28542
rect 6962 28478 6974 28530
rect 7026 28478 7038 28530
rect 13682 28478 13694 28530
rect 13746 28478 13758 28530
rect 23538 28478 23550 28530
rect 23602 28478 23614 28530
rect 27918 28466 27970 28478
rect 31950 28530 32002 28542
rect 31950 28466 32002 28478
rect 35758 28530 35810 28542
rect 42802 28478 42814 28530
rect 42866 28478 42878 28530
rect 35758 28466 35810 28478
rect 28030 28418 28082 28430
rect 40574 28418 40626 28430
rect 10770 28366 10782 28418
rect 10834 28366 10846 28418
rect 17042 28366 17054 28418
rect 17106 28366 17118 28418
rect 27122 28366 27134 28418
rect 27186 28366 27198 28418
rect 40002 28366 40014 28418
rect 40066 28366 40078 28418
rect 28030 28354 28082 28366
rect 40574 28354 40626 28366
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 2046 28082 2098 28094
rect 10782 28082 10834 28094
rect 3042 28030 3054 28082
rect 3106 28030 3118 28082
rect 2046 28018 2098 28030
rect 10782 28018 10834 28030
rect 15262 28082 15314 28094
rect 15262 28018 15314 28030
rect 16718 28082 16770 28094
rect 32622 28082 32674 28094
rect 28018 28030 28030 28082
rect 28082 28030 28094 28082
rect 16718 28018 16770 28030
rect 32622 28018 32674 28030
rect 14478 27970 14530 27982
rect 23998 27970 24050 27982
rect 6626 27918 6638 27970
rect 6690 27918 6702 27970
rect 18834 27918 18846 27970
rect 18898 27918 18910 27970
rect 14478 27906 14530 27918
rect 23998 27906 24050 27918
rect 31838 27970 31890 27982
rect 31838 27906 31890 27918
rect 33742 27970 33794 27982
rect 33742 27906 33794 27918
rect 39678 27970 39730 27982
rect 39678 27906 39730 27918
rect 40462 27970 40514 27982
rect 42914 27918 42926 27970
rect 42978 27918 42990 27970
rect 40462 27906 40514 27918
rect 1710 27858 1762 27870
rect 5742 27858 5794 27870
rect 11566 27858 11618 27870
rect 21310 27858 21362 27870
rect 25118 27858 25170 27870
rect 36654 27858 36706 27870
rect 5282 27806 5294 27858
rect 5346 27806 5358 27858
rect 10770 27806 10782 27858
rect 10834 27806 10846 27858
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 21746 27806 21758 27858
rect 21810 27806 21822 27858
rect 25778 27806 25790 27858
rect 25842 27806 25854 27858
rect 29026 27806 29038 27858
rect 29090 27806 29102 27858
rect 29474 27806 29486 27858
rect 29538 27806 29550 27858
rect 35970 27806 35982 27858
rect 36034 27806 36046 27858
rect 1710 27794 1762 27806
rect 5742 27794 5794 27806
rect 11566 27794 11618 27806
rect 21310 27794 21362 27806
rect 25118 27794 25170 27806
rect 36654 27794 36706 27806
rect 36990 27858 37042 27870
rect 37426 27806 37438 27858
rect 37490 27806 37502 27858
rect 36990 27794 37042 27806
rect 9886 27746 9938 27758
rect 7970 27694 7982 27746
rect 8034 27694 8046 27746
rect 9538 27694 9550 27746
rect 9602 27694 9614 27746
rect 9886 27682 9938 27694
rect 15710 27746 15762 27758
rect 15710 27682 15762 27694
rect 16830 27746 16882 27758
rect 16830 27682 16882 27694
rect 17726 27746 17778 27758
rect 20974 27746 21026 27758
rect 18050 27694 18062 27746
rect 18114 27694 18126 27746
rect 19842 27694 19854 27746
rect 19906 27694 19918 27746
rect 41906 27694 41918 27746
rect 41970 27694 41982 27746
rect 17726 27682 17778 27694
rect 20974 27682 21026 27694
rect 2270 27634 2322 27646
rect 2270 27570 2322 27582
rect 24782 27634 24834 27646
rect 24782 27570 24834 27582
rect 28814 27634 28866 27646
rect 28814 27570 28866 27582
rect 32958 27634 33010 27646
rect 32958 27570 33010 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 9214 27298 9266 27310
rect 9214 27234 9266 27246
rect 13022 27298 13074 27310
rect 13022 27234 13074 27246
rect 22094 27298 22146 27310
rect 22094 27234 22146 27246
rect 27358 27298 27410 27310
rect 27358 27234 27410 27246
rect 34190 27298 34242 27310
rect 34190 27234 34242 27246
rect 40574 27298 40626 27310
rect 40574 27234 40626 27246
rect 1822 27186 1874 27198
rect 19406 27186 19458 27198
rect 4050 27134 4062 27186
rect 4114 27134 4126 27186
rect 14130 27134 14142 27186
rect 14194 27134 14206 27186
rect 23426 27134 23438 27186
rect 23490 27134 23502 27186
rect 35522 27134 35534 27186
rect 35586 27134 35598 27186
rect 41794 27134 41806 27186
rect 41858 27134 41870 27186
rect 1822 27122 1874 27134
rect 19406 27122 19458 27134
rect 5518 27074 5570 27086
rect 9326 27074 9378 27086
rect 15934 27074 15986 27086
rect 23886 27074 23938 27086
rect 30494 27074 30546 27086
rect 37102 27074 37154 27086
rect 6178 27022 6190 27074
rect 6242 27022 6254 27074
rect 9986 27022 9998 27074
rect 10050 27022 10062 27074
rect 13906 27022 13918 27074
rect 13970 27022 13982 27074
rect 16370 27022 16382 27074
rect 16434 27022 16446 27074
rect 19842 27022 19854 27074
rect 19906 27022 19918 27074
rect 20626 27022 20638 27074
rect 20690 27022 20702 27074
rect 24322 27022 24334 27074
rect 24386 27022 24398 27074
rect 31154 27022 31166 27074
rect 31218 27022 31230 27074
rect 34850 27022 34862 27074
rect 34914 27022 34926 27074
rect 37538 27022 37550 27074
rect 37602 27022 37614 27074
rect 5518 27010 5570 27022
rect 9326 27010 9378 27022
rect 15934 27010 15986 27022
rect 23886 27010 23938 27022
rect 30494 27010 30546 27022
rect 37102 27010 37154 27022
rect 12238 26962 12290 26974
rect 2706 26910 2718 26962
rect 2770 26910 2782 26962
rect 12238 26898 12290 26910
rect 14478 26962 14530 26974
rect 18622 26962 18674 26974
rect 23102 26962 23154 26974
rect 14802 26910 14814 26962
rect 14866 26910 14878 26962
rect 19618 26910 19630 26962
rect 19682 26910 19694 26962
rect 20402 26910 20414 26962
rect 20466 26910 20478 26962
rect 21522 26910 21534 26962
rect 21586 26910 21598 26962
rect 14478 26898 14530 26910
rect 18622 26898 18674 26910
rect 23102 26898 23154 26910
rect 26574 26962 26626 26974
rect 27918 26962 27970 26974
rect 27570 26910 27582 26962
rect 27634 26910 27646 26962
rect 26574 26898 26626 26910
rect 27918 26898 27970 26910
rect 29262 26962 29314 26974
rect 29262 26898 29314 26910
rect 36318 26962 36370 26974
rect 43598 26962 43650 26974
rect 42802 26910 42814 26962
rect 42866 26910 42878 26962
rect 43922 26910 43934 26962
rect 43986 26910 43998 26962
rect 36318 26898 36370 26910
rect 43598 26898 43650 26910
rect 15486 26850 15538 26862
rect 8642 26798 8654 26850
rect 8706 26798 8718 26850
rect 15486 26786 15538 26798
rect 29374 26850 29426 26862
rect 33394 26798 33406 26850
rect 33458 26798 33470 26850
rect 40002 26798 40014 26850
rect 40066 26798 40078 26850
rect 29374 26786 29426 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 7646 26514 7698 26526
rect 6962 26462 6974 26514
rect 7026 26462 7038 26514
rect 7646 26450 7698 26462
rect 33406 26514 33458 26526
rect 43822 26514 43874 26526
rect 36866 26462 36878 26514
rect 36930 26462 36942 26514
rect 33406 26450 33458 26462
rect 43822 26450 43874 26462
rect 37550 26402 37602 26414
rect 3042 26350 3054 26402
rect 3106 26350 3118 26402
rect 8642 26350 8654 26402
rect 8706 26350 8718 26402
rect 9762 26350 9774 26402
rect 9826 26350 9838 26402
rect 28578 26350 28590 26402
rect 28642 26350 28654 26402
rect 39778 26350 39790 26402
rect 39842 26350 39854 26402
rect 42914 26350 42926 26402
rect 42978 26350 42990 26402
rect 37550 26338 37602 26350
rect 2494 26290 2546 26302
rect 3950 26290 4002 26302
rect 34078 26290 34130 26302
rect 2818 26238 2830 26290
rect 2882 26238 2894 26290
rect 4498 26238 4510 26290
rect 4562 26238 4574 26290
rect 8866 26238 8878 26290
rect 8930 26238 8942 26290
rect 14802 26238 14814 26290
rect 14866 26238 14878 26290
rect 16706 26238 16718 26290
rect 16770 26238 16782 26290
rect 21858 26238 21870 26290
rect 21922 26238 21934 26290
rect 23202 26238 23214 26290
rect 23266 26238 23278 26290
rect 32162 26238 32174 26290
rect 32226 26238 32238 26290
rect 33394 26238 33406 26290
rect 33458 26238 33470 26290
rect 34514 26238 34526 26290
rect 34578 26238 34590 26290
rect 2494 26226 2546 26238
rect 3950 26226 4002 26238
rect 34078 26226 34130 26238
rect 3726 26178 3778 26190
rect 3378 26126 3390 26178
rect 3442 26126 3454 26178
rect 3726 26114 3778 26126
rect 8318 26178 8370 26190
rect 15486 26178 15538 26190
rect 15138 26126 15150 26178
rect 15202 26126 15214 26178
rect 8318 26114 8370 26126
rect 15486 26114 15538 26126
rect 15822 26178 15874 26190
rect 23774 26178 23826 26190
rect 16146 26126 16158 26178
rect 16210 26126 16222 26178
rect 16482 26126 16494 26178
rect 16546 26126 16558 26178
rect 19618 26126 19630 26178
rect 19682 26126 19694 26178
rect 22978 26126 22990 26178
rect 23042 26126 23054 26178
rect 15822 26114 15874 26126
rect 23774 26114 23826 26126
rect 26798 26178 26850 26190
rect 43710 26178 43762 26190
rect 38882 26126 38894 26178
rect 38946 26126 38958 26178
rect 41906 26126 41918 26178
rect 41970 26126 41982 26178
rect 26798 26114 26850 26126
rect 43710 26114 43762 26126
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 5518 25730 5570 25742
rect 5518 25666 5570 25678
rect 19854 25730 19906 25742
rect 19854 25666 19906 25678
rect 4510 25618 4562 25630
rect 20526 25618 20578 25630
rect 36430 25618 36482 25630
rect 3826 25566 3838 25618
rect 3890 25566 3902 25618
rect 14914 25566 14926 25618
rect 14978 25566 14990 25618
rect 20290 25566 20302 25618
rect 20354 25566 20366 25618
rect 22866 25566 22878 25618
rect 22930 25566 22942 25618
rect 25666 25566 25678 25618
rect 25730 25566 25742 25618
rect 30146 25566 30158 25618
rect 30210 25566 30222 25618
rect 32946 25566 32958 25618
rect 33010 25566 33022 25618
rect 35634 25566 35646 25618
rect 35698 25566 35710 25618
rect 4510 25554 4562 25566
rect 20526 25554 20578 25566
rect 36430 25554 36482 25566
rect 36990 25618 37042 25630
rect 42466 25566 42478 25618
rect 42530 25566 42542 25618
rect 36990 25554 37042 25566
rect 9214 25506 9266 25518
rect 12798 25506 12850 25518
rect 37550 25506 37602 25518
rect 8642 25454 8654 25506
rect 8706 25454 8718 25506
rect 12338 25454 12350 25506
rect 12402 25454 12414 25506
rect 16258 25454 16270 25506
rect 16322 25454 16334 25506
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 34850 25454 34862 25506
rect 34914 25454 34926 25506
rect 38210 25454 38222 25506
rect 38274 25454 38286 25506
rect 9214 25442 9266 25454
rect 12798 25442 12850 25454
rect 37550 25442 37602 25454
rect 6302 25394 6354 25406
rect 19070 25394 19122 25406
rect 41246 25394 41298 25406
rect 2706 25342 2718 25394
rect 2770 25342 2782 25394
rect 13570 25342 13582 25394
rect 13634 25342 13646 25394
rect 23874 25342 23886 25394
rect 23938 25342 23950 25394
rect 26898 25342 26910 25394
rect 26962 25342 26974 25394
rect 31490 25342 31502 25394
rect 31554 25342 31566 25394
rect 33954 25342 33966 25394
rect 34018 25342 34030 25394
rect 43698 25342 43710 25394
rect 43762 25342 43774 25394
rect 6302 25330 6354 25342
rect 19070 25330 19122 25342
rect 41246 25330 41298 25342
rect 9326 25282 9378 25294
rect 15486 25282 15538 25294
rect 10098 25230 10110 25282
rect 10162 25230 10174 25282
rect 9326 25218 9378 25230
rect 15486 25218 15538 25230
rect 15934 25282 15986 25294
rect 15934 25218 15986 25230
rect 32174 25282 32226 25294
rect 32174 25218 32226 25230
rect 32734 25282 32786 25294
rect 32734 25218 32786 25230
rect 37102 25282 37154 25294
rect 40674 25230 40686 25282
rect 40738 25230 40750 25282
rect 37102 25218 37154 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 2046 24946 2098 24958
rect 13134 24946 13186 24958
rect 2818 24894 2830 24946
rect 2882 24894 2894 24946
rect 12562 24894 12574 24946
rect 12626 24894 12638 24946
rect 2046 24882 2098 24894
rect 13134 24882 13186 24894
rect 13246 24946 13298 24958
rect 23326 24946 23378 24958
rect 14018 24894 14030 24946
rect 14082 24894 14094 24946
rect 22754 24894 22766 24946
rect 22818 24894 22830 24946
rect 29362 24894 29374 24946
rect 29426 24894 29438 24946
rect 13246 24882 13298 24894
rect 23326 24882 23378 24894
rect 31390 24834 31442 24846
rect 6962 24782 6974 24834
rect 7026 24782 7038 24834
rect 31714 24782 31726 24834
rect 31778 24782 31790 24834
rect 39330 24782 39342 24834
rect 39394 24782 39406 24834
rect 40002 24782 40014 24834
rect 40066 24782 40078 24834
rect 43138 24782 43150 24834
rect 43202 24782 43214 24834
rect 31390 24770 31442 24782
rect 9438 24722 9490 24734
rect 16942 24722 16994 24734
rect 19854 24722 19906 24734
rect 26462 24722 26514 24734
rect 31054 24722 31106 24734
rect 39678 24722 39730 24734
rect 5170 24670 5182 24722
rect 5234 24670 5246 24722
rect 5618 24670 5630 24722
rect 5682 24670 5694 24722
rect 10098 24670 10110 24722
rect 10162 24670 10174 24722
rect 16258 24670 16270 24722
rect 16322 24670 16334 24722
rect 18386 24670 18398 24722
rect 18450 24670 18462 24722
rect 20290 24670 20302 24722
rect 20354 24670 20366 24722
rect 27010 24670 27022 24722
rect 27074 24670 27086 24722
rect 32274 24670 32286 24722
rect 32338 24670 32350 24722
rect 33618 24670 33630 24722
rect 33682 24670 33694 24722
rect 9438 24658 9490 24670
rect 16942 24658 16994 24670
rect 19854 24658 19906 24670
rect 26462 24658 26514 24670
rect 31054 24658 31106 24670
rect 39678 24658 39730 24670
rect 19406 24610 19458 24622
rect 23886 24610 23938 24622
rect 7970 24558 7982 24610
rect 8034 24558 8046 24610
rect 19058 24558 19070 24610
rect 19122 24558 19134 24610
rect 23538 24558 23550 24610
rect 23602 24558 23614 24610
rect 19406 24546 19458 24558
rect 23886 24546 23938 24558
rect 30158 24610 30210 24622
rect 39006 24610 39058 24622
rect 32498 24558 32510 24610
rect 32562 24558 32574 24610
rect 35634 24558 35646 24610
rect 35698 24558 35710 24610
rect 41906 24558 41918 24610
rect 41970 24558 41982 24610
rect 30158 24546 30210 24558
rect 39006 24546 39058 24558
rect 17614 24498 17666 24510
rect 17614 24434 17666 24446
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 11902 24162 11954 24174
rect 11902 24098 11954 24110
rect 17166 24162 17218 24174
rect 17166 24098 17218 24110
rect 6750 24050 6802 24062
rect 4050 23998 4062 24050
rect 4114 23998 4126 24050
rect 6750 23986 6802 23998
rect 11006 24050 11058 24062
rect 16382 24050 16434 24062
rect 24334 24050 24386 24062
rect 13458 23998 13470 24050
rect 13522 23998 13534 24050
rect 15922 23998 15934 24050
rect 15986 23998 15998 24050
rect 23314 23998 23326 24050
rect 23378 23998 23390 24050
rect 36978 23998 36990 24050
rect 37042 23998 37054 24050
rect 43474 23998 43486 24050
rect 43538 23998 43550 24050
rect 11006 23986 11058 23998
rect 16382 23986 16434 23998
rect 24334 23986 24386 23998
rect 10446 23938 10498 23950
rect 20862 23938 20914 23950
rect 9986 23886 9998 23938
rect 10050 23886 10062 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 20178 23886 20190 23938
rect 20242 23886 20254 23938
rect 10446 23874 10498 23886
rect 20862 23874 20914 23886
rect 24558 23938 24610 23950
rect 29038 23938 29090 23950
rect 32846 23938 32898 23950
rect 38110 23938 38162 23950
rect 25218 23886 25230 23938
rect 25282 23886 25294 23938
rect 29698 23886 29710 23938
rect 29762 23886 29774 23938
rect 33506 23886 33518 23938
rect 33570 23886 33582 23938
rect 37202 23886 37214 23938
rect 37266 23886 37278 23938
rect 38770 23886 38782 23938
rect 38834 23886 38846 23938
rect 42242 23886 42254 23938
rect 42306 23886 42318 23938
rect 24558 23874 24610 23886
rect 29038 23874 29090 23886
rect 32846 23874 32898 23886
rect 38110 23874 38162 23886
rect 17950 23826 18002 23838
rect 3042 23774 3054 23826
rect 3106 23774 3118 23826
rect 6402 23774 6414 23826
rect 6466 23774 6478 23826
rect 11330 23774 11342 23826
rect 11394 23774 11406 23826
rect 12898 23774 12910 23826
rect 12962 23774 12974 23826
rect 14914 23774 14926 23826
rect 14978 23774 14990 23826
rect 22306 23774 22318 23826
rect 22370 23774 22382 23826
rect 42018 23774 42030 23826
rect 42082 23774 42094 23826
rect 17950 23762 18002 23774
rect 6974 23714 7026 23726
rect 16942 23714 16994 23726
rect 28254 23714 28306 23726
rect 32734 23714 32786 23726
rect 36542 23714 36594 23726
rect 41806 23714 41858 23726
rect 7634 23662 7646 23714
rect 7698 23662 7710 23714
rect 27682 23662 27694 23714
rect 27746 23662 27758 23714
rect 32162 23662 32174 23714
rect 32226 23662 32238 23714
rect 35970 23662 35982 23714
rect 36034 23662 36046 23714
rect 41234 23662 41246 23714
rect 41298 23662 41310 23714
rect 6974 23650 7026 23662
rect 16942 23650 16994 23662
rect 28254 23650 28306 23662
rect 32734 23650 32786 23662
rect 36542 23650 36594 23662
rect 41806 23650 41858 23662
rect 42926 23714 42978 23726
rect 42926 23650 42978 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 16942 23378 16994 23390
rect 32958 23378 33010 23390
rect 16146 23326 16158 23378
rect 16210 23326 16222 23378
rect 23426 23326 23438 23378
rect 23490 23326 23502 23378
rect 29922 23326 29934 23378
rect 29986 23326 29998 23378
rect 33506 23326 33518 23378
rect 33570 23326 33582 23378
rect 16942 23314 16994 23326
rect 32958 23314 33010 23326
rect 9438 23266 9490 23278
rect 4050 23214 4062 23266
rect 4114 23214 4126 23266
rect 6962 23214 6974 23266
rect 7026 23214 7038 23266
rect 9438 23202 9490 23214
rect 10222 23266 10274 23278
rect 39678 23266 39730 23278
rect 43710 23266 43762 23278
rect 18050 23214 18062 23266
rect 18114 23214 18126 23266
rect 31490 23214 31502 23266
rect 31554 23214 31566 23266
rect 32162 23214 32174 23266
rect 32226 23214 32238 23266
rect 42914 23214 42926 23266
rect 42978 23214 42990 23266
rect 10222 23202 10274 23214
rect 39678 23202 39730 23214
rect 43710 23202 43762 23214
rect 13134 23154 13186 23166
rect 20302 23154 20354 23166
rect 27134 23154 27186 23166
rect 36430 23154 36482 23166
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 13346 23102 13358 23154
rect 13410 23102 13422 23154
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 20850 23102 20862 23154
rect 20914 23102 20926 23154
rect 24546 23102 24558 23154
rect 24610 23102 24622 23154
rect 26226 23102 26238 23154
rect 26290 23102 26302 23154
rect 27570 23102 27582 23154
rect 27634 23102 27646 23154
rect 31714 23102 31726 23154
rect 31778 23102 31790 23154
rect 36082 23102 36094 23154
rect 36146 23102 36158 23154
rect 13134 23090 13186 23102
rect 20302 23090 20354 23102
rect 27134 23090 27186 23102
rect 36430 23090 36482 23102
rect 36766 23154 36818 23166
rect 37426 23102 37438 23154
rect 37490 23102 37502 23154
rect 36766 23090 36818 23102
rect 25454 23042 25506 23054
rect 31166 23042 31218 23054
rect 5170 22990 5182 23042
rect 5234 22990 5246 23042
rect 7970 22990 7982 23042
rect 8034 22990 8046 23042
rect 19058 22990 19070 23042
rect 19122 22990 19134 23042
rect 24322 22990 24334 23042
rect 24386 22990 24398 23042
rect 30818 22990 30830 23042
rect 30882 22990 30894 23042
rect 25454 22978 25506 22990
rect 31166 22978 31218 22990
rect 32510 23042 32562 23054
rect 41906 22990 41918 23042
rect 41970 22990 41982 23042
rect 43922 22990 43934 23042
rect 43986 22990 43998 23042
rect 32510 22978 32562 22990
rect 23998 22930 24050 22942
rect 23998 22866 24050 22878
rect 30606 22930 30658 22942
rect 30606 22866 30658 22878
rect 40462 22930 40514 22942
rect 40462 22866 40514 22878
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 9214 22594 9266 22606
rect 9214 22530 9266 22542
rect 33518 22594 33570 22606
rect 33518 22530 33570 22542
rect 13582 22482 13634 22494
rect 15822 22482 15874 22494
rect 4050 22430 4062 22482
rect 4114 22430 4126 22482
rect 15362 22430 15374 22482
rect 15426 22430 15438 22482
rect 13582 22418 13634 22430
rect 15822 22418 15874 22430
rect 27918 22482 27970 22494
rect 28478 22482 28530 22494
rect 28130 22430 28142 22482
rect 28194 22430 28206 22482
rect 34738 22430 34750 22482
rect 34802 22430 34814 22482
rect 41794 22430 41806 22482
rect 41858 22430 41870 22482
rect 27918 22418 27970 22430
rect 28478 22418 28530 22430
rect 5518 22370 5570 22382
rect 9326 22370 9378 22382
rect 20302 22370 20354 22382
rect 30046 22370 30098 22382
rect 36878 22370 36930 22382
rect 6066 22318 6078 22370
rect 6130 22318 6142 22370
rect 9874 22318 9886 22370
rect 9938 22318 9950 22370
rect 19730 22318 19742 22370
rect 19794 22318 19806 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 29362 22318 29374 22370
rect 29426 22318 29438 22370
rect 30482 22318 30494 22370
rect 30546 22318 30558 22370
rect 37538 22318 37550 22370
rect 37602 22318 37614 22370
rect 5518 22306 5570 22318
rect 9326 22306 9378 22318
rect 20302 22306 20354 22318
rect 30046 22306 30098 22318
rect 36878 22306 36930 22318
rect 16606 22258 16658 22270
rect 43598 22258 43650 22270
rect 3042 22206 3054 22258
rect 3106 22206 3118 22258
rect 14354 22206 14366 22258
rect 14418 22206 14430 22258
rect 23538 22206 23550 22258
rect 23602 22206 23614 22258
rect 29586 22206 29598 22258
rect 29650 22206 29662 22258
rect 35746 22206 35758 22258
rect 35810 22206 35822 22258
rect 42802 22206 42814 22258
rect 42866 22206 42878 22258
rect 16606 22194 16658 22206
rect 43598 22194 43650 22206
rect 13022 22146 13074 22158
rect 20862 22146 20914 22158
rect 33854 22146 33906 22158
rect 8642 22094 8654 22146
rect 8706 22094 8718 22146
rect 12338 22094 12350 22146
rect 12402 22094 12414 22146
rect 17378 22094 17390 22146
rect 17442 22094 17454 22146
rect 32946 22094 32958 22146
rect 33010 22094 33022 22146
rect 13022 22082 13074 22094
rect 20862 22082 20914 22094
rect 33854 22082 33906 22094
rect 34302 22146 34354 22158
rect 40574 22146 40626 22158
rect 40002 22094 40014 22146
rect 40066 22094 40078 22146
rect 34302 22082 34354 22094
rect 40574 22082 40626 22094
rect 41470 22146 41522 22158
rect 41470 22082 41522 22094
rect 43710 22146 43762 22158
rect 43710 22082 43762 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 12574 21810 12626 21822
rect 16942 21810 16994 21822
rect 21982 21810 22034 21822
rect 29822 21810 29874 21822
rect 2146 21758 2158 21810
rect 2210 21758 2222 21810
rect 6178 21758 6190 21810
rect 6242 21758 6254 21810
rect 16370 21758 16382 21810
rect 16434 21758 16446 21810
rect 21298 21758 21310 21810
rect 21362 21758 21374 21810
rect 28914 21758 28926 21810
rect 28978 21758 28990 21810
rect 37314 21758 37326 21810
rect 37378 21758 37390 21810
rect 12574 21746 12626 21758
rect 16942 21746 16994 21758
rect 21982 21746 22034 21758
rect 29822 21746 29874 21758
rect 38446 21698 38498 21710
rect 10994 21646 11006 21698
rect 11058 21646 11070 21698
rect 22642 21646 22654 21698
rect 22706 21646 22718 21698
rect 31938 21646 31950 21698
rect 32002 21646 32014 21698
rect 33058 21646 33070 21698
rect 33122 21646 33134 21698
rect 38446 21634 38498 21646
rect 39454 21698 39506 21710
rect 42914 21646 42926 21698
rect 42978 21646 42990 21698
rect 39454 21634 39506 21646
rect 5294 21586 5346 21598
rect 9102 21586 9154 21598
rect 25790 21586 25842 21598
rect 33406 21586 33458 21598
rect 4722 21534 4734 21586
rect 4786 21534 4798 21586
rect 8418 21534 8430 21586
rect 8482 21534 8494 21586
rect 9986 21534 9998 21586
rect 10050 21534 10062 21586
rect 13346 21534 13358 21586
rect 13410 21534 13422 21586
rect 13794 21534 13806 21586
rect 13858 21534 13870 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 18834 21534 18846 21586
rect 18898 21534 18910 21586
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 26450 21534 26462 21586
rect 26514 21534 26526 21586
rect 5294 21522 5346 21534
rect 9102 21522 9154 21534
rect 25790 21522 25842 21534
rect 33406 21522 33458 21534
rect 33854 21586 33906 21598
rect 33854 21522 33906 21534
rect 34190 21586 34242 21598
rect 43710 21586 43762 21598
rect 34850 21534 34862 21586
rect 34914 21534 34926 21586
rect 38098 21534 38110 21586
rect 38162 21534 38174 21586
rect 34190 21522 34242 21534
rect 43710 21522 43762 21534
rect 39118 21474 39170 21486
rect 10210 21422 10222 21474
rect 10274 21422 10286 21474
rect 12002 21422 12014 21474
rect 12066 21422 12078 21474
rect 23650 21422 23662 21474
rect 23714 21422 23726 21474
rect 25554 21422 25566 21474
rect 25618 21422 25630 21474
rect 30706 21422 30718 21474
rect 30770 21422 30782 21474
rect 38770 21422 38782 21474
rect 38834 21422 38846 21474
rect 39666 21422 39678 21474
rect 39730 21422 39742 21474
rect 41906 21422 41918 21474
rect 41970 21422 41982 21474
rect 43922 21422 43934 21474
rect 43986 21422 43998 21474
rect 39118 21410 39170 21422
rect 1598 21362 1650 21374
rect 1598 21298 1650 21310
rect 5406 21362 5458 21374
rect 5406 21298 5458 21310
rect 29486 21362 29538 21374
rect 29486 21298 29538 21310
rect 37886 21362 37938 21374
rect 37886 21298 37938 21310
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 13358 21026 13410 21038
rect 13358 20962 13410 20974
rect 22318 21026 22370 21038
rect 22318 20962 22370 20974
rect 35758 21026 35810 21038
rect 35758 20962 35810 20974
rect 22094 20914 22146 20926
rect 4050 20862 4062 20914
rect 4114 20862 4126 20914
rect 7634 20862 7646 20914
rect 7698 20862 7710 20914
rect 11890 20862 11902 20914
rect 11954 20862 11966 20914
rect 12562 20862 12574 20914
rect 12626 20862 12638 20914
rect 21858 20862 21870 20914
rect 21922 20862 21934 20914
rect 22094 20850 22146 20862
rect 29374 20914 29426 20926
rect 36430 20914 36482 20926
rect 37326 20914 37378 20926
rect 30146 20862 30158 20914
rect 30210 20862 30222 20914
rect 33170 20862 33182 20914
rect 33234 20862 33246 20914
rect 36978 20862 36990 20914
rect 37042 20862 37054 20914
rect 29374 20850 29426 20862
rect 36430 20850 36482 20862
rect 37326 20850 37378 20862
rect 42478 20914 42530 20926
rect 42690 20862 42702 20914
rect 42754 20862 42766 20914
rect 42478 20850 42530 20862
rect 7982 20802 8034 20814
rect 17054 20802 17106 20814
rect 8530 20750 8542 20802
rect 8594 20750 8606 20802
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 12786 20750 12798 20802
rect 12850 20750 12862 20802
rect 16370 20750 16382 20802
rect 16434 20750 16446 20802
rect 7982 20738 8034 20750
rect 17054 20738 17106 20750
rect 17390 20802 17442 20814
rect 25790 20802 25842 20814
rect 37774 20802 37826 20814
rect 17714 20750 17726 20802
rect 17778 20750 17790 20802
rect 25330 20750 25342 20802
rect 25394 20750 25406 20802
rect 28354 20750 28366 20802
rect 28418 20750 28430 20802
rect 34738 20750 34750 20802
rect 34802 20750 34814 20802
rect 38434 20750 38446 20802
rect 38498 20750 38510 20802
rect 17390 20738 17442 20750
rect 25790 20738 25842 20750
rect 37774 20738 37826 20750
rect 5966 20690 6018 20702
rect 3042 20638 3054 20690
rect 3106 20638 3118 20690
rect 5618 20638 5630 20690
rect 5682 20638 5694 20690
rect 5966 20626 6018 20638
rect 7422 20690 7474 20702
rect 7422 20626 7474 20638
rect 10894 20690 10946 20702
rect 10894 20626 10946 20638
rect 23102 20690 23154 20702
rect 31154 20638 31166 20690
rect 31218 20638 31230 20690
rect 33954 20638 33966 20690
rect 34018 20638 34030 20690
rect 43698 20638 43710 20690
rect 43762 20638 43774 20690
rect 23102 20626 23154 20638
rect 11678 20578 11730 20590
rect 20862 20578 20914 20590
rect 13906 20526 13918 20578
rect 13970 20526 13982 20578
rect 20290 20526 20302 20578
rect 20354 20526 20366 20578
rect 11678 20514 11730 20526
rect 20862 20514 20914 20526
rect 28366 20578 28418 20590
rect 41470 20578 41522 20590
rect 40898 20526 40910 20578
rect 40962 20526 40974 20578
rect 28366 20514 28418 20526
rect 41470 20514 41522 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 21858 20190 21870 20242
rect 21922 20190 21934 20242
rect 3278 20130 3330 20142
rect 3278 20066 3330 20078
rect 6750 20130 6802 20142
rect 8990 20130 9042 20142
rect 20190 20130 20242 20142
rect 8642 20078 8654 20130
rect 8706 20078 8718 20130
rect 9762 20078 9774 20130
rect 9826 20078 9838 20130
rect 6750 20066 6802 20078
rect 8990 20066 9042 20078
rect 20190 20066 20242 20078
rect 28814 20130 28866 20142
rect 36206 20130 36258 20142
rect 31938 20078 31950 20130
rect 32002 20078 32014 20130
rect 39218 20078 39230 20130
rect 39282 20078 39294 20130
rect 42914 20078 42926 20130
rect 42978 20078 42990 20130
rect 28814 20066 28866 20078
rect 36206 20066 36258 20078
rect 4062 20018 4114 20030
rect 17502 20018 17554 20030
rect 24558 20018 24610 20030
rect 33518 20018 33570 20030
rect 4386 19966 4398 20018
rect 4450 19966 4462 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 16146 19966 16158 20018
rect 16210 19966 16222 20018
rect 17938 19966 17950 20018
rect 18002 19966 18014 20018
rect 24098 19966 24110 20018
rect 24162 19966 24174 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 26002 19966 26014 20018
rect 26066 19966 26078 20018
rect 26450 19966 26462 20018
rect 26514 19966 26526 20018
rect 33954 19966 33966 20018
rect 34018 19966 34030 20018
rect 4062 19954 4114 19966
rect 17502 19954 17554 19966
rect 24558 19954 24610 19966
rect 33518 19954 33570 19966
rect 7982 19906 8034 19918
rect 16830 19906 16882 19918
rect 30046 19906 30098 19918
rect 3602 19854 3614 19906
rect 3666 19854 3678 19906
rect 8306 19854 8318 19906
rect 8370 19854 8382 19906
rect 25218 19854 25230 19906
rect 25282 19854 25294 19906
rect 7982 19842 8034 19854
rect 16830 19842 16882 19854
rect 30046 19842 30098 19854
rect 30494 19906 30546 19918
rect 37326 19906 37378 19918
rect 30818 19854 30830 19906
rect 30882 19854 30894 19906
rect 38210 19854 38222 19906
rect 38274 19854 38286 19906
rect 41906 19854 41918 19906
rect 41970 19854 41982 19906
rect 30494 19842 30546 19854
rect 37326 19842 37378 19854
rect 7534 19794 7586 19806
rect 7534 19730 7586 19742
rect 15822 19794 15874 19806
rect 15822 19730 15874 19742
rect 20974 19794 21026 19806
rect 20974 19730 21026 19742
rect 21086 19794 21138 19806
rect 21086 19730 21138 19742
rect 29598 19794 29650 19806
rect 29598 19730 29650 19742
rect 36990 19794 37042 19806
rect 36990 19730 37042 19742
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 12462 19458 12514 19470
rect 12462 19394 12514 19406
rect 42814 19458 42866 19470
rect 42814 19394 42866 19406
rect 6974 19346 7026 19358
rect 21646 19346 21698 19358
rect 3938 19294 3950 19346
rect 4002 19294 4014 19346
rect 6290 19294 6302 19346
rect 6354 19294 6366 19346
rect 19954 19294 19966 19346
rect 20018 19294 20030 19346
rect 21298 19294 21310 19346
rect 21362 19294 21374 19346
rect 22082 19294 22094 19346
rect 22146 19294 22158 19346
rect 37874 19294 37886 19346
rect 37938 19294 37950 19346
rect 6974 19282 7026 19294
rect 21646 19282 21698 19294
rect 7198 19234 7250 19246
rect 20302 19234 20354 19246
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 7746 19182 7758 19234
rect 7810 19182 7822 19234
rect 15026 19182 15038 19234
rect 15090 19182 15102 19234
rect 7198 19170 7250 19182
rect 20302 19170 20354 19182
rect 22430 19234 22482 19246
rect 22430 19170 22482 19182
rect 23886 19234 23938 19246
rect 32734 19234 32786 19246
rect 36542 19234 36594 19246
rect 39118 19234 39170 19246
rect 24322 19182 24334 19234
rect 24386 19182 24398 19234
rect 32162 19182 32174 19234
rect 32226 19182 32238 19234
rect 35970 19182 35982 19234
rect 36034 19182 36046 19234
rect 37202 19182 37214 19234
rect 37266 19182 37278 19234
rect 39778 19182 39790 19234
rect 39842 19182 39854 19234
rect 23886 19170 23938 19182
rect 32734 19170 32786 19182
rect 36542 19170 36594 19182
rect 39118 19170 39170 19182
rect 10110 19122 10162 19134
rect 13806 19122 13858 19134
rect 26574 19122 26626 19134
rect 2034 19070 2046 19122
rect 2098 19070 2110 19122
rect 3042 19070 3054 19122
rect 3106 19070 3118 19122
rect 6626 19070 6638 19122
rect 6690 19070 6702 19122
rect 11442 19070 11454 19122
rect 11506 19070 11518 19122
rect 13458 19070 13470 19122
rect 13522 19070 13534 19122
rect 18386 19070 18398 19122
rect 18450 19070 18462 19122
rect 10110 19058 10162 19070
rect 13806 19058 13858 19070
rect 26574 19058 26626 19070
rect 28254 19122 28306 19134
rect 28254 19058 28306 19070
rect 33630 19122 33682 19134
rect 33630 19058 33682 19070
rect 38894 19122 38946 19134
rect 38894 19058 38946 19070
rect 1710 19010 1762 19022
rect 1710 18946 1762 18958
rect 10894 19010 10946 19022
rect 10894 18946 10946 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 27358 19010 27410 19022
rect 27358 18946 27410 18958
rect 27694 19010 27746 19022
rect 27694 18946 27746 18958
rect 28366 19010 28418 19022
rect 28366 18946 28418 18958
rect 29038 19010 29090 19022
rect 32846 19010 32898 19022
rect 29698 18958 29710 19010
rect 29762 18958 29774 19010
rect 29038 18946 29090 18958
rect 32846 18946 32898 18958
rect 38782 19010 38834 19022
rect 42242 18958 42254 19010
rect 42306 18958 42318 19010
rect 38782 18946 38834 18958
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 1822 18674 1874 18686
rect 4946 18622 4958 18674
rect 5010 18622 5022 18674
rect 15586 18622 15598 18674
rect 15650 18622 15662 18674
rect 20514 18622 20526 18674
rect 20578 18622 20590 18674
rect 1822 18610 1874 18622
rect 21646 18562 21698 18574
rect 6962 18510 6974 18562
rect 7026 18510 7038 18562
rect 9986 18510 9998 18562
rect 10050 18510 10062 18562
rect 24546 18510 24558 18562
rect 24610 18510 24622 18562
rect 30034 18510 30046 18562
rect 30098 18510 30110 18562
rect 42914 18510 42926 18562
rect 42978 18510 42990 18562
rect 21646 18498 21698 18510
rect 2270 18450 2322 18462
rect 12686 18450 12738 18462
rect 17614 18450 17666 18462
rect 26462 18450 26514 18462
rect 32510 18450 32562 18462
rect 2706 18398 2718 18450
rect 2770 18398 2782 18450
rect 13010 18398 13022 18450
rect 13074 18398 13086 18450
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 32050 18398 32062 18450
rect 32114 18398 32126 18450
rect 33058 18398 33070 18450
rect 33122 18398 33134 18450
rect 38770 18398 38782 18450
rect 38834 18398 38846 18450
rect 39330 18398 39342 18450
rect 39394 18398 39406 18450
rect 39554 18398 39566 18450
rect 39618 18398 39630 18450
rect 40226 18398 40238 18450
rect 40290 18398 40302 18450
rect 2270 18386 2322 18398
rect 12686 18386 12738 18398
rect 17614 18386 17666 18398
rect 26462 18386 26514 18398
rect 32510 18386 32562 18398
rect 16830 18338 16882 18350
rect 22094 18338 22146 18350
rect 25342 18338 25394 18350
rect 7970 18286 7982 18338
rect 8034 18286 8046 18338
rect 11218 18286 11230 18338
rect 11282 18286 11294 18338
rect 16482 18286 16494 18338
rect 16546 18286 16558 18338
rect 21410 18286 21422 18338
rect 21474 18286 21486 18338
rect 23202 18286 23214 18338
rect 23266 18286 23278 18338
rect 16830 18274 16882 18286
rect 22094 18274 22146 18286
rect 25342 18274 25394 18286
rect 26014 18338 26066 18350
rect 36530 18286 36542 18338
rect 36594 18286 36606 18338
rect 38994 18286 39006 18338
rect 39058 18286 39070 18338
rect 40002 18286 40014 18338
rect 40066 18286 40078 18338
rect 41906 18286 41918 18338
rect 41970 18286 41982 18338
rect 26014 18274 26066 18286
rect 5742 18226 5794 18238
rect 5742 18162 5794 18174
rect 16158 18226 16210 18238
rect 16158 18162 16210 18174
rect 21086 18226 21138 18238
rect 21086 18162 21138 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 5518 17890 5570 17902
rect 5518 17826 5570 17838
rect 26014 17890 26066 17902
rect 26014 17826 26066 17838
rect 43598 17778 43650 17790
rect 2146 17726 2158 17778
rect 2210 17726 2222 17778
rect 3938 17726 3950 17778
rect 4002 17726 4014 17778
rect 21410 17726 21422 17778
rect 21474 17726 21486 17778
rect 41794 17726 41806 17778
rect 41858 17726 41870 17778
rect 43598 17714 43650 17726
rect 9214 17666 9266 17678
rect 17054 17666 17106 17678
rect 20862 17666 20914 17678
rect 8530 17614 8542 17666
rect 8594 17614 8606 17666
rect 9426 17614 9438 17666
rect 9490 17614 9502 17666
rect 9874 17614 9886 17666
rect 9938 17614 9950 17666
rect 16482 17614 16494 17666
rect 16546 17614 16558 17666
rect 20178 17614 20190 17666
rect 20242 17614 20254 17666
rect 9214 17602 9266 17614
rect 17054 17602 17106 17614
rect 20862 17602 20914 17614
rect 22318 17666 22370 17678
rect 32510 17666 32562 17678
rect 36542 17666 36594 17678
rect 22978 17614 22990 17666
rect 23042 17614 23054 17666
rect 27346 17614 27358 17666
rect 27410 17614 27422 17666
rect 32162 17614 32174 17666
rect 32226 17614 32238 17666
rect 35970 17614 35982 17666
rect 36034 17614 36046 17666
rect 36978 17614 36990 17666
rect 37042 17614 37054 17666
rect 37538 17614 37550 17666
rect 37602 17614 37614 17666
rect 22318 17602 22370 17614
rect 32510 17602 32562 17614
rect 36542 17602 36594 17614
rect 1934 17554 1986 17566
rect 14142 17554 14194 17566
rect 3042 17502 3054 17554
rect 3106 17502 3118 17554
rect 1934 17490 1986 17502
rect 14142 17490 14194 17502
rect 21646 17554 21698 17566
rect 21646 17490 21698 17502
rect 25230 17554 25282 17566
rect 26910 17554 26962 17566
rect 39790 17554 39842 17566
rect 26562 17502 26574 17554
rect 26626 17502 26638 17554
rect 28130 17502 28142 17554
rect 28194 17502 28206 17554
rect 42802 17502 42814 17554
rect 42866 17502 42878 17554
rect 43922 17502 43934 17554
rect 43986 17502 43998 17554
rect 25230 17490 25282 17502
rect 26910 17490 26962 17502
rect 39790 17490 39842 17502
rect 13022 17442 13074 17454
rect 6290 17390 6302 17442
rect 6354 17390 6366 17442
rect 12450 17390 12462 17442
rect 12514 17390 12526 17442
rect 13022 17378 13074 17390
rect 13358 17442 13410 17454
rect 13358 17378 13410 17390
rect 17166 17442 17218 17454
rect 22094 17442 22146 17454
rect 17714 17390 17726 17442
rect 17778 17390 17790 17442
rect 17166 17378 17218 17390
rect 22094 17378 22146 17390
rect 29038 17442 29090 17454
rect 32846 17442 32898 17454
rect 40574 17442 40626 17454
rect 29586 17390 29598 17442
rect 29650 17390 29662 17442
rect 33618 17390 33630 17442
rect 33682 17390 33694 17442
rect 29038 17378 29090 17390
rect 32846 17378 32898 17390
rect 40574 17378 40626 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 32622 17106 32674 17118
rect 36654 17106 36706 17118
rect 2146 17054 2158 17106
rect 2210 17054 2222 17106
rect 6178 17054 6190 17106
rect 6242 17054 6254 17106
rect 12562 17054 12574 17106
rect 12626 17054 12638 17106
rect 16370 17054 16382 17106
rect 16434 17054 16446 17106
rect 36082 17054 36094 17106
rect 36146 17054 36158 17106
rect 39890 17054 39902 17106
rect 39954 17054 39966 17106
rect 32622 17042 32674 17054
rect 36654 17042 36706 17054
rect 18846 16994 18898 17006
rect 25902 16994 25954 17006
rect 22530 16942 22542 16994
rect 22594 16942 22606 16994
rect 18846 16930 18898 16942
rect 25902 16930 25954 16942
rect 31838 16994 31890 17006
rect 43710 16994 43762 17006
rect 42914 16942 42926 16994
rect 42978 16942 42990 16994
rect 31838 16930 31890 16942
rect 43710 16930 43762 16942
rect 5070 16882 5122 16894
rect 8878 16882 8930 16894
rect 4722 16830 4734 16882
rect 4786 16830 4798 16882
rect 8418 16830 8430 16882
rect 8482 16830 8494 16882
rect 5070 16818 5122 16830
rect 8878 16818 8930 16830
rect 9438 16882 9490 16894
rect 13246 16882 13298 16894
rect 21758 16882 21810 16894
rect 28590 16882 28642 16894
rect 10098 16830 10110 16882
rect 10162 16830 10174 16882
rect 13906 16830 13918 16882
rect 13970 16830 13982 16882
rect 21186 16830 21198 16882
rect 21250 16830 21262 16882
rect 28242 16830 28254 16882
rect 28306 16830 28318 16882
rect 9438 16818 9490 16830
rect 13246 16818 13298 16830
rect 21758 16818 21810 16830
rect 28590 16818 28642 16830
rect 28926 16882 28978 16894
rect 33182 16882 33234 16894
rect 36990 16882 37042 16894
rect 29586 16830 29598 16882
rect 29650 16830 29662 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 37426 16830 37438 16882
rect 37490 16830 37502 16882
rect 28926 16818 28978 16830
rect 33182 16818 33234 16830
rect 36990 16818 37042 16830
rect 17838 16770 17890 16782
rect 17490 16718 17502 16770
rect 17554 16718 17566 16770
rect 23426 16718 23438 16770
rect 23490 16718 23502 16770
rect 41906 16718 41918 16770
rect 41970 16718 41982 16770
rect 44034 16718 44046 16770
rect 44098 16718 44110 16770
rect 17838 16706 17890 16718
rect 1598 16658 1650 16670
rect 1598 16594 1650 16606
rect 5406 16658 5458 16670
rect 5406 16594 5458 16606
rect 13134 16658 13186 16670
rect 13134 16594 13186 16606
rect 16942 16658 16994 16670
rect 16942 16594 16994 16606
rect 18062 16658 18114 16670
rect 18062 16594 18114 16606
rect 25118 16658 25170 16670
rect 25118 16594 25170 16606
rect 40462 16658 40514 16670
rect 40462 16594 40514 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 26910 16210 26962 16222
rect 28590 16210 28642 16222
rect 3826 16158 3838 16210
rect 3890 16158 3902 16210
rect 15474 16158 15486 16210
rect 15538 16158 15550 16210
rect 27794 16158 27806 16210
rect 27858 16158 27870 16210
rect 41794 16158 41806 16210
rect 41858 16158 41870 16210
rect 26910 16146 26962 16158
rect 28590 16146 28642 16158
rect 1934 16098 1986 16110
rect 11342 16098 11394 16110
rect 20190 16098 20242 16110
rect 29038 16098 29090 16110
rect 33070 16098 33122 16110
rect 40350 16098 40402 16110
rect 10770 16046 10782 16098
rect 10834 16046 10846 16098
rect 11554 16046 11566 16098
rect 11618 16046 11630 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 22754 16046 22766 16098
rect 22818 16046 22830 16098
rect 23314 16046 23326 16098
rect 23378 16046 23390 16098
rect 29698 16046 29710 16098
rect 29762 16046 29774 16098
rect 33506 16046 33518 16098
rect 33570 16046 33582 16098
rect 40002 16046 40014 16098
rect 40066 16046 40078 16098
rect 1934 16034 1986 16046
rect 11342 16034 11394 16046
rect 20190 16034 20242 16046
rect 29038 16034 29090 16046
rect 33070 16034 33122 16046
rect 40350 16034 40402 16046
rect 6302 15986 6354 15998
rect 17502 15986 17554 15998
rect 2706 15934 2718 15986
rect 2770 15934 2782 15986
rect 5954 15934 5966 15986
rect 6018 15934 6030 15986
rect 14354 15934 14366 15986
rect 14418 15934 14430 15986
rect 6302 15922 6354 15934
rect 17502 15922 17554 15934
rect 21982 15986 22034 15998
rect 21982 15922 22034 15934
rect 27470 15986 27522 15998
rect 27470 15922 27522 15934
rect 28142 15986 28194 15998
rect 28142 15922 28194 15934
rect 37662 15986 37714 15998
rect 42802 15934 42814 15986
rect 42866 15934 42878 15986
rect 37662 15922 37714 15934
rect 2046 15874 2098 15886
rect 2046 15810 2098 15822
rect 7646 15874 7698 15886
rect 12126 15874 12178 15886
rect 8418 15822 8430 15874
rect 8482 15822 8494 15874
rect 7646 15810 7698 15822
rect 12126 15810 12178 15822
rect 16718 15874 16770 15886
rect 16718 15810 16770 15822
rect 22094 15874 22146 15886
rect 26350 15874 26402 15886
rect 25778 15822 25790 15874
rect 25842 15822 25854 15874
rect 22094 15810 22146 15822
rect 26350 15810 26402 15822
rect 27358 15874 27410 15886
rect 32734 15874 32786 15886
rect 36542 15874 36594 15886
rect 32050 15822 32062 15874
rect 32114 15822 32126 15874
rect 35970 15822 35982 15874
rect 36034 15822 36046 15874
rect 27358 15810 27410 15822
rect 32734 15810 32786 15822
rect 36542 15810 36594 15822
rect 36878 15874 36930 15886
rect 36878 15810 36930 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 25342 15538 25394 15550
rect 32510 15538 32562 15550
rect 4946 15486 4958 15538
rect 5010 15486 5022 15538
rect 24210 15486 24222 15538
rect 24274 15486 24286 15538
rect 30258 15486 30270 15538
rect 30322 15486 30334 15538
rect 38098 15486 38110 15538
rect 38162 15486 38174 15538
rect 25342 15474 25394 15486
rect 32510 15474 32562 15486
rect 10222 15426 10274 15438
rect 11454 15426 11506 15438
rect 7970 15374 7982 15426
rect 8034 15374 8046 15426
rect 9874 15374 9886 15426
rect 9938 15374 9950 15426
rect 11106 15374 11118 15426
rect 11170 15374 11182 15426
rect 10222 15362 10274 15374
rect 11454 15362 11506 15374
rect 12462 15426 12514 15438
rect 26126 15426 26178 15438
rect 31390 15426 31442 15438
rect 15586 15374 15598 15426
rect 15650 15374 15662 15426
rect 17714 15374 17726 15426
rect 17778 15374 17790 15426
rect 20738 15374 20750 15426
rect 20802 15374 20814 15426
rect 25778 15374 25790 15426
rect 25842 15374 25854 15426
rect 26450 15374 26462 15426
rect 26514 15374 26526 15426
rect 31042 15374 31054 15426
rect 31106 15374 31118 15426
rect 12462 15362 12514 15374
rect 26126 15362 26178 15374
rect 31390 15362 31442 15374
rect 31726 15426 31778 15438
rect 32050 15374 32062 15426
rect 32114 15374 32126 15426
rect 33058 15374 33070 15426
rect 33122 15374 33134 15426
rect 34402 15374 34414 15426
rect 34466 15374 34478 15426
rect 38882 15374 38894 15426
rect 38946 15374 38958 15426
rect 42914 15374 42926 15426
rect 42978 15374 42990 15426
rect 31726 15362 31778 15374
rect 2270 15314 2322 15326
rect 15374 15314 15426 15326
rect 2706 15262 2718 15314
rect 2770 15262 2782 15314
rect 14802 15262 14814 15314
rect 14866 15262 14878 15314
rect 2270 15250 2322 15262
rect 15374 15250 15426 15262
rect 21310 15314 21362 15326
rect 27134 15314 27186 15326
rect 33742 15314 33794 15326
rect 21746 15262 21758 15314
rect 21810 15262 21822 15314
rect 26674 15262 26686 15314
rect 26738 15262 26750 15314
rect 27794 15262 27806 15314
rect 27858 15262 27870 15314
rect 33282 15262 33294 15314
rect 33346 15262 33358 15314
rect 21310 15250 21362 15262
rect 27134 15250 27186 15262
rect 33742 15250 33794 15262
rect 34974 15314 35026 15326
rect 35634 15262 35646 15314
rect 35698 15262 35710 15314
rect 39106 15262 39118 15314
rect 39170 15262 39182 15314
rect 34974 15250 35026 15262
rect 15934 15202 15986 15214
rect 6962 15150 6974 15202
rect 7026 15150 7038 15202
rect 15934 15138 15986 15150
rect 18062 15202 18114 15214
rect 34750 15202 34802 15214
rect 19618 15150 19630 15202
rect 19682 15150 19694 15202
rect 33954 15150 33966 15202
rect 34018 15150 34030 15202
rect 41906 15150 41918 15202
rect 41970 15150 41982 15202
rect 18062 15138 18114 15150
rect 34750 15138 34802 15150
rect 5742 15090 5794 15102
rect 5742 15026 5794 15038
rect 11678 15090 11730 15102
rect 11678 15026 11730 15038
rect 24782 15090 24834 15102
rect 24782 15026 24834 15038
rect 30830 15090 30882 15102
rect 30830 15026 30882 15038
rect 38670 15090 38722 15102
rect 38670 15026 38722 15038
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 28130 14751 28142 14754
rect 27585 14705 28142 14751
rect 14366 14642 14418 14654
rect 15038 14642 15090 14654
rect 27246 14642 27298 14654
rect 27585 14642 27631 14705
rect 28130 14702 28142 14705
rect 28194 14751 28206 14754
rect 28578 14751 28590 14754
rect 28194 14705 28590 14751
rect 28194 14702 28206 14705
rect 28578 14702 28590 14705
rect 28642 14702 28654 14754
rect 27694 14642 27746 14654
rect 3490 14590 3502 14642
rect 3554 14590 3566 14642
rect 7410 14590 7422 14642
rect 7474 14590 7486 14642
rect 11442 14590 11454 14642
rect 11506 14590 11518 14642
rect 14018 14590 14030 14642
rect 14082 14590 14094 14642
rect 14690 14590 14702 14642
rect 14754 14590 14766 14642
rect 16818 14590 16830 14642
rect 16882 14590 16894 14642
rect 19730 14590 19742 14642
rect 19794 14590 19806 14642
rect 21410 14590 21422 14642
rect 21474 14590 21486 14642
rect 27570 14590 27582 14642
rect 27634 14590 27646 14642
rect 14366 14578 14418 14590
rect 15038 14578 15090 14590
rect 27246 14578 27298 14590
rect 27694 14578 27746 14590
rect 28142 14642 28194 14654
rect 28142 14578 28194 14590
rect 28590 14642 28642 14654
rect 34290 14590 34302 14642
rect 34354 14590 34366 14642
rect 36082 14590 36094 14642
rect 36146 14590 36158 14642
rect 41794 14590 41806 14642
rect 41858 14590 41870 14642
rect 28590 14578 28642 14590
rect 23438 14530 23490 14542
rect 33070 14530 33122 14542
rect 40350 14530 40402 14542
rect 23874 14478 23886 14530
rect 23938 14478 23950 14530
rect 32498 14478 32510 14530
rect 32562 14478 32574 14530
rect 36306 14478 36318 14530
rect 36370 14478 36382 14530
rect 40002 14478 40014 14530
rect 40066 14478 40078 14530
rect 23438 14466 23490 14478
rect 33070 14466 33122 14478
rect 40350 14466 40402 14478
rect 21646 14418 21698 14430
rect 2370 14366 2382 14418
rect 2434 14366 2446 14418
rect 6066 14366 6078 14418
rect 6130 14366 6142 14418
rect 12450 14366 12462 14418
rect 12514 14366 12526 14418
rect 15922 14366 15934 14418
rect 15986 14366 15998 14418
rect 18498 14366 18510 14418
rect 18562 14366 18574 14418
rect 21646 14354 21698 14366
rect 30158 14418 30210 14430
rect 37662 14418 37714 14430
rect 35298 14366 35310 14418
rect 35362 14366 35374 14418
rect 42914 14366 42926 14418
rect 42978 14366 42990 14418
rect 30158 14354 30210 14366
rect 37662 14354 37714 14366
rect 26910 14306 26962 14318
rect 26338 14254 26350 14306
rect 26402 14254 26414 14306
rect 26910 14242 26962 14254
rect 29374 14306 29426 14318
rect 29374 14242 29426 14254
rect 36878 14306 36930 14318
rect 36878 14242 36930 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 5394 13918 5406 13970
rect 5458 13918 5470 13970
rect 8418 13806 8430 13858
rect 8482 13806 8494 13858
rect 12786 13806 12798 13858
rect 12850 13806 12862 13858
rect 15250 13806 15262 13858
rect 15314 13806 15326 13858
rect 20962 13806 20974 13858
rect 21026 13806 21038 13858
rect 21634 13806 21646 13858
rect 21698 13806 21710 13858
rect 29250 13806 29262 13858
rect 29314 13806 29326 13858
rect 31938 13806 31950 13858
rect 32002 13806 32014 13858
rect 35746 13806 35758 13858
rect 35810 13806 35822 13858
rect 38210 13806 38222 13858
rect 38274 13806 38286 13858
rect 2270 13746 2322 13758
rect 2930 13694 2942 13746
rect 2994 13694 3006 13746
rect 2270 13682 2322 13694
rect 7186 13582 7198 13634
rect 7250 13582 7262 13634
rect 11442 13582 11454 13634
rect 11506 13582 11518 13634
rect 14242 13582 14254 13634
rect 14306 13582 14318 13634
rect 19730 13582 19742 13634
rect 19794 13582 19806 13634
rect 22978 13582 22990 13634
rect 23042 13582 23054 13634
rect 28354 13582 28366 13634
rect 28418 13582 28430 13634
rect 30930 13582 30942 13634
rect 30994 13582 31006 13634
rect 34402 13582 34414 13634
rect 34466 13582 34478 13634
rect 37202 13582 37214 13634
rect 37266 13582 37278 13634
rect 5966 13522 6018 13534
rect 5966 13458 6018 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 26686 13074 26738 13086
rect 3602 13022 3614 13074
rect 3666 13022 3678 13074
rect 11554 13022 11566 13074
rect 11618 13022 11630 13074
rect 15250 13022 15262 13074
rect 15314 13022 15326 13074
rect 19058 13022 19070 13074
rect 19122 13022 19134 13074
rect 30146 13022 30158 13074
rect 30210 13022 30222 13074
rect 34290 13022 34302 13074
rect 34354 13022 34366 13074
rect 37986 13022 37998 13074
rect 38050 13022 38062 13074
rect 40786 13022 40798 13074
rect 40850 13022 40862 13074
rect 26686 13010 26738 13022
rect 26238 12962 26290 12974
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 26238 12898 26290 12910
rect 23326 12850 23378 12862
rect 4946 12798 4958 12850
rect 5010 12798 5022 12850
rect 12450 12798 12462 12850
rect 12514 12798 12526 12850
rect 16594 12798 16606 12850
rect 16658 12798 16670 12850
rect 17826 12798 17838 12850
rect 17890 12798 17902 12850
rect 31154 12798 31166 12850
rect 31218 12798 31230 12850
rect 35634 12798 35646 12850
rect 35698 12798 35710 12850
rect 38994 12798 39006 12850
rect 39058 12798 39070 12850
rect 42018 12798 42030 12850
rect 42082 12798 42094 12850
rect 23326 12786 23378 12798
rect 22542 12738 22594 12750
rect 22542 12674 22594 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 14242 12238 14254 12290
rect 14306 12238 14318 12290
rect 17490 12238 17502 12290
rect 17554 12238 17566 12290
rect 23538 12238 23550 12290
rect 23602 12238 23614 12290
rect 27234 12238 27246 12290
rect 27298 12238 27310 12290
rect 30370 12238 30382 12290
rect 30434 12238 30446 12290
rect 35410 12238 35422 12290
rect 35474 12238 35486 12290
rect 15362 12014 15374 12066
rect 15426 12014 15438 12066
rect 18722 12014 18734 12066
rect 18786 12014 18798 12066
rect 22306 12014 22318 12066
rect 22370 12014 22382 12066
rect 26226 12014 26238 12066
rect 26290 12014 26302 12066
rect 29026 12014 29038 12066
rect 29090 12014 29102 12066
rect 34066 12014 34078 12066
rect 34130 12014 34142 12066
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 24098 11454 24110 11506
rect 24162 11454 24174 11506
rect 26674 11454 26686 11506
rect 26738 11454 26750 11506
rect 33506 11454 33518 11506
rect 33570 11454 33582 11506
rect 22978 11230 22990 11282
rect 23042 11230 23054 11282
rect 28018 11230 28030 11282
rect 28082 11230 28094 11282
rect 34850 11230 34862 11282
rect 34914 11230 34926 11282
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 20078 9154 20130 9166
rect 20078 9090 20130 9102
rect 20862 9154 20914 9166
rect 20862 9090 20914 9102
rect 43822 9154 43874 9166
rect 43822 9090 43874 9102
rect 19742 9042 19794 9054
rect 44158 9042 44210 9054
rect 20626 8990 20638 9042
rect 20690 8990 20702 9042
rect 19742 8978 19794 8990
rect 44158 8978 44210 8990
rect 43598 8930 43650 8942
rect 43598 8866 43650 8878
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 27010 8206 27022 8258
rect 27074 8206 27086 8258
rect 42914 8206 42926 8258
rect 42978 8206 42990 8258
rect 44034 8094 44046 8146
rect 44098 8094 44110 8146
rect 27246 8034 27298 8046
rect 27246 7970 27298 7982
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 42590 7586 42642 7598
rect 42590 7522 42642 7534
rect 44046 7474 44098 7486
rect 42914 7422 42926 7474
rect 42978 7422 42990 7474
rect 44046 7410 44098 7422
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 43138 6638 43150 6690
rect 43202 6638 43214 6690
rect 24446 6578 24498 6590
rect 44034 6526 44046 6578
rect 44098 6526 44110 6578
rect 24446 6514 24498 6526
rect 24782 6466 24834 6478
rect 24782 6402 24834 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 42914 5854 42926 5906
rect 42978 5854 42990 5906
rect 42254 5794 42306 5806
rect 42254 5730 42306 5742
rect 42702 5794 42754 5806
rect 44034 5742 44046 5794
rect 44098 5742 44110 5794
rect 42702 5730 42754 5742
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 43822 5122 43874 5134
rect 25106 5070 25118 5122
rect 25170 5070 25182 5122
rect 33394 5070 33406 5122
rect 33458 5070 33470 5122
rect 37426 5070 37438 5122
rect 37490 5070 37502 5122
rect 38098 5070 38110 5122
rect 38162 5070 38174 5122
rect 38658 5070 38670 5122
rect 38722 5070 38734 5122
rect 43822 5058 43874 5070
rect 31838 5010 31890 5022
rect 31838 4946 31890 4958
rect 37886 5010 37938 5022
rect 37886 4946 37938 4958
rect 39230 5010 39282 5022
rect 39230 4946 39282 4958
rect 41470 5010 41522 5022
rect 41470 4946 41522 4958
rect 41806 5010 41858 5022
rect 41806 4946 41858 4958
rect 42142 5010 42194 5022
rect 42142 4946 42194 4958
rect 42478 5010 42530 5022
rect 42478 4946 42530 4958
rect 42814 5010 42866 5022
rect 42814 4946 42866 4958
rect 43150 5010 43202 5022
rect 43150 4946 43202 4958
rect 43486 5010 43538 5022
rect 43486 4946 43538 4958
rect 25342 4898 25394 4910
rect 25342 4834 25394 4846
rect 32174 4898 32226 4910
rect 32174 4834 32226 4846
rect 33630 4898 33682 4910
rect 33630 4834 33682 4846
rect 35870 4898 35922 4910
rect 35870 4834 35922 4846
rect 36542 4898 36594 4910
rect 36542 4834 36594 4846
rect 37214 4898 37266 4910
rect 37214 4834 37266 4846
rect 38894 4898 38946 4910
rect 38894 4834 38946 4846
rect 39566 4898 39618 4910
rect 39566 4834 39618 4846
rect 40686 4898 40738 4910
rect 40686 4834 40738 4846
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 20078 4562 20130 4574
rect 20078 4498 20130 4510
rect 20750 4562 20802 4574
rect 20750 4498 20802 4510
rect 25230 4562 25282 4574
rect 25230 4498 25282 4510
rect 27134 4562 27186 4574
rect 27134 4498 27186 4510
rect 33518 4562 33570 4574
rect 33518 4498 33570 4510
rect 35758 4562 35810 4574
rect 35758 4498 35810 4510
rect 36430 4562 36482 4574
rect 36430 4498 36482 4510
rect 37102 4562 37154 4574
rect 37102 4498 37154 4510
rect 38894 4562 38946 4574
rect 38894 4498 38946 4510
rect 40910 4562 40962 4574
rect 40910 4498 40962 4510
rect 42814 4562 42866 4574
rect 42814 4498 42866 4510
rect 43822 4562 43874 4574
rect 43822 4498 43874 4510
rect 19070 4450 19122 4462
rect 19070 4386 19122 4398
rect 26462 4450 26514 4462
rect 26462 4386 26514 4398
rect 32398 4450 32450 4462
rect 32398 4386 32450 4398
rect 38222 4450 38274 4462
rect 38222 4386 38274 4398
rect 39902 4450 39954 4462
rect 39902 4386 39954 4398
rect 41582 4450 41634 4462
rect 41582 4386 41634 4398
rect 42366 4450 42418 4462
rect 42366 4386 42418 4398
rect 43150 4450 43202 4462
rect 43150 4386 43202 4398
rect 19742 4338 19794 4350
rect 19742 4274 19794 4286
rect 20414 4338 20466 4350
rect 20414 4274 20466 4286
rect 25566 4338 25618 4350
rect 33182 4338 33234 4350
rect 27346 4286 27358 4338
rect 27410 4286 27422 4338
rect 25566 4274 25618 4286
rect 33182 4274 33234 4286
rect 36094 4338 36146 4350
rect 36094 4274 36146 4286
rect 36766 4338 36818 4350
rect 38558 4338 38610 4350
rect 37986 4286 37998 4338
rect 38050 4286 38062 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 41794 4286 41806 4338
rect 41858 4286 41870 4338
rect 43362 4286 43374 4338
rect 43426 4286 43438 4338
rect 44034 4286 44046 4338
rect 44098 4286 44110 4338
rect 36766 4274 36818 4286
rect 38558 4274 38610 4286
rect 19518 4226 19570 4238
rect 19518 4162 19570 4174
rect 24222 4226 24274 4238
rect 24222 4162 24274 4174
rect 24782 4226 24834 4238
rect 24782 4162 24834 4174
rect 26238 4226 26290 4238
rect 26238 4162 26290 4174
rect 32174 4226 32226 4238
rect 32174 4162 32226 4174
rect 37662 4226 37714 4238
rect 37662 4162 37714 4174
rect 34974 4114 35026 4126
rect 34974 4050 35026 4062
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 21522 3614 21534 3666
rect 21586 3614 21598 3666
rect 26562 3614 26574 3666
rect 26626 3614 26638 3666
rect 28802 3614 28814 3666
rect 28866 3614 28878 3666
rect 32610 3614 32622 3666
rect 32674 3614 32686 3666
rect 34290 3614 34302 3666
rect 34354 3614 34366 3666
rect 40226 3614 40238 3666
rect 40290 3614 40302 3666
rect 42242 3614 42254 3666
rect 42306 3614 42318 3666
rect 21086 3554 21138 3566
rect 26126 3554 26178 3566
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 23762 3502 23774 3554
rect 23826 3502 23838 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 21086 3490 21138 3502
rect 26126 3490 26178 3502
rect 28366 3554 28418 3566
rect 28366 3490 28418 3502
rect 32174 3554 32226 3566
rect 32174 3490 32226 3502
rect 33854 3554 33906 3566
rect 33854 3490 33906 3502
rect 37214 3554 37266 3566
rect 39790 3554 39842 3566
rect 39106 3502 39118 3554
rect 39170 3502 39182 3554
rect 37214 3490 37266 3502
rect 39790 3490 39842 3502
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 30942 3442 30994 3454
rect 30942 3378 30994 3390
rect 31166 3442 31218 3454
rect 31166 3378 31218 3390
rect 31502 3442 31554 3454
rect 31502 3378 31554 3390
rect 41246 3442 41298 3454
rect 41246 3378 41298 3390
rect 41806 3442 41858 3454
rect 41806 3378 41858 3390
rect 43150 3442 43202 3454
rect 43150 3378 43202 3390
rect 43822 3442 43874 3454
rect 43822 3378 43874 3390
rect 44158 3442 44210 3454
rect 44158 3378 44210 3390
rect 19406 3330 19458 3342
rect 19406 3266 19458 3278
rect 22654 3330 22706 3342
rect 22654 3266 22706 3278
rect 24558 3330 24610 3342
rect 24558 3266 24610 3278
rect 36430 3330 36482 3342
rect 36430 3266 36482 3278
rect 37550 3330 37602 3342
rect 37550 3266 37602 3278
rect 38446 3330 38498 3342
rect 38446 3266 38498 3278
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 15598 42142 15650 42194
rect 19406 42142 19458 42194
rect 31166 42142 31218 42194
rect 33182 42142 33234 42194
rect 34750 42142 34802 42194
rect 36654 42142 36706 42194
rect 38446 42142 38498 42194
rect 41358 42142 41410 42194
rect 14142 42030 14194 42082
rect 14814 42030 14866 42082
rect 28366 42030 28418 42082
rect 32846 42030 32898 42082
rect 36318 42030 36370 42082
rect 37550 42030 37602 42082
rect 43822 42030 43874 42082
rect 13918 41918 13970 41970
rect 14590 41918 14642 41970
rect 15262 41918 15314 41970
rect 16270 41918 16322 41970
rect 16942 41918 16994 41970
rect 20078 41918 20130 41970
rect 20862 41918 20914 41970
rect 22430 41918 22482 41970
rect 24558 41918 24610 41970
rect 26462 41918 26514 41970
rect 27918 41918 27970 41970
rect 28590 41918 28642 41970
rect 32510 41918 32562 41970
rect 33854 41918 33906 41970
rect 35534 41918 35586 41970
rect 35982 41918 36034 41970
rect 37214 41918 37266 41970
rect 39230 41918 39282 41970
rect 39790 41918 39842 41970
rect 41806 41918 41858 41970
rect 44158 41918 44210 41970
rect 17390 41806 17442 41858
rect 21310 41806 21362 41858
rect 22878 41806 22930 41858
rect 25006 41806 25058 41858
rect 26910 41806 26962 41858
rect 40350 41806 40402 41858
rect 42366 41806 42418 41858
rect 43150 41806 43202 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 14366 41246 14418 41298
rect 19294 41246 19346 41298
rect 20190 41246 20242 41298
rect 21534 41246 21586 41298
rect 23550 41246 23602 41298
rect 24894 41246 24946 41298
rect 27582 41246 27634 41298
rect 32510 41246 32562 41298
rect 37214 41246 37266 41298
rect 37662 41246 37714 41298
rect 40350 41246 40402 41298
rect 42030 41246 42082 41298
rect 44046 41246 44098 41298
rect 17726 41134 17778 41186
rect 20414 41134 20466 41186
rect 21982 41134 22034 41186
rect 23774 41134 23826 41186
rect 26014 41134 26066 41186
rect 37886 41134 37938 41186
rect 42478 41134 42530 41186
rect 42926 41134 42978 41186
rect 17054 41022 17106 41074
rect 25118 41022 25170 41074
rect 31838 41022 31890 41074
rect 16830 40910 16882 40962
rect 18062 40910 18114 40962
rect 18846 40910 18898 40962
rect 20750 40910 20802 40962
rect 21758 40910 21810 40962
rect 24110 40910 24162 40962
rect 25790 40910 25842 40962
rect 27134 40910 27186 40962
rect 38222 40910 38274 40962
rect 39566 40910 39618 40962
rect 39902 40910 39954 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 15150 40574 15202 40626
rect 15822 40574 15874 40626
rect 18846 40574 18898 40626
rect 19742 40574 19794 40626
rect 33406 40574 33458 40626
rect 39454 40574 39506 40626
rect 42590 40574 42642 40626
rect 43710 40574 43762 40626
rect 44158 40574 44210 40626
rect 14814 40462 14866 40514
rect 15486 40462 15538 40514
rect 18510 40462 18562 40514
rect 20078 40462 20130 40514
rect 33070 40462 33122 40514
rect 38782 40462 38834 40514
rect 39118 40462 39170 40514
rect 39790 40462 39842 40514
rect 40350 40462 40402 40514
rect 40910 40462 40962 40514
rect 41918 40462 41970 40514
rect 42926 40462 42978 40514
rect 19518 40350 19570 40402
rect 20302 40350 20354 40402
rect 41134 40350 41186 40402
rect 41694 40350 41746 40402
rect 42366 40350 42418 40402
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 44158 39790 44210 39842
rect 19854 39678 19906 39730
rect 40686 39678 40738 39730
rect 39118 39566 39170 39618
rect 39902 39566 39954 39618
rect 41806 39566 41858 39618
rect 39454 39454 39506 39506
rect 40126 39454 40178 39506
rect 41470 39454 41522 39506
rect 42142 39454 42194 39506
rect 42478 39454 42530 39506
rect 42814 39454 42866 39506
rect 43374 39342 43426 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 42366 39006 42418 39058
rect 43150 39006 43202 39058
rect 43822 39006 43874 39058
rect 42814 38894 42866 38946
rect 43486 38894 43538 38946
rect 44046 38782 44098 38834
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 43150 38110 43202 38162
rect 44046 37998 44098 38050
rect 43822 37886 43874 37938
rect 43486 37774 43538 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 43822 37438 43874 37490
rect 44158 37326 44210 37378
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 43710 36318 43762 36370
rect 44158 36206 44210 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 20750 35870 20802 35922
rect 21646 35870 21698 35922
rect 24446 35870 24498 35922
rect 25790 35870 25842 35922
rect 26462 35870 26514 35922
rect 24110 35758 24162 35810
rect 44158 35758 44210 35810
rect 20526 35646 20578 35698
rect 21422 35646 21474 35698
rect 25566 35646 25618 35698
rect 26238 35646 26290 35698
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 11454 31838 11506 31890
rect 18510 31838 18562 31890
rect 22318 31838 22370 31890
rect 42926 31726 42978 31778
rect 12462 31614 12514 31666
rect 17390 31614 17442 31666
rect 23550 31614 23602 31666
rect 44046 31614 44098 31666
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 42702 31166 42754 31218
rect 14142 31054 14194 31106
rect 22542 31054 22594 31106
rect 28702 31054 28754 31106
rect 31502 31054 31554 31106
rect 34638 31054 34690 31106
rect 43822 31054 43874 31106
rect 19630 30942 19682 30994
rect 20302 30942 20354 30994
rect 42478 30942 42530 30994
rect 43598 30942 43650 30994
rect 44158 30942 44210 30994
rect 12910 30830 12962 30882
rect 27806 30830 27858 30882
rect 30494 30830 30546 30882
rect 35982 30830 36034 30882
rect 23326 30718 23378 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 6638 30270 6690 30322
rect 11230 30270 11282 30322
rect 19182 30270 19234 30322
rect 23102 30270 23154 30322
rect 25902 30270 25954 30322
rect 31054 30270 31106 30322
rect 33854 30270 33906 30322
rect 37998 30270 38050 30322
rect 14478 30158 14530 30210
rect 14926 30158 14978 30210
rect 7646 30046 7698 30098
rect 9886 30046 9938 30098
rect 17950 30046 18002 30098
rect 20190 30046 20242 30098
rect 21310 30046 21362 30098
rect 21646 30046 21698 30098
rect 24110 30046 24162 30098
rect 26910 30046 26962 30098
rect 27694 30046 27746 30098
rect 28030 30046 28082 30098
rect 29486 30046 29538 30098
rect 32062 30046 32114 30098
rect 34862 30046 34914 30098
rect 35646 30046 35698 30098
rect 39006 30046 39058 30098
rect 17166 29934 17218 29986
rect 29374 29934 29426 29986
rect 35758 29934 35810 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5294 29598 5346 29650
rect 20414 29598 20466 29650
rect 20974 29598 21026 29650
rect 24222 29598 24274 29650
rect 24782 29598 24834 29650
rect 25342 29598 25394 29650
rect 29374 29598 29426 29650
rect 4510 29486 4562 29538
rect 8542 29486 8594 29538
rect 13582 29486 13634 29538
rect 16382 29486 16434 29538
rect 25230 29486 25282 29538
rect 35310 29486 35362 29538
rect 37886 29486 37938 29538
rect 1822 29374 1874 29426
rect 2158 29374 2210 29426
rect 17502 29374 17554 29426
rect 17950 29374 18002 29426
rect 21310 29374 21362 29426
rect 21758 29374 21810 29426
rect 26238 29374 26290 29426
rect 26910 29374 26962 29426
rect 7534 29262 7586 29314
rect 12574 29262 12626 29314
rect 15374 29262 15426 29314
rect 31502 29262 31554 29314
rect 31838 29262 31890 29314
rect 34078 29262 34130 29314
rect 36878 29262 36930 29314
rect 29934 29150 29986 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 11566 28814 11618 28866
rect 16270 28814 16322 28866
rect 27694 28814 27746 28866
rect 32734 28814 32786 28866
rect 36542 28814 36594 28866
rect 4958 28702 5010 28754
rect 15038 28702 15090 28754
rect 20638 28702 20690 28754
rect 22318 28702 22370 28754
rect 41806 28702 41858 28754
rect 4846 28590 4898 28642
rect 5742 28590 5794 28642
rect 6750 28590 6802 28642
rect 7422 28590 7474 28642
rect 7870 28590 7922 28642
rect 8430 28590 8482 28642
rect 19406 28590 19458 28642
rect 19742 28590 19794 28642
rect 20526 28590 20578 28642
rect 23998 28590 24050 28642
rect 24670 28590 24722 28642
rect 29038 28590 29090 28642
rect 29710 28590 29762 28642
rect 33070 28590 33122 28642
rect 33518 28590 33570 28642
rect 36990 28590 37042 28642
rect 37550 28590 37602 28642
rect 6974 28478 7026 28530
rect 13694 28478 13746 28530
rect 23550 28478 23602 28530
rect 27918 28478 27970 28530
rect 31950 28478 32002 28530
rect 35758 28478 35810 28530
rect 42814 28478 42866 28530
rect 10782 28366 10834 28418
rect 17054 28366 17106 28418
rect 27134 28366 27186 28418
rect 28030 28366 28082 28418
rect 40014 28366 40066 28418
rect 40574 28366 40626 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 2046 28030 2098 28082
rect 3054 28030 3106 28082
rect 10782 28030 10834 28082
rect 15262 28030 15314 28082
rect 16718 28030 16770 28082
rect 28030 28030 28082 28082
rect 32622 28030 32674 28082
rect 6638 27918 6690 27970
rect 14478 27918 14530 27970
rect 18846 27918 18898 27970
rect 23998 27918 24050 27970
rect 31838 27918 31890 27970
rect 33742 27918 33794 27970
rect 39678 27918 39730 27970
rect 40462 27918 40514 27970
rect 42926 27918 42978 27970
rect 1710 27806 1762 27858
rect 5294 27806 5346 27858
rect 5742 27806 5794 27858
rect 10782 27806 10834 27858
rect 11566 27806 11618 27858
rect 12238 27806 12290 27858
rect 21310 27806 21362 27858
rect 21758 27806 21810 27858
rect 25118 27806 25170 27858
rect 25790 27806 25842 27858
rect 29038 27806 29090 27858
rect 29486 27806 29538 27858
rect 35982 27806 36034 27858
rect 36654 27806 36706 27858
rect 36990 27806 37042 27858
rect 37438 27806 37490 27858
rect 7982 27694 8034 27746
rect 9550 27694 9602 27746
rect 9886 27694 9938 27746
rect 15710 27694 15762 27746
rect 16830 27694 16882 27746
rect 17726 27694 17778 27746
rect 18062 27694 18114 27746
rect 19854 27694 19906 27746
rect 20974 27694 21026 27746
rect 41918 27694 41970 27746
rect 2270 27582 2322 27634
rect 24782 27582 24834 27634
rect 28814 27582 28866 27634
rect 32958 27582 33010 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 9214 27246 9266 27298
rect 13022 27246 13074 27298
rect 22094 27246 22146 27298
rect 27358 27246 27410 27298
rect 34190 27246 34242 27298
rect 40574 27246 40626 27298
rect 1822 27134 1874 27186
rect 4062 27134 4114 27186
rect 14142 27134 14194 27186
rect 19406 27134 19458 27186
rect 23438 27134 23490 27186
rect 35534 27134 35586 27186
rect 41806 27134 41858 27186
rect 5518 27022 5570 27074
rect 6190 27022 6242 27074
rect 9326 27022 9378 27074
rect 9998 27022 10050 27074
rect 13918 27022 13970 27074
rect 15934 27022 15986 27074
rect 16382 27022 16434 27074
rect 19854 27022 19906 27074
rect 20638 27022 20690 27074
rect 23886 27022 23938 27074
rect 24334 27022 24386 27074
rect 30494 27022 30546 27074
rect 31166 27022 31218 27074
rect 34862 27022 34914 27074
rect 37102 27022 37154 27074
rect 37550 27022 37602 27074
rect 2718 26910 2770 26962
rect 12238 26910 12290 26962
rect 14478 26910 14530 26962
rect 14814 26910 14866 26962
rect 18622 26910 18674 26962
rect 19630 26910 19682 26962
rect 20414 26910 20466 26962
rect 21534 26910 21586 26962
rect 23102 26910 23154 26962
rect 26574 26910 26626 26962
rect 27582 26910 27634 26962
rect 27918 26910 27970 26962
rect 29262 26910 29314 26962
rect 36318 26910 36370 26962
rect 42814 26910 42866 26962
rect 43598 26910 43650 26962
rect 43934 26910 43986 26962
rect 8654 26798 8706 26850
rect 15486 26798 15538 26850
rect 29374 26798 29426 26850
rect 33406 26798 33458 26850
rect 40014 26798 40066 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 6974 26462 7026 26514
rect 7646 26462 7698 26514
rect 33406 26462 33458 26514
rect 36878 26462 36930 26514
rect 43822 26462 43874 26514
rect 3054 26350 3106 26402
rect 8654 26350 8706 26402
rect 9774 26350 9826 26402
rect 28590 26350 28642 26402
rect 37550 26350 37602 26402
rect 39790 26350 39842 26402
rect 42926 26350 42978 26402
rect 2494 26238 2546 26290
rect 2830 26238 2882 26290
rect 3950 26238 4002 26290
rect 4510 26238 4562 26290
rect 8878 26238 8930 26290
rect 14814 26238 14866 26290
rect 16718 26238 16770 26290
rect 21870 26238 21922 26290
rect 23214 26238 23266 26290
rect 32174 26238 32226 26290
rect 33406 26238 33458 26290
rect 34078 26238 34130 26290
rect 34526 26238 34578 26290
rect 3390 26126 3442 26178
rect 3726 26126 3778 26178
rect 8318 26126 8370 26178
rect 15150 26126 15202 26178
rect 15486 26126 15538 26178
rect 15822 26126 15874 26178
rect 16158 26126 16210 26178
rect 16494 26126 16546 26178
rect 19630 26126 19682 26178
rect 22990 26126 23042 26178
rect 23774 26126 23826 26178
rect 26798 26126 26850 26178
rect 38894 26126 38946 26178
rect 41918 26126 41970 26178
rect 43710 26126 43762 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 5518 25678 5570 25730
rect 19854 25678 19906 25730
rect 3838 25566 3890 25618
rect 4510 25566 4562 25618
rect 14926 25566 14978 25618
rect 20302 25566 20354 25618
rect 20526 25566 20578 25618
rect 22878 25566 22930 25618
rect 25678 25566 25730 25618
rect 30158 25566 30210 25618
rect 32958 25566 33010 25618
rect 35646 25566 35698 25618
rect 36430 25566 36482 25618
rect 36990 25566 37042 25618
rect 42478 25566 42530 25618
rect 8654 25454 8706 25506
rect 9214 25454 9266 25506
rect 12350 25454 12402 25506
rect 12798 25454 12850 25506
rect 16270 25454 16322 25506
rect 16830 25454 16882 25506
rect 34862 25454 34914 25506
rect 37550 25454 37602 25506
rect 38222 25454 38274 25506
rect 2718 25342 2770 25394
rect 6302 25342 6354 25394
rect 13582 25342 13634 25394
rect 19070 25342 19122 25394
rect 23886 25342 23938 25394
rect 26910 25342 26962 25394
rect 31502 25342 31554 25394
rect 33966 25342 34018 25394
rect 41246 25342 41298 25394
rect 43710 25342 43762 25394
rect 9326 25230 9378 25282
rect 10110 25230 10162 25282
rect 15486 25230 15538 25282
rect 15934 25230 15986 25282
rect 32174 25230 32226 25282
rect 32734 25230 32786 25282
rect 37102 25230 37154 25282
rect 40686 25230 40738 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2046 24894 2098 24946
rect 2830 24894 2882 24946
rect 12574 24894 12626 24946
rect 13134 24894 13186 24946
rect 13246 24894 13298 24946
rect 14030 24894 14082 24946
rect 22766 24894 22818 24946
rect 23326 24894 23378 24946
rect 29374 24894 29426 24946
rect 6974 24782 7026 24834
rect 31390 24782 31442 24834
rect 31726 24782 31778 24834
rect 39342 24782 39394 24834
rect 40014 24782 40066 24834
rect 43150 24782 43202 24834
rect 5182 24670 5234 24722
rect 5630 24670 5682 24722
rect 9438 24670 9490 24722
rect 10110 24670 10162 24722
rect 16270 24670 16322 24722
rect 16942 24670 16994 24722
rect 18398 24670 18450 24722
rect 19854 24670 19906 24722
rect 20302 24670 20354 24722
rect 26462 24670 26514 24722
rect 27022 24670 27074 24722
rect 31054 24670 31106 24722
rect 32286 24670 32338 24722
rect 33630 24670 33682 24722
rect 39678 24670 39730 24722
rect 7982 24558 8034 24610
rect 19070 24558 19122 24610
rect 19406 24558 19458 24610
rect 23550 24558 23602 24610
rect 23886 24558 23938 24610
rect 30158 24558 30210 24610
rect 32510 24558 32562 24610
rect 35646 24558 35698 24610
rect 39006 24558 39058 24610
rect 41918 24558 41970 24610
rect 17614 24446 17666 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 11902 24110 11954 24162
rect 17166 24110 17218 24162
rect 4062 23998 4114 24050
rect 6750 23998 6802 24050
rect 11006 23998 11058 24050
rect 13470 23998 13522 24050
rect 15934 23998 15986 24050
rect 16382 23998 16434 24050
rect 23326 23998 23378 24050
rect 24334 23998 24386 24050
rect 36990 23998 37042 24050
rect 43486 23998 43538 24050
rect 9998 23886 10050 23938
rect 10446 23886 10498 23938
rect 13694 23886 13746 23938
rect 20190 23886 20242 23938
rect 20862 23886 20914 23938
rect 24558 23886 24610 23938
rect 25230 23886 25282 23938
rect 29038 23886 29090 23938
rect 29710 23886 29762 23938
rect 32846 23886 32898 23938
rect 33518 23886 33570 23938
rect 37214 23886 37266 23938
rect 38110 23886 38162 23938
rect 38782 23886 38834 23938
rect 42254 23886 42306 23938
rect 3054 23774 3106 23826
rect 6414 23774 6466 23826
rect 11342 23774 11394 23826
rect 12910 23774 12962 23826
rect 14926 23774 14978 23826
rect 17950 23774 18002 23826
rect 22318 23774 22370 23826
rect 42030 23774 42082 23826
rect 6974 23662 7026 23714
rect 7646 23662 7698 23714
rect 16942 23662 16994 23714
rect 27694 23662 27746 23714
rect 28254 23662 28306 23714
rect 32174 23662 32226 23714
rect 32734 23662 32786 23714
rect 35982 23662 36034 23714
rect 36542 23662 36594 23714
rect 41246 23662 41298 23714
rect 41806 23662 41858 23714
rect 42926 23662 42978 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 16158 23326 16210 23378
rect 16942 23326 16994 23378
rect 23438 23326 23490 23378
rect 29934 23326 29986 23378
rect 32958 23326 33010 23378
rect 33518 23326 33570 23378
rect 4062 23214 4114 23266
rect 6974 23214 7026 23266
rect 9438 23214 9490 23266
rect 10222 23214 10274 23266
rect 18062 23214 18114 23266
rect 31502 23214 31554 23266
rect 32174 23214 32226 23266
rect 39678 23214 39730 23266
rect 42926 23214 42978 23266
rect 43710 23214 43762 23266
rect 12462 23102 12514 23154
rect 13134 23102 13186 23154
rect 13358 23102 13410 23154
rect 13806 23102 13858 23154
rect 20302 23102 20354 23154
rect 20862 23102 20914 23154
rect 24558 23102 24610 23154
rect 26238 23102 26290 23154
rect 27134 23102 27186 23154
rect 27582 23102 27634 23154
rect 31726 23102 31778 23154
rect 36094 23102 36146 23154
rect 36430 23102 36482 23154
rect 36766 23102 36818 23154
rect 37438 23102 37490 23154
rect 5182 22990 5234 23042
rect 7982 22990 8034 23042
rect 19070 22990 19122 23042
rect 24334 22990 24386 23042
rect 25454 22990 25506 23042
rect 30830 22990 30882 23042
rect 31166 22990 31218 23042
rect 32510 22990 32562 23042
rect 41918 22990 41970 23042
rect 43934 22990 43986 23042
rect 23998 22878 24050 22930
rect 30606 22878 30658 22930
rect 40462 22878 40514 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 9214 22542 9266 22594
rect 33518 22542 33570 22594
rect 4062 22430 4114 22482
rect 13582 22430 13634 22482
rect 15374 22430 15426 22482
rect 15822 22430 15874 22482
rect 27918 22430 27970 22482
rect 28142 22430 28194 22482
rect 28478 22430 28530 22482
rect 34750 22430 34802 22482
rect 41806 22430 41858 22482
rect 5518 22318 5570 22370
rect 6078 22318 6130 22370
rect 9326 22318 9378 22370
rect 9886 22318 9938 22370
rect 19742 22318 19794 22370
rect 20302 22318 20354 22370
rect 21422 22318 21474 22370
rect 29374 22318 29426 22370
rect 30046 22318 30098 22370
rect 30494 22318 30546 22370
rect 36878 22318 36930 22370
rect 37550 22318 37602 22370
rect 3054 22206 3106 22258
rect 14366 22206 14418 22258
rect 16606 22206 16658 22258
rect 23550 22206 23602 22258
rect 29598 22206 29650 22258
rect 35758 22206 35810 22258
rect 42814 22206 42866 22258
rect 43598 22206 43650 22258
rect 8654 22094 8706 22146
rect 12350 22094 12402 22146
rect 13022 22094 13074 22146
rect 17390 22094 17442 22146
rect 20862 22094 20914 22146
rect 32958 22094 33010 22146
rect 33854 22094 33906 22146
rect 34302 22094 34354 22146
rect 40014 22094 40066 22146
rect 40574 22094 40626 22146
rect 41470 22094 41522 22146
rect 43710 22094 43762 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2158 21758 2210 21810
rect 6190 21758 6242 21810
rect 12574 21758 12626 21810
rect 16382 21758 16434 21810
rect 16942 21758 16994 21810
rect 21310 21758 21362 21810
rect 21982 21758 22034 21810
rect 28926 21758 28978 21810
rect 29822 21758 29874 21810
rect 37326 21758 37378 21810
rect 11006 21646 11058 21698
rect 22654 21646 22706 21698
rect 31950 21646 32002 21698
rect 33070 21646 33122 21698
rect 38446 21646 38498 21698
rect 39454 21646 39506 21698
rect 42926 21646 42978 21698
rect 4734 21534 4786 21586
rect 5294 21534 5346 21586
rect 8430 21534 8482 21586
rect 9102 21534 9154 21586
rect 9998 21534 10050 21586
rect 13358 21534 13410 21586
rect 13806 21534 13858 21586
rect 18398 21534 18450 21586
rect 18846 21534 18898 21586
rect 25342 21534 25394 21586
rect 25790 21534 25842 21586
rect 26462 21534 26514 21586
rect 33406 21534 33458 21586
rect 33854 21534 33906 21586
rect 34190 21534 34242 21586
rect 34862 21534 34914 21586
rect 38110 21534 38162 21586
rect 43710 21534 43762 21586
rect 10222 21422 10274 21474
rect 12014 21422 12066 21474
rect 23662 21422 23714 21474
rect 25566 21422 25618 21474
rect 30718 21422 30770 21474
rect 38782 21422 38834 21474
rect 39118 21422 39170 21474
rect 39678 21422 39730 21474
rect 41918 21422 41970 21474
rect 43934 21422 43986 21474
rect 1598 21310 1650 21362
rect 5406 21310 5458 21362
rect 29486 21310 29538 21362
rect 37886 21310 37938 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 13358 20974 13410 21026
rect 22318 20974 22370 21026
rect 35758 20974 35810 21026
rect 4062 20862 4114 20914
rect 7646 20862 7698 20914
rect 11902 20862 11954 20914
rect 12574 20862 12626 20914
rect 21870 20862 21922 20914
rect 22094 20862 22146 20914
rect 29374 20862 29426 20914
rect 30158 20862 30210 20914
rect 33182 20862 33234 20914
rect 36430 20862 36482 20914
rect 36990 20862 37042 20914
rect 37326 20862 37378 20914
rect 42478 20862 42530 20914
rect 42702 20862 42754 20914
rect 7982 20750 8034 20802
rect 8542 20750 8594 20802
rect 12126 20750 12178 20802
rect 12798 20750 12850 20802
rect 16382 20750 16434 20802
rect 17054 20750 17106 20802
rect 17390 20750 17442 20802
rect 17726 20750 17778 20802
rect 25342 20750 25394 20802
rect 25790 20750 25842 20802
rect 28366 20750 28418 20802
rect 34750 20750 34802 20802
rect 37774 20750 37826 20802
rect 38446 20750 38498 20802
rect 3054 20638 3106 20690
rect 5630 20638 5682 20690
rect 5966 20638 6018 20690
rect 7422 20638 7474 20690
rect 10894 20638 10946 20690
rect 23102 20638 23154 20690
rect 31166 20638 31218 20690
rect 33966 20638 34018 20690
rect 43710 20638 43762 20690
rect 11678 20526 11730 20578
rect 13918 20526 13970 20578
rect 20302 20526 20354 20578
rect 20862 20526 20914 20578
rect 28366 20526 28418 20578
rect 40910 20526 40962 20578
rect 41470 20526 41522 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 21870 20190 21922 20242
rect 3278 20078 3330 20130
rect 6750 20078 6802 20130
rect 8654 20078 8706 20130
rect 8990 20078 9042 20130
rect 9774 20078 9826 20130
rect 20190 20078 20242 20130
rect 28814 20078 28866 20130
rect 31950 20078 32002 20130
rect 36206 20078 36258 20130
rect 39230 20078 39282 20130
rect 42926 20078 42978 20130
rect 4062 19966 4114 20018
rect 4398 19966 4450 20018
rect 14814 19966 14866 20018
rect 16158 19966 16210 20018
rect 17502 19966 17554 20018
rect 17950 19966 18002 20018
rect 24110 19966 24162 20018
rect 24558 19966 24610 20018
rect 25454 19966 25506 20018
rect 26014 19966 26066 20018
rect 26462 19966 26514 20018
rect 33518 19966 33570 20018
rect 33966 19966 34018 20018
rect 3614 19854 3666 19906
rect 7982 19854 8034 19906
rect 8318 19854 8370 19906
rect 16830 19854 16882 19906
rect 25230 19854 25282 19906
rect 30046 19854 30098 19906
rect 30494 19854 30546 19906
rect 30830 19854 30882 19906
rect 37326 19854 37378 19906
rect 38222 19854 38274 19906
rect 41918 19854 41970 19906
rect 7534 19742 7586 19794
rect 15822 19742 15874 19794
rect 20974 19742 21026 19794
rect 21086 19742 21138 19794
rect 29598 19742 29650 19794
rect 36990 19742 37042 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 12462 19406 12514 19458
rect 42814 19406 42866 19458
rect 3950 19294 4002 19346
rect 6302 19294 6354 19346
rect 6974 19294 7026 19346
rect 19966 19294 20018 19346
rect 21310 19294 21362 19346
rect 21646 19294 21698 19346
rect 22094 19294 22146 19346
rect 37886 19294 37938 19346
rect 6078 19182 6130 19234
rect 7198 19182 7250 19234
rect 7758 19182 7810 19234
rect 15038 19182 15090 19234
rect 20302 19182 20354 19234
rect 22430 19182 22482 19234
rect 23886 19182 23938 19234
rect 24334 19182 24386 19234
rect 32174 19182 32226 19234
rect 32734 19182 32786 19234
rect 35982 19182 36034 19234
rect 36542 19182 36594 19234
rect 37214 19182 37266 19234
rect 39118 19182 39170 19234
rect 39790 19182 39842 19234
rect 2046 19070 2098 19122
rect 3054 19070 3106 19122
rect 6638 19070 6690 19122
rect 10110 19070 10162 19122
rect 11454 19070 11506 19122
rect 13470 19070 13522 19122
rect 13806 19070 13858 19122
rect 18398 19070 18450 19122
rect 26574 19070 26626 19122
rect 28254 19070 28306 19122
rect 33630 19070 33682 19122
rect 38894 19070 38946 19122
rect 1710 18958 1762 19010
rect 10894 18958 10946 19010
rect 20750 18958 20802 19010
rect 27358 18958 27410 19010
rect 27694 18958 27746 19010
rect 28366 18958 28418 19010
rect 29038 18958 29090 19010
rect 29710 18958 29762 19010
rect 32846 18958 32898 19010
rect 38782 18958 38834 19010
rect 42254 18958 42306 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 1822 18622 1874 18674
rect 4958 18622 5010 18674
rect 15598 18622 15650 18674
rect 20526 18622 20578 18674
rect 6974 18510 7026 18562
rect 9998 18510 10050 18562
rect 21646 18510 21698 18562
rect 24558 18510 24610 18562
rect 30046 18510 30098 18562
rect 42926 18510 42978 18562
rect 2270 18398 2322 18450
rect 2718 18398 2770 18450
rect 12686 18398 12738 18450
rect 13022 18398 13074 18450
rect 17614 18398 17666 18450
rect 18062 18398 18114 18450
rect 26462 18398 26514 18450
rect 32062 18398 32114 18450
rect 32510 18398 32562 18450
rect 33070 18398 33122 18450
rect 38782 18398 38834 18450
rect 39342 18398 39394 18450
rect 39566 18398 39618 18450
rect 40238 18398 40290 18450
rect 7982 18286 8034 18338
rect 11230 18286 11282 18338
rect 16494 18286 16546 18338
rect 16830 18286 16882 18338
rect 21422 18286 21474 18338
rect 22094 18286 22146 18338
rect 23214 18286 23266 18338
rect 25342 18286 25394 18338
rect 26014 18286 26066 18338
rect 36542 18286 36594 18338
rect 39006 18286 39058 18338
rect 40014 18286 40066 18338
rect 41918 18286 41970 18338
rect 5742 18174 5794 18226
rect 16158 18174 16210 18226
rect 21086 18174 21138 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 5518 17838 5570 17890
rect 26014 17838 26066 17890
rect 2158 17726 2210 17778
rect 3950 17726 4002 17778
rect 21422 17726 21474 17778
rect 41806 17726 41858 17778
rect 43598 17726 43650 17778
rect 8542 17614 8594 17666
rect 9214 17614 9266 17666
rect 9438 17614 9490 17666
rect 9886 17614 9938 17666
rect 16494 17614 16546 17666
rect 17054 17614 17106 17666
rect 20190 17614 20242 17666
rect 20862 17614 20914 17666
rect 22318 17614 22370 17666
rect 22990 17614 23042 17666
rect 27358 17614 27410 17666
rect 32174 17614 32226 17666
rect 32510 17614 32562 17666
rect 35982 17614 36034 17666
rect 36542 17614 36594 17666
rect 36990 17614 37042 17666
rect 37550 17614 37602 17666
rect 1934 17502 1986 17554
rect 3054 17502 3106 17554
rect 14142 17502 14194 17554
rect 21646 17502 21698 17554
rect 25230 17502 25282 17554
rect 26574 17502 26626 17554
rect 26910 17502 26962 17554
rect 28142 17502 28194 17554
rect 39790 17502 39842 17554
rect 42814 17502 42866 17554
rect 43934 17502 43986 17554
rect 6302 17390 6354 17442
rect 12462 17390 12514 17442
rect 13022 17390 13074 17442
rect 13358 17390 13410 17442
rect 17166 17390 17218 17442
rect 17726 17390 17778 17442
rect 22094 17390 22146 17442
rect 29038 17390 29090 17442
rect 29598 17390 29650 17442
rect 32846 17390 32898 17442
rect 33630 17390 33682 17442
rect 40574 17390 40626 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 2158 17054 2210 17106
rect 6190 17054 6242 17106
rect 12574 17054 12626 17106
rect 16382 17054 16434 17106
rect 32622 17054 32674 17106
rect 36094 17054 36146 17106
rect 36654 17054 36706 17106
rect 39902 17054 39954 17106
rect 18846 16942 18898 16994
rect 22542 16942 22594 16994
rect 25902 16942 25954 16994
rect 31838 16942 31890 16994
rect 42926 16942 42978 16994
rect 43710 16942 43762 16994
rect 4734 16830 4786 16882
rect 5070 16830 5122 16882
rect 8430 16830 8482 16882
rect 8878 16830 8930 16882
rect 9438 16830 9490 16882
rect 10110 16830 10162 16882
rect 13246 16830 13298 16882
rect 13918 16830 13970 16882
rect 21198 16830 21250 16882
rect 21758 16830 21810 16882
rect 28254 16830 28306 16882
rect 28590 16830 28642 16882
rect 28926 16830 28978 16882
rect 29598 16830 29650 16882
rect 33182 16830 33234 16882
rect 33630 16830 33682 16882
rect 36990 16830 37042 16882
rect 37438 16830 37490 16882
rect 17502 16718 17554 16770
rect 17838 16718 17890 16770
rect 23438 16718 23490 16770
rect 41918 16718 41970 16770
rect 44046 16718 44098 16770
rect 1598 16606 1650 16658
rect 5406 16606 5458 16658
rect 13134 16606 13186 16658
rect 16942 16606 16994 16658
rect 18062 16606 18114 16658
rect 25118 16606 25170 16658
rect 40462 16606 40514 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 3838 16158 3890 16210
rect 15486 16158 15538 16210
rect 26910 16158 26962 16210
rect 27806 16158 27858 16210
rect 28590 16158 28642 16210
rect 41806 16158 41858 16210
rect 1934 16046 1986 16098
rect 10782 16046 10834 16098
rect 11342 16046 11394 16098
rect 11566 16046 11618 16098
rect 19742 16046 19794 16098
rect 20190 16046 20242 16098
rect 22766 16046 22818 16098
rect 23326 16046 23378 16098
rect 29038 16046 29090 16098
rect 29710 16046 29762 16098
rect 33070 16046 33122 16098
rect 33518 16046 33570 16098
rect 40014 16046 40066 16098
rect 40350 16046 40402 16098
rect 2718 15934 2770 15986
rect 5966 15934 6018 15986
rect 6302 15934 6354 15986
rect 14366 15934 14418 15986
rect 17502 15934 17554 15986
rect 21982 15934 22034 15986
rect 27470 15934 27522 15986
rect 28142 15934 28194 15986
rect 37662 15934 37714 15986
rect 42814 15934 42866 15986
rect 2046 15822 2098 15874
rect 7646 15822 7698 15874
rect 8430 15822 8482 15874
rect 12126 15822 12178 15874
rect 16718 15822 16770 15874
rect 22094 15822 22146 15874
rect 25790 15822 25842 15874
rect 26350 15822 26402 15874
rect 27358 15822 27410 15874
rect 32062 15822 32114 15874
rect 32734 15822 32786 15874
rect 35982 15822 36034 15874
rect 36542 15822 36594 15874
rect 36878 15822 36930 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 4958 15486 5010 15538
rect 24222 15486 24274 15538
rect 25342 15486 25394 15538
rect 30270 15486 30322 15538
rect 32510 15486 32562 15538
rect 38110 15486 38162 15538
rect 7982 15374 8034 15426
rect 9886 15374 9938 15426
rect 10222 15374 10274 15426
rect 11118 15374 11170 15426
rect 11454 15374 11506 15426
rect 12462 15374 12514 15426
rect 15598 15374 15650 15426
rect 17726 15374 17778 15426
rect 20750 15374 20802 15426
rect 25790 15374 25842 15426
rect 26126 15374 26178 15426
rect 26462 15374 26514 15426
rect 31054 15374 31106 15426
rect 31390 15374 31442 15426
rect 31726 15374 31778 15426
rect 32062 15374 32114 15426
rect 33070 15374 33122 15426
rect 34414 15374 34466 15426
rect 38894 15374 38946 15426
rect 42926 15374 42978 15426
rect 2270 15262 2322 15314
rect 2718 15262 2770 15314
rect 14814 15262 14866 15314
rect 15374 15262 15426 15314
rect 21310 15262 21362 15314
rect 21758 15262 21810 15314
rect 26686 15262 26738 15314
rect 27134 15262 27186 15314
rect 27806 15262 27858 15314
rect 33294 15262 33346 15314
rect 33742 15262 33794 15314
rect 34974 15262 35026 15314
rect 35646 15262 35698 15314
rect 39118 15262 39170 15314
rect 6974 15150 7026 15202
rect 15934 15150 15986 15202
rect 18062 15150 18114 15202
rect 19630 15150 19682 15202
rect 33966 15150 34018 15202
rect 34750 15150 34802 15202
rect 41918 15150 41970 15202
rect 5742 15038 5794 15090
rect 11678 15038 11730 15090
rect 24782 15038 24834 15090
rect 30830 15038 30882 15090
rect 38670 15038 38722 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 28142 14702 28194 14754
rect 28590 14702 28642 14754
rect 3502 14590 3554 14642
rect 7422 14590 7474 14642
rect 11454 14590 11506 14642
rect 14030 14590 14082 14642
rect 14366 14590 14418 14642
rect 14702 14590 14754 14642
rect 15038 14590 15090 14642
rect 16830 14590 16882 14642
rect 19742 14590 19794 14642
rect 21422 14590 21474 14642
rect 27246 14590 27298 14642
rect 27582 14590 27634 14642
rect 27694 14590 27746 14642
rect 28142 14590 28194 14642
rect 28590 14590 28642 14642
rect 34302 14590 34354 14642
rect 36094 14590 36146 14642
rect 41806 14590 41858 14642
rect 23438 14478 23490 14530
rect 23886 14478 23938 14530
rect 32510 14478 32562 14530
rect 33070 14478 33122 14530
rect 36318 14478 36370 14530
rect 40014 14478 40066 14530
rect 40350 14478 40402 14530
rect 2382 14366 2434 14418
rect 6078 14366 6130 14418
rect 12462 14366 12514 14418
rect 15934 14366 15986 14418
rect 18510 14366 18562 14418
rect 21646 14366 21698 14418
rect 30158 14366 30210 14418
rect 35310 14366 35362 14418
rect 37662 14366 37714 14418
rect 42926 14366 42978 14418
rect 26350 14254 26402 14306
rect 26910 14254 26962 14306
rect 29374 14254 29426 14306
rect 36878 14254 36930 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 5406 13918 5458 13970
rect 8430 13806 8482 13858
rect 12798 13806 12850 13858
rect 15262 13806 15314 13858
rect 20974 13806 21026 13858
rect 21646 13806 21698 13858
rect 29262 13806 29314 13858
rect 31950 13806 32002 13858
rect 35758 13806 35810 13858
rect 38222 13806 38274 13858
rect 2270 13694 2322 13746
rect 2942 13694 2994 13746
rect 7198 13582 7250 13634
rect 11454 13582 11506 13634
rect 14254 13582 14306 13634
rect 19742 13582 19794 13634
rect 22990 13582 23042 13634
rect 28366 13582 28418 13634
rect 30942 13582 30994 13634
rect 34414 13582 34466 13634
rect 37214 13582 37266 13634
rect 5966 13470 6018 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 3614 13022 3666 13074
rect 11566 13022 11618 13074
rect 15262 13022 15314 13074
rect 19070 13022 19122 13074
rect 26686 13022 26738 13074
rect 30158 13022 30210 13074
rect 34302 13022 34354 13074
rect 37998 13022 38050 13074
rect 40798 13022 40850 13074
rect 25678 12910 25730 12962
rect 26238 12910 26290 12962
rect 4958 12798 5010 12850
rect 12462 12798 12514 12850
rect 16606 12798 16658 12850
rect 17838 12798 17890 12850
rect 23326 12798 23378 12850
rect 31166 12798 31218 12850
rect 35646 12798 35698 12850
rect 39006 12798 39058 12850
rect 42030 12798 42082 12850
rect 22542 12686 22594 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 14254 12238 14306 12290
rect 17502 12238 17554 12290
rect 23550 12238 23602 12290
rect 27246 12238 27298 12290
rect 30382 12238 30434 12290
rect 35422 12238 35474 12290
rect 15374 12014 15426 12066
rect 18734 12014 18786 12066
rect 22318 12014 22370 12066
rect 26238 12014 26290 12066
rect 29038 12014 29090 12066
rect 34078 12014 34130 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 24110 11454 24162 11506
rect 26686 11454 26738 11506
rect 33518 11454 33570 11506
rect 22990 11230 23042 11282
rect 28030 11230 28082 11282
rect 34862 11230 34914 11282
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 20078 9102 20130 9154
rect 20862 9102 20914 9154
rect 43822 9102 43874 9154
rect 19742 8990 19794 9042
rect 20638 8990 20690 9042
rect 44158 8990 44210 9042
rect 43598 8878 43650 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 27022 8206 27074 8258
rect 42926 8206 42978 8258
rect 44046 8094 44098 8146
rect 27246 7982 27298 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 42590 7534 42642 7586
rect 42926 7422 42978 7474
rect 44046 7422 44098 7474
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 43150 6638 43202 6690
rect 24446 6526 24498 6578
rect 44046 6526 44098 6578
rect 24782 6414 24834 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 42926 5854 42978 5906
rect 42254 5742 42306 5794
rect 42702 5742 42754 5794
rect 44046 5742 44098 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 25118 5070 25170 5122
rect 33406 5070 33458 5122
rect 37438 5070 37490 5122
rect 38110 5070 38162 5122
rect 38670 5070 38722 5122
rect 43822 5070 43874 5122
rect 31838 4958 31890 5010
rect 37886 4958 37938 5010
rect 39230 4958 39282 5010
rect 41470 4958 41522 5010
rect 41806 4958 41858 5010
rect 42142 4958 42194 5010
rect 42478 4958 42530 5010
rect 42814 4958 42866 5010
rect 43150 4958 43202 5010
rect 43486 4958 43538 5010
rect 25342 4846 25394 4898
rect 32174 4846 32226 4898
rect 33630 4846 33682 4898
rect 35870 4846 35922 4898
rect 36542 4846 36594 4898
rect 37214 4846 37266 4898
rect 38894 4846 38946 4898
rect 39566 4846 39618 4898
rect 40686 4846 40738 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 20078 4510 20130 4562
rect 20750 4510 20802 4562
rect 25230 4510 25282 4562
rect 27134 4510 27186 4562
rect 33518 4510 33570 4562
rect 35758 4510 35810 4562
rect 36430 4510 36482 4562
rect 37102 4510 37154 4562
rect 38894 4510 38946 4562
rect 40910 4510 40962 4562
rect 42814 4510 42866 4562
rect 43822 4510 43874 4562
rect 19070 4398 19122 4450
rect 26462 4398 26514 4450
rect 32398 4398 32450 4450
rect 38222 4398 38274 4450
rect 39902 4398 39954 4450
rect 41582 4398 41634 4450
rect 42366 4398 42418 4450
rect 43150 4398 43202 4450
rect 19742 4286 19794 4338
rect 20414 4286 20466 4338
rect 25566 4286 25618 4338
rect 27358 4286 27410 4338
rect 33182 4286 33234 4338
rect 36094 4286 36146 4338
rect 36766 4286 36818 4338
rect 37998 4286 38050 4338
rect 38558 4286 38610 4338
rect 41134 4286 41186 4338
rect 41806 4286 41858 4338
rect 43374 4286 43426 4338
rect 44046 4286 44098 4338
rect 19518 4174 19570 4226
rect 24222 4174 24274 4226
rect 24782 4174 24834 4226
rect 26238 4174 26290 4226
rect 32174 4174 32226 4226
rect 37662 4174 37714 4226
rect 34974 4062 35026 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 21534 3614 21586 3666
rect 26574 3614 26626 3666
rect 28814 3614 28866 3666
rect 32622 3614 32674 3666
rect 34302 3614 34354 3666
rect 40238 3614 40290 3666
rect 42254 3614 42306 3666
rect 20078 3502 20130 3554
rect 21086 3502 21138 3554
rect 23774 3502 23826 3554
rect 25230 3502 25282 3554
rect 26126 3502 26178 3554
rect 28366 3502 28418 3554
rect 32174 3502 32226 3554
rect 33854 3502 33906 3554
rect 37214 3502 37266 3554
rect 39118 3502 39170 3554
rect 39790 3502 39842 3554
rect 23998 3390 24050 3442
rect 30942 3390 30994 3442
rect 31166 3390 31218 3442
rect 31502 3390 31554 3442
rect 41246 3390 41298 3442
rect 41806 3390 41858 3442
rect 43150 3390 43202 3442
rect 43822 3390 43874 3442
rect 44158 3390 44210 3442
rect 19406 3278 19458 3330
rect 22654 3278 22706 3330
rect 24558 3278 24610 3330
rect 36430 3278 36482 3330
rect 37550 3278 37602 3330
rect 38446 3278 38498 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 14112 45200 14224 46000
rect 14784 45200 14896 46000
rect 15456 45200 15568 46000
rect 16128 45200 16240 46000
rect 16800 45200 16912 46000
rect 17472 45200 17584 46000
rect 18144 45200 18256 46000
rect 18816 45200 18928 46000
rect 19488 45200 19600 46000
rect 20160 45200 20272 46000
rect 20832 45200 20944 46000
rect 21504 45200 21616 46000
rect 22176 45200 22288 46000
rect 22540 45276 22932 45332
rect 14140 43708 14196 45200
rect 14812 43708 14868 45200
rect 13916 43652 14196 43708
rect 14588 43652 14868 43708
rect 15484 43708 15540 45200
rect 16156 43708 16212 45200
rect 16828 43708 16884 45200
rect 17500 43708 17556 45200
rect 15484 43652 15652 43708
rect 16156 43652 16436 43708
rect 16828 43652 17108 43708
rect 17500 43652 17780 43708
rect 13916 41972 13972 43652
rect 14140 42082 14196 42094
rect 14140 42030 14142 42082
rect 14194 42030 14196 42082
rect 14140 41972 14196 42030
rect 14588 41972 14644 43652
rect 15596 42194 15652 43652
rect 15596 42142 15598 42194
rect 15650 42142 15652 42194
rect 15596 42130 15652 42142
rect 13916 41970 14084 41972
rect 13916 41918 13918 41970
rect 13970 41918 14084 41970
rect 13916 41916 14084 41918
rect 14140 41916 14532 41972
rect 13916 41906 13972 41916
rect 14028 41860 14084 41916
rect 14028 41804 14420 41860
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 14364 41298 14420 41804
rect 14364 41246 14366 41298
rect 14418 41246 14420 41298
rect 14364 41234 14420 41246
rect 14476 40516 14532 41916
rect 14588 41878 14644 41916
rect 14812 42082 14868 42094
rect 14812 42030 14814 42082
rect 14866 42030 14868 42082
rect 14476 40450 14532 40460
rect 14812 40514 14868 42030
rect 15260 41972 15316 41982
rect 16268 41972 16324 41982
rect 15260 41878 15316 41916
rect 15820 41970 16324 41972
rect 15820 41918 16270 41970
rect 16322 41918 16324 41970
rect 15820 41916 16324 41918
rect 15148 41188 15204 41198
rect 15148 40626 15204 41132
rect 15148 40574 15150 40626
rect 15202 40574 15204 40626
rect 15148 40562 15204 40574
rect 15820 40626 15876 41916
rect 16268 41906 16324 41916
rect 16380 41972 16436 43652
rect 16380 41906 16436 41916
rect 16940 41970 16996 41982
rect 16940 41918 16942 41970
rect 16994 41918 16996 41970
rect 16940 41188 16996 41918
rect 16940 41122 16996 41132
rect 17052 41074 17108 43652
rect 17388 41972 17444 41982
rect 17388 41858 17444 41916
rect 17388 41806 17390 41858
rect 17442 41806 17444 41858
rect 17388 41794 17444 41806
rect 17724 41188 17780 43652
rect 18172 41412 18228 45200
rect 18172 41346 18228 41356
rect 17052 41022 17054 41074
rect 17106 41022 17108 41074
rect 17052 41010 17108 41022
rect 17164 41186 17780 41188
rect 17164 41134 17726 41186
rect 17778 41134 17780 41186
rect 17164 41132 17780 41134
rect 16828 40962 16884 40974
rect 16828 40910 16830 40962
rect 16882 40910 16884 40962
rect 16828 40852 16884 40910
rect 17164 40852 17220 41132
rect 17724 41122 17780 41132
rect 18844 41188 18900 45200
rect 19516 43708 19572 45200
rect 19404 43652 19572 43708
rect 19404 42194 19460 43652
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19404 42142 19406 42194
rect 19458 42142 19460 42194
rect 19404 42130 19460 42142
rect 20076 41972 20132 41982
rect 19516 41970 20132 41972
rect 19516 41918 20078 41970
rect 20130 41918 20132 41970
rect 19516 41916 20132 41918
rect 19292 41412 19348 41422
rect 19292 41298 19348 41356
rect 19292 41246 19294 41298
rect 19346 41246 19348 41298
rect 19292 41234 19348 41246
rect 18844 41122 18900 41132
rect 18060 40964 18116 40974
rect 18060 40962 18564 40964
rect 18060 40910 18062 40962
rect 18114 40910 18564 40962
rect 18060 40908 18564 40910
rect 18060 40898 18116 40908
rect 16828 40796 17220 40852
rect 15820 40574 15822 40626
rect 15874 40574 15876 40626
rect 15820 40562 15876 40574
rect 14812 40462 14814 40514
rect 14866 40462 14868 40514
rect 14812 40450 14868 40462
rect 15484 40516 15540 40526
rect 15484 40422 15540 40460
rect 18508 40514 18564 40908
rect 18844 40962 18900 40974
rect 18844 40910 18846 40962
rect 18898 40910 18900 40962
rect 18844 40626 18900 40910
rect 18844 40574 18846 40626
rect 18898 40574 18900 40626
rect 18844 40562 18900 40574
rect 19516 40628 19572 41916
rect 20076 41906 20132 41916
rect 20188 41300 20244 45200
rect 20860 43708 20916 45200
rect 20860 43652 21364 43708
rect 20860 41970 20916 41982
rect 20860 41918 20862 41970
rect 20914 41918 20916 41970
rect 20188 41298 20468 41300
rect 20188 41246 20190 41298
rect 20242 41246 20468 41298
rect 20188 41244 20468 41246
rect 20188 41234 20244 41244
rect 20412 41186 20468 41244
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 20412 41122 20468 41134
rect 20188 41076 20244 41086
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19740 40628 19796 40638
rect 19516 40626 19796 40628
rect 19516 40574 19742 40626
rect 19794 40574 19796 40626
rect 19516 40572 19796 40574
rect 19740 40562 19796 40572
rect 18508 40462 18510 40514
rect 18562 40462 18564 40514
rect 18508 40450 18564 40462
rect 20076 40514 20132 40526
rect 20076 40462 20078 40514
rect 20130 40462 20132 40514
rect 19516 40404 19572 40414
rect 20076 40404 20132 40462
rect 19516 40402 20132 40404
rect 19516 40350 19518 40402
rect 19570 40350 20132 40402
rect 19516 40348 20132 40350
rect 20188 40404 20244 41020
rect 20748 40964 20804 40974
rect 20524 40962 20804 40964
rect 20524 40910 20750 40962
rect 20802 40910 20804 40962
rect 20524 40908 20804 40910
rect 20300 40404 20356 40414
rect 20188 40402 20356 40404
rect 20188 40350 20302 40402
rect 20354 40350 20356 40402
rect 20188 40348 20356 40350
rect 19516 40338 19572 40348
rect 20188 40292 20244 40348
rect 20300 40338 20356 40348
rect 19852 40236 20244 40292
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 19852 39730 19908 40236
rect 19852 39678 19854 39730
rect 19906 39678 19908 39730
rect 19852 39666 19908 39678
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20524 35698 20580 40908
rect 20748 40898 20804 40908
rect 20748 35924 20804 35934
rect 20860 35924 20916 41918
rect 21308 41858 21364 43652
rect 21308 41806 21310 41858
rect 21362 41806 21364 41858
rect 21308 41794 21364 41806
rect 21532 41300 21588 45200
rect 22204 45108 22260 45200
rect 22540 45108 22596 45276
rect 22204 45052 22596 45108
rect 22428 41970 22484 41982
rect 22428 41918 22430 41970
rect 22482 41918 22484 41970
rect 21532 41298 22036 41300
rect 21532 41246 21534 41298
rect 21586 41246 22036 41298
rect 21532 41244 22036 41246
rect 21532 41234 21588 41244
rect 21980 41186 22036 41244
rect 21980 41134 21982 41186
rect 22034 41134 22036 41186
rect 21980 41122 22036 41134
rect 21756 40964 21812 40974
rect 21644 40962 21812 40964
rect 21644 40910 21758 40962
rect 21810 40910 21812 40962
rect 21644 40908 21812 40910
rect 21644 38276 21700 40908
rect 21756 40898 21812 40908
rect 20748 35922 20916 35924
rect 20748 35870 20750 35922
rect 20802 35870 20916 35922
rect 20748 35868 20916 35870
rect 21420 38220 21700 38276
rect 20748 35858 20804 35868
rect 20524 35646 20526 35698
rect 20578 35646 20580 35698
rect 20524 35634 20580 35646
rect 21420 35698 21476 38220
rect 21644 35924 21700 35934
rect 21644 35830 21700 35868
rect 22428 35924 22484 41918
rect 22876 41858 22932 45276
rect 23520 45200 23632 46000
rect 24192 45200 24304 46000
rect 24864 45200 24976 46000
rect 25536 45200 25648 46000
rect 26208 45200 26320 46000
rect 26880 45200 26992 46000
rect 27552 45200 27664 46000
rect 30912 45200 31024 46000
rect 31584 45200 31696 46000
rect 32256 45200 32368 46000
rect 32928 45200 33040 46000
rect 34272 45200 34384 46000
rect 35616 45200 35728 46000
rect 36288 45200 36400 46000
rect 36960 45200 37072 46000
rect 37632 45200 37744 46000
rect 38304 45200 38416 46000
rect 38976 45200 39088 46000
rect 39648 45200 39760 46000
rect 40320 45200 40432 46000
rect 40992 45200 41104 46000
rect 41664 45200 41776 46000
rect 41916 45780 41972 45790
rect 22876 41806 22878 41858
rect 22930 41806 22932 41858
rect 22876 41794 22932 41806
rect 23548 41300 23604 45200
rect 24220 43708 24276 45200
rect 24892 43708 24948 45200
rect 25564 43708 25620 45200
rect 24220 43652 24836 43708
rect 24892 43652 25172 43708
rect 25564 43652 26068 43708
rect 24780 42756 24836 43652
rect 24780 42700 25060 42756
rect 24556 41970 24612 41982
rect 24556 41918 24558 41970
rect 24610 41918 24612 41970
rect 23548 41298 23828 41300
rect 23548 41246 23550 41298
rect 23602 41246 23828 41298
rect 23548 41244 23828 41246
rect 23548 41234 23604 41244
rect 23772 41186 23828 41244
rect 23772 41134 23774 41186
rect 23826 41134 23828 41186
rect 23772 41122 23828 41134
rect 22428 35858 22484 35868
rect 24108 40962 24164 40974
rect 24108 40910 24110 40962
rect 24162 40910 24164 40962
rect 24108 35810 24164 40910
rect 24444 35924 24500 35934
rect 24556 35924 24612 41918
rect 25004 41858 25060 42700
rect 25004 41806 25006 41858
rect 25058 41806 25060 41858
rect 25004 41794 25060 41806
rect 24892 41300 24948 41310
rect 24892 41206 24948 41244
rect 25116 41074 25172 43652
rect 26012 41300 26068 43652
rect 26236 41972 26292 45200
rect 26908 43708 26964 45200
rect 27580 43708 27636 45200
rect 30940 43708 30996 45200
rect 31612 43708 31668 45200
rect 32284 43708 32340 45200
rect 32956 43708 33012 45200
rect 34300 43708 34356 45200
rect 26908 43652 27524 43708
rect 27580 43652 27972 43708
rect 30940 43652 31220 43708
rect 31612 43652 31892 43708
rect 32284 43652 32564 43708
rect 32956 43652 33236 43708
rect 34300 43652 34804 43708
rect 26460 41972 26516 41982
rect 26236 41906 26292 41916
rect 26348 41970 26516 41972
rect 26348 41918 26462 41970
rect 26514 41918 26516 41970
rect 26348 41916 26516 41918
rect 26012 41186 26068 41244
rect 26012 41134 26014 41186
rect 26066 41134 26068 41186
rect 26012 41122 26068 41134
rect 25116 41022 25118 41074
rect 25170 41022 25172 41074
rect 25116 41010 25172 41022
rect 25788 40964 25844 40974
rect 24444 35922 24612 35924
rect 24444 35870 24446 35922
rect 24498 35870 24612 35922
rect 24444 35868 24612 35870
rect 25564 40962 25844 40964
rect 25564 40910 25790 40962
rect 25842 40910 25844 40962
rect 25564 40908 25844 40910
rect 24444 35858 24500 35868
rect 24108 35758 24110 35810
rect 24162 35758 24164 35810
rect 24108 35746 24164 35758
rect 21420 35646 21422 35698
rect 21474 35646 21476 35698
rect 21420 35634 21476 35646
rect 25564 35698 25620 40908
rect 25788 40898 25844 40908
rect 26348 38948 26404 41916
rect 26460 41906 26516 41916
rect 26908 41972 26964 41982
rect 26908 41858 26964 41916
rect 26908 41806 26910 41858
rect 26962 41806 26964 41858
rect 26908 41794 26964 41806
rect 27468 41300 27524 43652
rect 27916 41972 27972 43652
rect 31164 42194 31220 43652
rect 31164 42142 31166 42194
rect 31218 42142 31220 42194
rect 31164 42130 31220 42142
rect 27916 41878 27972 41916
rect 28364 42082 28420 42094
rect 28364 42030 28366 42082
rect 28418 42030 28420 42082
rect 27580 41300 27636 41310
rect 27468 41298 27636 41300
rect 27468 41246 27582 41298
rect 27634 41246 27636 41298
rect 27468 41244 27636 41246
rect 27580 41234 27636 41244
rect 25788 38892 26404 38948
rect 27132 40962 27188 40974
rect 27132 40910 27134 40962
rect 27186 40910 27188 40962
rect 25788 35922 25844 38892
rect 25788 35870 25790 35922
rect 25842 35870 25844 35922
rect 25788 35858 25844 35870
rect 26236 38612 26292 38622
rect 25564 35646 25566 35698
rect 25618 35646 25620 35698
rect 25564 35634 25620 35646
rect 26236 35698 26292 38556
rect 26460 35924 26516 35934
rect 26460 35830 26516 35868
rect 27132 35924 27188 40910
rect 28364 38612 28420 42030
rect 28588 41972 28644 41982
rect 28588 41878 28644 41916
rect 31836 41074 31892 43652
rect 32508 41970 32564 43652
rect 33180 42194 33236 43652
rect 33180 42142 33182 42194
rect 33234 42142 33236 42194
rect 33180 42130 33236 42142
rect 34748 42194 34804 43652
rect 34748 42142 34750 42194
rect 34802 42142 34804 42194
rect 34748 42130 34804 42142
rect 32508 41918 32510 41970
rect 32562 41918 32564 41970
rect 32508 41298 32564 41918
rect 32508 41246 32510 41298
rect 32562 41246 32564 41298
rect 32508 41234 32564 41246
rect 32844 42082 32900 42094
rect 32844 42030 32846 42082
rect 32898 42030 32900 42082
rect 31836 41022 31838 41074
rect 31890 41022 31892 41074
rect 31836 41010 31892 41022
rect 32844 40516 32900 42030
rect 33852 41972 33908 41982
rect 33404 41970 33908 41972
rect 33404 41918 33854 41970
rect 33906 41918 33908 41970
rect 33404 41916 33908 41918
rect 33404 40626 33460 41916
rect 33852 41906 33908 41916
rect 35532 41972 35588 41982
rect 35644 41972 35700 45200
rect 36316 43708 36372 45200
rect 36988 43708 37044 45200
rect 36316 43652 36708 43708
rect 36988 43652 37268 43708
rect 36652 42194 36708 43652
rect 36652 42142 36654 42194
rect 36706 42142 36708 42194
rect 36652 42130 36708 42142
rect 36316 42082 36372 42094
rect 36316 42030 36318 42082
rect 36370 42030 36372 42082
rect 35980 41972 36036 41982
rect 35532 41970 36036 41972
rect 35532 41918 35534 41970
rect 35586 41918 35982 41970
rect 36034 41918 36036 41970
rect 35532 41916 36036 41918
rect 35532 41906 35588 41916
rect 35980 41906 36036 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 33404 40574 33406 40626
rect 33458 40574 33460 40626
rect 33404 40562 33460 40574
rect 33068 40516 33124 40526
rect 32844 40514 33124 40516
rect 32844 40462 33070 40514
rect 33122 40462 33124 40514
rect 32844 40460 33124 40462
rect 33068 40450 33124 40460
rect 36316 40516 36372 42030
rect 37212 41970 37268 43652
rect 37212 41918 37214 41970
rect 37266 41918 37268 41970
rect 37212 41298 37268 41918
rect 37212 41246 37214 41298
rect 37266 41246 37268 41298
rect 37212 41234 37268 41246
rect 37548 42082 37604 42094
rect 37548 42030 37550 42082
rect 37602 42030 37604 42082
rect 36316 40450 36372 40460
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 37548 39620 37604 42030
rect 37660 41300 37716 45200
rect 38332 43708 38388 45200
rect 38332 43652 38500 43708
rect 38444 42194 38500 43652
rect 38444 42142 38446 42194
rect 38498 42142 38500 42194
rect 38444 42130 38500 42142
rect 39004 41972 39060 45200
rect 39676 43708 39732 45200
rect 40348 43708 40404 45200
rect 41020 43708 41076 45200
rect 41692 43708 41748 45200
rect 39676 43652 40292 43708
rect 40348 43652 40964 43708
rect 41020 43652 41412 43708
rect 39004 41906 39060 41916
rect 39228 41972 39284 41982
rect 39788 41972 39844 41982
rect 39228 41970 39508 41972
rect 39228 41918 39230 41970
rect 39282 41918 39508 41970
rect 39228 41916 39508 41918
rect 39228 41906 39284 41916
rect 37660 41298 37940 41300
rect 37660 41246 37662 41298
rect 37714 41246 37940 41298
rect 37660 41244 37940 41246
rect 37660 41234 37716 41244
rect 37884 41186 37940 41244
rect 37884 41134 37886 41186
rect 37938 41134 37940 41186
rect 37884 41122 37940 41134
rect 38220 40964 38276 40974
rect 38220 40870 38276 40908
rect 39452 40626 39508 41916
rect 39676 41970 39844 41972
rect 39676 41918 39790 41970
rect 39842 41918 39844 41970
rect 39676 41916 39844 41918
rect 39452 40574 39454 40626
rect 39506 40574 39508 40626
rect 39452 40562 39508 40574
rect 39564 40962 39620 40974
rect 39564 40910 39566 40962
rect 39618 40910 39620 40962
rect 39564 40628 39620 40910
rect 39564 40562 39620 40572
rect 38780 40516 38836 40526
rect 38780 40422 38836 40460
rect 39116 40514 39172 40526
rect 39116 40462 39118 40514
rect 39170 40462 39172 40514
rect 39116 40404 39172 40462
rect 39676 40404 39732 41916
rect 39788 41906 39844 41916
rect 40236 41300 40292 43652
rect 40348 41972 40404 41982
rect 40348 41858 40404 41916
rect 40348 41806 40350 41858
rect 40402 41806 40404 41858
rect 40348 41794 40404 41806
rect 40348 41300 40404 41310
rect 40236 41298 40404 41300
rect 40236 41246 40350 41298
rect 40402 41246 40404 41298
rect 40236 41244 40404 41246
rect 40348 41234 40404 41244
rect 40908 41188 40964 43652
rect 41356 42194 41412 43652
rect 41356 42142 41358 42194
rect 41410 42142 41412 42194
rect 41356 42130 41412 42142
rect 41468 43652 41748 43708
rect 40684 41132 41188 41188
rect 39788 40964 39844 40974
rect 39788 40514 39844 40908
rect 39788 40462 39790 40514
rect 39842 40462 39844 40514
rect 39788 40450 39844 40462
rect 39900 40962 39956 40974
rect 39900 40910 39902 40962
rect 39954 40910 39956 40962
rect 39116 40348 39732 40404
rect 39900 40180 39956 40910
rect 39452 40124 39956 40180
rect 40124 40852 40180 40862
rect 37548 39554 37604 39564
rect 39116 39620 39172 39630
rect 39116 39526 39172 39564
rect 39452 39506 39508 40124
rect 39900 39620 39956 39630
rect 39900 39526 39956 39564
rect 39452 39454 39454 39506
rect 39506 39454 39508 39506
rect 39452 39442 39508 39454
rect 40124 39506 40180 40796
rect 40348 40514 40404 40526
rect 40348 40462 40350 40514
rect 40402 40462 40404 40514
rect 40348 39732 40404 40462
rect 40348 39666 40404 39676
rect 40684 39730 40740 41132
rect 40684 39678 40686 39730
rect 40738 39678 40740 39730
rect 40684 39666 40740 39678
rect 40908 40514 40964 40526
rect 40908 40462 40910 40514
rect 40962 40462 40964 40514
rect 40908 39620 40964 40462
rect 41132 40402 41188 41132
rect 41132 40350 41134 40402
rect 41186 40350 41188 40402
rect 41132 40338 41188 40350
rect 40908 39554 40964 39564
rect 40124 39454 40126 39506
rect 40178 39454 40180 39506
rect 40124 39442 40180 39454
rect 41468 39506 41524 43652
rect 41804 41970 41860 41982
rect 41804 41918 41806 41970
rect 41858 41918 41860 41970
rect 41692 40964 41748 40974
rect 41692 40628 41748 40908
rect 41804 40852 41860 41918
rect 41916 41300 41972 45724
rect 42336 45200 42448 46000
rect 42364 41858 42420 45200
rect 44268 45108 44324 45118
rect 43932 44436 43988 44446
rect 43708 43764 43764 43774
rect 43484 42420 43540 42430
rect 43372 42364 43484 42420
rect 42364 41806 42366 41858
rect 42418 41806 42420 41858
rect 42364 41794 42420 41806
rect 43148 41860 43204 41870
rect 43148 41766 43204 41804
rect 42028 41300 42084 41310
rect 41916 41298 42084 41300
rect 41916 41246 42030 41298
rect 42082 41246 42084 41298
rect 41916 41244 42084 41246
rect 42028 41234 42084 41244
rect 41804 40786 41860 40796
rect 42476 41186 42532 41198
rect 42924 41188 42980 41198
rect 42476 41134 42478 41186
rect 42530 41134 42532 41186
rect 41692 40572 41860 40628
rect 41692 40404 41748 40414
rect 41692 40310 41748 40348
rect 41804 39618 41860 40572
rect 41916 40516 41972 40526
rect 41916 40422 41972 40460
rect 41804 39566 41806 39618
rect 41858 39566 41860 39618
rect 41804 39554 41860 39566
rect 42364 40402 42420 40414
rect 42364 40350 42366 40402
rect 42418 40350 42420 40402
rect 41468 39454 41470 39506
rect 41522 39454 41524 39506
rect 41468 39442 41524 39454
rect 42140 39506 42196 39518
rect 42140 39454 42142 39506
rect 42194 39454 42196 39506
rect 42140 39396 42196 39454
rect 42252 39396 42308 39406
rect 42140 39340 42252 39396
rect 42252 39330 42308 39340
rect 42364 39284 42420 40350
rect 42476 39506 42532 41134
rect 42588 41186 42980 41188
rect 42588 41134 42926 41186
rect 42978 41134 42980 41186
rect 42588 41132 42980 41134
rect 42588 40626 42644 41132
rect 42924 41122 42980 41132
rect 42588 40574 42590 40626
rect 42642 40574 42644 40626
rect 42588 40562 42644 40574
rect 42924 40516 42980 40526
rect 42924 40422 42980 40460
rect 43372 39844 43428 42364
rect 43484 42354 43540 42364
rect 43708 40626 43764 43708
rect 43708 40574 43710 40626
rect 43762 40574 43764 40626
rect 43708 40562 43764 40574
rect 43820 42082 43876 42094
rect 43820 42030 43822 42082
rect 43874 42030 43876 42082
rect 43820 40628 43876 42030
rect 43932 40628 43988 44380
rect 44156 41970 44212 41982
rect 44156 41918 44158 41970
rect 44210 41918 44212 41970
rect 44156 41860 44212 41918
rect 44156 41794 44212 41804
rect 44044 41748 44100 41758
rect 44044 41298 44100 41692
rect 44044 41246 44046 41298
rect 44098 41246 44100 41298
rect 44044 41234 44100 41246
rect 44156 40628 44212 40638
rect 43932 40626 44212 40628
rect 43932 40574 44158 40626
rect 44210 40574 44212 40626
rect 43932 40572 44212 40574
rect 43820 40562 43876 40572
rect 43484 40404 43540 40414
rect 43540 40348 43764 40404
rect 43484 40338 43540 40348
rect 43372 39788 43540 39844
rect 42476 39454 42478 39506
rect 42530 39454 42532 39506
rect 42476 39442 42532 39454
rect 42812 39508 42868 39518
rect 42812 39414 42868 39452
rect 43372 39396 43428 39406
rect 43372 39302 43428 39340
rect 42364 39228 43204 39284
rect 42364 39060 42420 39070
rect 42364 38966 42420 39004
rect 43148 39058 43204 39228
rect 43148 39006 43150 39058
rect 43202 39006 43204 39058
rect 43148 38994 43204 39006
rect 28364 38546 28420 38556
rect 42812 38946 42868 38958
rect 42812 38894 42814 38946
rect 42866 38894 42868 38946
rect 42812 38612 42868 38894
rect 43484 38948 43540 39788
rect 43484 38946 43652 38948
rect 43484 38894 43486 38946
rect 43538 38894 43652 38946
rect 43484 38892 43652 38894
rect 43484 38882 43540 38892
rect 42812 38546 42868 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 43148 38164 43204 38174
rect 43148 38070 43204 38108
rect 43484 37828 43540 37838
rect 43484 37734 43540 37772
rect 43596 37716 43652 38892
rect 43708 37940 43764 40348
rect 43820 39508 43876 39518
rect 43820 39058 43876 39452
rect 43820 39006 43822 39058
rect 43874 39006 43876 39058
rect 43820 38994 43876 39006
rect 44044 38834 44100 40572
rect 44156 40562 44212 40572
rect 44156 39844 44212 39854
rect 44268 39844 44324 45052
rect 44156 39842 44324 39844
rect 44156 39790 44158 39842
rect 44210 39790 44324 39842
rect 44156 39788 44324 39790
rect 44380 43092 44436 43102
rect 44156 39778 44212 39788
rect 44044 38782 44046 38834
rect 44098 38782 44100 38834
rect 44044 38770 44100 38782
rect 44044 38164 44100 38174
rect 44044 38050 44100 38108
rect 44380 38164 44436 43036
rect 44492 41860 44548 41870
rect 44492 41076 44548 41804
rect 44492 41010 44548 41020
rect 44380 38098 44436 38108
rect 44044 37998 44046 38050
rect 44098 37998 44100 38050
rect 44044 37986 44100 37998
rect 43820 37940 43876 37950
rect 43708 37938 43876 37940
rect 43708 37886 43822 37938
rect 43874 37886 43876 37938
rect 43708 37884 43876 37886
rect 43820 37874 43876 37884
rect 43596 37660 43764 37716
rect 43708 37492 43764 37660
rect 43820 37492 43876 37502
rect 43708 37490 43876 37492
rect 43708 37438 43822 37490
rect 43874 37438 43876 37490
rect 43708 37436 43876 37438
rect 43820 37426 43876 37436
rect 44156 37378 44212 37390
rect 44156 37326 44158 37378
rect 44210 37326 44212 37378
rect 44156 37044 44212 37326
rect 44156 36978 44212 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 43708 36372 43764 36382
rect 43708 36278 43764 36316
rect 44156 36260 44212 36270
rect 44156 36258 44324 36260
rect 44156 36206 44158 36258
rect 44210 36206 44324 36258
rect 44156 36204 44324 36206
rect 44156 36194 44212 36204
rect 27132 35858 27188 35868
rect 44156 35812 44212 35822
rect 44156 35718 44212 35756
rect 26236 35646 26238 35698
rect 26290 35646 26292 35698
rect 26236 35634 26292 35646
rect 44268 35700 44324 36204
rect 44268 35634 44324 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 11452 31890 11508 31902
rect 18508 31892 18564 31902
rect 11452 31838 11454 31890
rect 11506 31838 11508 31890
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 6636 30324 6692 30334
rect 5180 30322 6692 30324
rect 5180 30270 6638 30322
rect 6690 30270 6692 30322
rect 5180 30268 6692 30270
rect 4508 29540 4564 29550
rect 4284 29538 4564 29540
rect 4284 29486 4510 29538
rect 4562 29486 4564 29538
rect 4284 29484 4564 29486
rect 1820 29426 1876 29438
rect 2156 29428 2212 29438
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 28644 1876 29374
rect 1820 28578 1876 28588
rect 2044 29426 2212 29428
rect 2044 29374 2158 29426
rect 2210 29374 2212 29426
rect 2044 29372 2212 29374
rect 2044 28082 2100 29372
rect 2156 29362 2212 29372
rect 3612 28980 3668 28990
rect 2044 28030 2046 28082
rect 2098 28030 2100 28082
rect 2044 28018 2100 28030
rect 3052 28756 3108 28766
rect 3052 28082 3108 28700
rect 3052 28030 3054 28082
rect 3106 28030 3108 28082
rect 3052 28018 3108 28030
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27636 1764 27806
rect 3052 27748 3108 27758
rect 1708 27188 1764 27580
rect 2268 27636 2324 27646
rect 2268 27634 2772 27636
rect 2268 27582 2270 27634
rect 2322 27582 2772 27634
rect 2268 27580 2772 27582
rect 2268 27570 2324 27580
rect 1820 27188 1876 27198
rect 1708 27186 1876 27188
rect 1708 27134 1822 27186
rect 1874 27134 1876 27186
rect 1708 27132 1876 27134
rect 1820 27122 1876 27132
rect 2716 26962 2772 27580
rect 2716 26910 2718 26962
rect 2770 26910 2772 26962
rect 2716 26898 2772 26910
rect 3052 26402 3108 27692
rect 3052 26350 3054 26402
rect 3106 26350 3108 26402
rect 3052 26338 3108 26350
rect 2492 26292 2548 26302
rect 2828 26292 2884 26302
rect 2492 26290 2884 26292
rect 2492 26238 2494 26290
rect 2546 26238 2830 26290
rect 2882 26238 2884 26290
rect 2492 26236 2884 26238
rect 2492 26226 2548 26236
rect 2828 26180 2884 26236
rect 3388 26180 3444 26190
rect 2828 26114 2884 26124
rect 3164 26178 3444 26180
rect 3164 26126 3390 26178
rect 3442 26126 3444 26178
rect 3164 26124 3444 26126
rect 3164 25508 3220 26124
rect 3388 26114 3444 26124
rect 2828 25452 3220 25508
rect 2716 25396 2772 25406
rect 2044 25394 2772 25396
rect 2044 25342 2718 25394
rect 2770 25342 2772 25394
rect 2044 25340 2772 25342
rect 2044 24946 2100 25340
rect 2716 25330 2772 25340
rect 2044 24894 2046 24946
rect 2098 24894 2100 24946
rect 2044 24882 2100 24894
rect 2828 24946 2884 25452
rect 2828 24894 2830 24946
rect 2882 24894 2884 24946
rect 2828 24882 2884 24894
rect 3052 23828 3108 23838
rect 3052 23734 3108 23772
rect 3052 22260 3108 22270
rect 3052 22166 3108 22204
rect 3612 22148 3668 28924
rect 3948 28532 4004 28542
rect 3836 27860 3892 27870
rect 3724 26180 3780 26190
rect 3724 25620 3780 26124
rect 3724 25554 3780 25564
rect 3836 25618 3892 27804
rect 3948 27076 4004 28476
rect 4284 27748 4340 29484
rect 4508 29474 4564 29484
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4956 28756 5012 28766
rect 4956 28662 5012 28700
rect 4844 28644 4900 28654
rect 4844 28550 4900 28588
rect 4284 27682 4340 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3948 26290 4004 27020
rect 3948 26238 3950 26290
rect 4002 26238 4004 26290
rect 3948 26226 4004 26238
rect 4060 27186 4116 27198
rect 4060 27134 4062 27186
rect 4114 27134 4116 27186
rect 4060 26292 4116 27134
rect 4508 26292 4564 26302
rect 4060 26290 4564 26292
rect 4060 26238 4510 26290
rect 4562 26238 4564 26290
rect 4060 26236 4564 26238
rect 4508 26226 4564 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3836 25566 3838 25618
rect 3890 25566 3892 25618
rect 3836 25554 3892 25566
rect 4508 25620 4564 25630
rect 4508 25526 4564 25564
rect 5180 24722 5236 30268
rect 6636 30258 6692 30268
rect 11228 30324 11284 30334
rect 11228 30230 11284 30268
rect 5292 30100 5348 30110
rect 5292 29650 5348 30044
rect 7644 30100 7700 30110
rect 9884 30100 9940 30110
rect 7644 30006 7700 30044
rect 9212 30098 9940 30100
rect 9212 30046 9886 30098
rect 9938 30046 9940 30098
rect 9212 30044 9940 30046
rect 5292 29598 5294 29650
rect 5346 29598 5348 29650
rect 5292 29586 5348 29598
rect 8540 29538 8596 29550
rect 8540 29486 8542 29538
rect 8594 29486 8596 29538
rect 6188 29316 6244 29326
rect 5740 28644 5796 28654
rect 5740 28550 5796 28588
rect 5516 27972 5572 27982
rect 5404 27916 5516 27972
rect 5292 27860 5348 27870
rect 5292 27766 5348 27804
rect 5404 25732 5460 27916
rect 5516 27906 5572 27916
rect 5740 27860 5796 27870
rect 5516 27076 5572 27086
rect 5740 27076 5796 27804
rect 5572 27020 5796 27076
rect 6188 27074 6244 29260
rect 7532 29316 7588 29326
rect 7532 29222 7588 29260
rect 6748 28644 6804 28654
rect 6748 28550 6804 28588
rect 7420 28644 7476 28654
rect 6972 28530 7028 28542
rect 6972 28478 6974 28530
rect 7026 28478 7028 28530
rect 6636 27972 6692 27982
rect 6636 27878 6692 27916
rect 6188 27022 6190 27074
rect 6242 27022 6244 27074
rect 5516 26982 5572 27020
rect 5516 25732 5572 25742
rect 5404 25730 5572 25732
rect 5404 25678 5518 25730
rect 5570 25678 5572 25730
rect 5404 25676 5572 25678
rect 5516 25666 5572 25676
rect 5180 24670 5182 24722
rect 5234 24670 5236 24722
rect 5180 24658 5236 24670
rect 5628 24722 5684 27020
rect 6188 27010 6244 27022
rect 6300 27076 6356 27086
rect 6300 25394 6356 27020
rect 6972 26514 7028 28478
rect 6972 26462 6974 26514
rect 7026 26462 7028 26514
rect 6972 26450 7028 26462
rect 7420 26068 7476 28588
rect 7868 28642 7924 28654
rect 8428 28644 8484 28654
rect 7868 28590 7870 28642
rect 7922 28590 7924 28642
rect 7868 27860 7924 28590
rect 7868 27794 7924 27804
rect 7980 28642 8484 28644
rect 7980 28590 8430 28642
rect 8482 28590 8484 28642
rect 7980 28588 8484 28590
rect 7644 27748 7700 27758
rect 7644 26514 7700 27692
rect 7980 27746 8036 28588
rect 8428 28578 8484 28588
rect 7980 27694 7982 27746
rect 8034 27694 8036 27746
rect 7980 27682 8036 27694
rect 8540 27748 8596 29486
rect 8540 27682 8596 27692
rect 9212 27298 9268 30044
rect 9884 30034 9940 30044
rect 9996 29428 10052 29438
rect 9212 27246 9214 27298
rect 9266 27246 9268 27298
rect 9212 27234 9268 27246
rect 9324 27860 9380 27870
rect 9324 27076 9380 27804
rect 9548 27746 9604 27758
rect 9548 27694 9550 27746
rect 9602 27694 9604 27746
rect 9548 27412 9604 27694
rect 9884 27748 9940 27758
rect 9884 27654 9940 27692
rect 9548 27346 9604 27356
rect 9324 27074 9828 27076
rect 9324 27022 9326 27074
rect 9378 27022 9828 27074
rect 9324 27020 9828 27022
rect 7644 26462 7646 26514
rect 7698 26462 7700 26514
rect 7644 26450 7700 26462
rect 8652 26850 8708 26862
rect 8652 26798 8654 26850
rect 8706 26798 8708 26850
rect 8652 26402 8708 26798
rect 8652 26350 8654 26402
rect 8706 26350 8708 26402
rect 8652 26338 8708 26350
rect 8876 26290 8932 26302
rect 8876 26238 8878 26290
rect 8930 26238 8932 26290
rect 7420 25620 7476 26012
rect 8316 26178 8372 26190
rect 8316 26126 8318 26178
rect 8370 26126 8372 26178
rect 8316 26068 8372 26126
rect 8876 26180 8932 26238
rect 8876 26114 8932 26124
rect 8316 26002 8372 26012
rect 8652 26068 8708 26078
rect 7420 25554 7476 25564
rect 8652 25506 8708 26012
rect 8652 25454 8654 25506
rect 8706 25454 8708 25506
rect 8652 25442 8708 25454
rect 9212 25508 9268 25518
rect 9324 25508 9380 27020
rect 9772 26852 9828 27020
rect 9996 27074 10052 29372
rect 11452 29428 11508 31838
rect 18060 31890 18564 31892
rect 18060 31838 18510 31890
rect 18562 31838 18564 31890
rect 18060 31836 18564 31838
rect 11452 29362 11508 29372
rect 11564 31668 11620 31678
rect 11564 28866 11620 31612
rect 12460 31668 12516 31678
rect 16604 31668 16660 31678
rect 12460 31574 12516 31612
rect 16492 31612 16604 31668
rect 14140 31108 14196 31118
rect 14140 31014 14196 31052
rect 12908 30882 12964 30894
rect 12908 30830 12910 30882
rect 12962 30830 12964 30882
rect 11564 28814 11566 28866
rect 11618 28814 11620 28866
rect 11564 28802 11620 28814
rect 12124 30324 12180 30334
rect 10780 28418 10836 28430
rect 10780 28366 10782 28418
rect 10834 28366 10836 28418
rect 10780 28082 10836 28366
rect 10780 28030 10782 28082
rect 10834 28030 10836 28082
rect 10780 28018 10836 28030
rect 9996 27022 9998 27074
rect 10050 27022 10052 27074
rect 9996 27010 10052 27022
rect 10780 27858 10836 27870
rect 10780 27806 10782 27858
rect 10834 27806 10836 27858
rect 10780 27748 10836 27806
rect 10780 27076 10836 27692
rect 10780 27010 10836 27020
rect 11564 27858 11620 27870
rect 11564 27806 11566 27858
rect 11618 27806 11620 27858
rect 9772 26402 9828 26796
rect 11564 26852 11620 27806
rect 11564 26786 11620 26796
rect 11900 27076 11956 27086
rect 9772 26350 9774 26402
rect 9826 26350 9828 26402
rect 9772 26338 9828 26350
rect 11004 26180 11060 26190
rect 9212 25506 9492 25508
rect 9212 25454 9214 25506
rect 9266 25454 9492 25506
rect 9212 25452 9492 25454
rect 9212 25442 9268 25452
rect 6300 25342 6302 25394
rect 6354 25342 6356 25394
rect 6300 25330 6356 25342
rect 6972 25284 7028 25294
rect 6972 24834 7028 25228
rect 9324 25284 9380 25294
rect 9324 25190 9380 25228
rect 6972 24782 6974 24834
rect 7026 24782 7028 24834
rect 6972 24770 7028 24782
rect 9436 24836 9492 25452
rect 10108 25282 10164 25294
rect 10108 25230 10110 25282
rect 10162 25230 10164 25282
rect 10108 24948 10164 25230
rect 10108 24882 10164 24892
rect 5628 24670 5630 24722
rect 5682 24670 5684 24722
rect 5628 24658 5684 24670
rect 7980 24724 8036 24734
rect 7980 24610 8036 24668
rect 9436 24722 9492 24780
rect 10220 24836 10276 24846
rect 10276 24780 10500 24836
rect 10220 24770 10276 24780
rect 9436 24670 9438 24722
rect 9490 24670 9492 24722
rect 9436 24658 9492 24670
rect 10108 24724 10164 24734
rect 10108 24630 10164 24668
rect 7980 24558 7982 24610
rect 8034 24558 8036 24610
rect 7980 24546 8036 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 6748 24164 6804 24174
rect 4060 24052 4116 24062
rect 4060 23958 4116 23996
rect 6748 24050 6804 24108
rect 6748 23998 6750 24050
rect 6802 23998 6804 24050
rect 6748 23986 6804 23998
rect 9996 23940 10052 23950
rect 9996 23846 10052 23884
rect 10444 23938 10500 24780
rect 11004 24052 11060 26124
rect 11900 24164 11956 27020
rect 12124 25508 12180 30268
rect 12572 29316 12628 29326
rect 12236 29314 12628 29316
rect 12236 29262 12574 29314
rect 12626 29262 12628 29314
rect 12236 29260 12628 29262
rect 12236 27858 12292 29260
rect 12572 29250 12628 29260
rect 12236 27806 12238 27858
rect 12290 27806 12292 27858
rect 12236 27794 12292 27806
rect 12236 26964 12292 26974
rect 12236 26870 12292 26908
rect 12796 26852 12852 26862
rect 12572 26180 12628 26190
rect 12348 25508 12404 25518
rect 12124 25506 12404 25508
rect 12124 25454 12350 25506
rect 12402 25454 12404 25506
rect 12124 25452 12404 25454
rect 12348 25442 12404 25452
rect 12572 24946 12628 26124
rect 12796 25506 12852 26796
rect 12908 26068 12964 30830
rect 14476 30210 14532 30222
rect 14476 30158 14478 30210
rect 14530 30158 14532 30210
rect 13580 29540 13636 29550
rect 13020 29538 13636 29540
rect 13020 29486 13582 29538
rect 13634 29486 13636 29538
rect 13020 29484 13636 29486
rect 13020 27298 13076 29484
rect 13580 29474 13636 29484
rect 14476 29428 14532 30158
rect 14476 29362 14532 29372
rect 14924 30210 14980 30222
rect 14924 30158 14926 30210
rect 14978 30158 14980 30210
rect 14924 29316 14980 30158
rect 16380 29540 16436 29550
rect 15484 29538 16436 29540
rect 15484 29486 16382 29538
rect 16434 29486 16436 29538
rect 15484 29484 16436 29486
rect 15372 29316 15428 29326
rect 14924 29314 15428 29316
rect 14924 29262 15374 29314
rect 15426 29262 15428 29314
rect 14924 29260 15428 29262
rect 15372 29250 15428 29260
rect 15036 28756 15092 28766
rect 15036 28754 15204 28756
rect 15036 28702 15038 28754
rect 15090 28702 15204 28754
rect 15036 28700 15204 28702
rect 15036 28690 15092 28700
rect 13692 28532 13748 28542
rect 13020 27246 13022 27298
rect 13074 27246 13076 27298
rect 13020 27234 13076 27246
rect 13468 28530 13748 28532
rect 13468 28478 13694 28530
rect 13746 28478 13748 28530
rect 13468 28476 13748 28478
rect 13468 26516 13524 28476
rect 13692 28466 13748 28476
rect 14476 27972 14532 27982
rect 14140 27970 14532 27972
rect 14140 27918 14478 27970
rect 14530 27918 14532 27970
rect 14140 27916 14532 27918
rect 14140 27186 14196 27916
rect 14476 27906 14532 27916
rect 15148 27860 15204 28700
rect 15484 28532 15540 29484
rect 16380 29474 16436 29484
rect 16268 28868 16324 28878
rect 16492 28868 16548 31612
rect 16604 31602 16660 31612
rect 17388 31668 17444 31678
rect 17388 31574 17444 31612
rect 17164 31108 17220 31118
rect 17220 31052 17332 31108
rect 17164 31042 17220 31052
rect 17164 29988 17220 29998
rect 16268 28866 16548 28868
rect 16268 28814 16270 28866
rect 16322 28814 16548 28866
rect 16268 28812 16548 28814
rect 16716 29986 17220 29988
rect 16716 29934 17166 29986
rect 17218 29934 17220 29986
rect 16716 29932 17220 29934
rect 16268 28802 16324 28812
rect 15260 28476 15540 28532
rect 16380 28532 16436 28542
rect 15260 28082 15316 28476
rect 15260 28030 15262 28082
rect 15314 28030 15316 28082
rect 15260 28018 15316 28030
rect 15372 27916 16324 27972
rect 15372 27860 15428 27916
rect 15148 27804 15428 27860
rect 15708 27748 15764 27758
rect 14140 27134 14142 27186
rect 14194 27134 14196 27186
rect 14140 27122 14196 27134
rect 15596 27746 15764 27748
rect 15596 27694 15710 27746
rect 15762 27694 15764 27746
rect 15596 27692 15764 27694
rect 13916 27076 13972 27086
rect 13916 26964 13972 27020
rect 14476 26964 14532 26974
rect 13916 26962 14532 26964
rect 13916 26910 14478 26962
rect 14530 26910 14532 26962
rect 13916 26908 14532 26910
rect 14476 26898 14532 26908
rect 14812 26964 14868 26974
rect 14812 26870 14868 26908
rect 12908 26002 12964 26012
rect 13132 26460 13524 26516
rect 15484 26850 15540 26862
rect 15484 26798 15486 26850
rect 15538 26798 15540 26850
rect 12796 25454 12798 25506
rect 12850 25454 12852 25506
rect 12796 25442 12852 25454
rect 12572 24894 12574 24946
rect 12626 24894 12628 24946
rect 12572 24882 12628 24894
rect 13132 24946 13188 26460
rect 14812 26292 14868 26302
rect 14812 26198 14868 26236
rect 15148 26180 15204 26190
rect 15148 26086 15204 26124
rect 15484 26178 15540 26798
rect 15596 26292 15652 27692
rect 15708 27682 15764 27692
rect 15932 27074 15988 27086
rect 15932 27022 15934 27074
rect 15986 27022 15988 27074
rect 15932 26404 15988 27022
rect 16268 26908 16324 27916
rect 16380 27074 16436 28476
rect 16716 28082 16772 29932
rect 17164 29922 17220 29932
rect 16716 28030 16718 28082
rect 16770 28030 16772 28082
rect 16716 28018 16772 28030
rect 17052 28418 17108 28430
rect 17052 28366 17054 28418
rect 17106 28366 17108 28418
rect 16828 27748 16884 27758
rect 16828 27654 16884 27692
rect 16380 27022 16382 27074
rect 16434 27022 16436 27074
rect 16380 27010 16436 27022
rect 16268 26852 16436 26908
rect 15932 26348 16324 26404
rect 15596 26226 15652 26236
rect 15484 26126 15486 26178
rect 15538 26126 15540 26178
rect 14028 25732 14084 25742
rect 13356 25508 13412 25518
rect 13132 24894 13134 24946
rect 13186 24894 13188 24946
rect 13132 24882 13188 24894
rect 13244 25396 13300 25406
rect 13244 24946 13300 25340
rect 13244 24894 13246 24946
rect 13298 24894 13300 24946
rect 13244 24882 13300 24894
rect 11004 23958 11060 23996
rect 11788 24108 11900 24164
rect 10444 23886 10446 23938
rect 10498 23886 10500 23938
rect 10444 23874 10500 23886
rect 6412 23828 6468 23838
rect 6188 23826 6468 23828
rect 6188 23774 6414 23826
rect 6466 23774 6468 23826
rect 6188 23772 6468 23774
rect 4060 23268 4116 23278
rect 4060 23174 4116 23212
rect 5180 23044 5236 23054
rect 5180 22950 5236 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4060 22484 4116 22494
rect 4060 22390 4116 22428
rect 5516 22372 5572 22382
rect 3612 22082 3668 22092
rect 5292 22370 5572 22372
rect 5292 22318 5518 22370
rect 5570 22318 5572 22370
rect 5292 22316 5572 22318
rect 4060 21924 4116 21934
rect 2156 21810 2212 21822
rect 2156 21758 2158 21810
rect 2210 21758 2212 21810
rect 1596 21362 1652 21374
rect 1596 21310 1598 21362
rect 1650 21310 1652 21362
rect 1596 16884 1652 21310
rect 2044 19124 2100 19134
rect 2044 19030 2100 19068
rect 1708 19010 1764 19022
rect 1708 18958 1710 19010
rect 1762 18958 1764 19010
rect 1708 18900 1764 18958
rect 1764 18844 1876 18900
rect 1708 18834 1764 18844
rect 1820 18674 1876 18844
rect 1820 18622 1822 18674
rect 1874 18622 1876 18674
rect 1820 18610 1876 18622
rect 2156 18004 2212 21758
rect 3052 21364 3108 21374
rect 3052 20690 3108 21308
rect 4060 20914 4116 21868
rect 4732 21588 4788 21598
rect 5292 21588 5348 22316
rect 5516 22306 5572 22316
rect 6076 22370 6132 22382
rect 6076 22318 6078 22370
rect 6130 22318 6132 22370
rect 6076 21924 6132 22318
rect 6076 21858 6132 21868
rect 6188 21810 6244 23772
rect 6412 23762 6468 23772
rect 9212 23828 9268 23838
rect 6972 23716 7028 23726
rect 6860 23714 7028 23716
rect 6860 23662 6974 23714
rect 7026 23662 7028 23714
rect 6860 23660 7028 23662
rect 6860 22260 6916 23660
rect 6972 23650 7028 23660
rect 7644 23714 7700 23726
rect 7644 23662 7646 23714
rect 7698 23662 7700 23714
rect 6972 23380 7028 23390
rect 6972 23266 7028 23324
rect 6972 23214 6974 23266
rect 7026 23214 7028 23266
rect 6972 23202 7028 23214
rect 6860 22194 6916 22204
rect 6188 21758 6190 21810
rect 6242 21758 6244 21810
rect 6188 21746 6244 21758
rect 4732 21494 4788 21532
rect 5068 21586 5348 21588
rect 5068 21534 5294 21586
rect 5346 21534 5348 21586
rect 5068 21532 5348 21534
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4060 20862 4062 20914
rect 4114 20862 4116 20914
rect 4060 20850 4116 20862
rect 3052 20638 3054 20690
rect 3106 20638 3108 20690
rect 3052 20626 3108 20638
rect 5068 20244 5124 21532
rect 5292 21522 5348 21532
rect 6860 21588 6916 21598
rect 5404 21364 5460 21374
rect 5404 21270 5460 21308
rect 5628 20690 5684 20702
rect 5628 20638 5630 20690
rect 5682 20638 5684 20690
rect 5628 20188 5684 20638
rect 3276 20132 3332 20142
rect 3276 20038 3332 20076
rect 4172 20132 5124 20188
rect 5180 20132 5684 20188
rect 5964 20690 6020 20702
rect 5964 20638 5966 20690
rect 6018 20638 6020 20690
rect 5964 20188 6020 20638
rect 5964 20132 6132 20188
rect 6748 20132 6804 20142
rect 4060 20020 4116 20030
rect 4172 20020 4228 20132
rect 4396 20020 4452 20030
rect 5180 20020 5236 20132
rect 5964 20066 6020 20076
rect 4060 20018 4228 20020
rect 4060 19966 4062 20018
rect 4114 19966 4228 20018
rect 4060 19964 4228 19966
rect 4060 19954 4116 19964
rect 3612 19908 3668 19918
rect 3612 19906 3892 19908
rect 3612 19854 3614 19906
rect 3666 19854 3892 19906
rect 3612 19852 3892 19854
rect 3612 19842 3668 19852
rect 3052 19122 3108 19134
rect 3052 19070 3054 19122
rect 3106 19070 3108 19122
rect 2044 17948 2212 18004
rect 2268 18450 2324 18462
rect 2268 18398 2270 18450
rect 2322 18398 2324 18450
rect 1932 17554 1988 17566
rect 1932 17502 1934 17554
rect 1986 17502 1988 17554
rect 1596 16828 1764 16884
rect 1596 16660 1652 16670
rect 1596 16566 1652 16604
rect 1708 15988 1764 16828
rect 1932 16100 1988 17502
rect 1932 16006 1988 16044
rect 1820 15988 1876 15998
rect 1708 15932 1820 15988
rect 1820 15922 1876 15932
rect 2044 15874 2100 17948
rect 2156 17778 2212 17790
rect 2156 17726 2158 17778
rect 2210 17726 2212 17778
rect 2156 17106 2212 17726
rect 2156 17054 2158 17106
rect 2210 17054 2212 17106
rect 2156 17042 2212 17054
rect 2044 15822 2046 15874
rect 2098 15822 2100 15874
rect 2044 15810 2100 15822
rect 2268 16884 2324 18398
rect 2268 15314 2324 16828
rect 2716 18450 2772 18462
rect 2716 18398 2718 18450
rect 2770 18398 2772 18450
rect 2268 15262 2270 15314
rect 2322 15262 2324 15314
rect 2268 13746 2324 15262
rect 2380 16660 2436 16670
rect 2380 14418 2436 16604
rect 2716 16548 2772 18398
rect 3052 18452 3108 19070
rect 3052 18386 3108 18396
rect 3052 18228 3108 18238
rect 3052 17554 3108 18172
rect 3052 17502 3054 17554
rect 3106 17502 3108 17554
rect 3052 17490 3108 17502
rect 3836 16660 3892 19852
rect 3948 19346 4004 19358
rect 3948 19294 3950 19346
rect 4002 19294 4004 19346
rect 3948 19236 4004 19294
rect 3948 19170 4004 19180
rect 3948 17780 4004 17790
rect 3948 17686 4004 17724
rect 4060 16884 4116 16894
rect 4172 16884 4228 19964
rect 4284 20018 4452 20020
rect 4284 19966 4398 20018
rect 4450 19966 4452 20018
rect 4284 19964 4452 19966
rect 4284 17780 4340 19964
rect 4396 19954 4452 19964
rect 4956 19964 5236 20020
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4956 18674 5012 19964
rect 4956 18622 4958 18674
rect 5010 18622 5012 18674
rect 4956 18610 5012 18622
rect 6076 19348 6132 20132
rect 6076 19234 6132 19292
rect 6300 20130 6804 20132
rect 6300 20078 6750 20130
rect 6802 20078 6804 20130
rect 6300 20076 6804 20078
rect 6300 19346 6356 20076
rect 6748 20066 6804 20076
rect 6300 19294 6302 19346
rect 6354 19294 6356 19346
rect 6300 19282 6356 19294
rect 6076 19182 6078 19234
rect 6130 19182 6132 19234
rect 5516 18452 5572 18462
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5516 17890 5572 18396
rect 5740 18228 5796 18238
rect 5740 18134 5796 18172
rect 5516 17838 5518 17890
rect 5570 17838 5572 17890
rect 5516 17826 5572 17838
rect 4284 17714 4340 17724
rect 4116 16828 4228 16884
rect 4732 16996 4788 17006
rect 4732 16882 4788 16940
rect 4732 16830 4734 16882
rect 4786 16830 4788 16882
rect 4060 16818 4116 16828
rect 4732 16818 4788 16830
rect 5068 16884 5124 16894
rect 6076 16884 6132 19182
rect 6636 19124 6692 19134
rect 6188 19122 6692 19124
rect 6188 19070 6638 19122
rect 6690 19070 6692 19122
rect 6188 19068 6692 19070
rect 6188 17106 6244 19068
rect 6636 19058 6692 19068
rect 6300 17444 6356 17454
rect 6300 17350 6356 17388
rect 6188 17054 6190 17106
rect 6242 17054 6244 17106
rect 6188 17042 6244 17054
rect 6076 16828 6244 16884
rect 5068 16790 5124 16828
rect 5404 16660 5460 16670
rect 3836 16604 5012 16660
rect 2716 16482 2772 16492
rect 3500 16548 3556 16558
rect 2940 16212 2996 16222
rect 2716 15988 2772 15998
rect 2716 15894 2772 15932
rect 2380 14366 2382 14418
rect 2434 14366 2436 14418
rect 2380 14354 2436 14366
rect 2716 15314 2772 15326
rect 2716 15262 2718 15314
rect 2770 15262 2772 15314
rect 2716 14196 2772 15262
rect 2716 14130 2772 14140
rect 2268 13694 2270 13746
rect 2322 13694 2324 13746
rect 2268 13682 2324 13694
rect 2940 13746 2996 16156
rect 3500 14642 3556 16492
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3836 16212 3892 16222
rect 3836 16118 3892 16156
rect 4956 15538 5012 16604
rect 5404 16658 6132 16660
rect 5404 16606 5406 16658
rect 5458 16606 6132 16658
rect 5404 16604 6132 16606
rect 5404 16594 5460 16604
rect 5964 15988 6020 15998
rect 4956 15486 4958 15538
rect 5010 15486 5012 15538
rect 4956 15474 5012 15486
rect 5404 15986 6020 15988
rect 5404 15934 5966 15986
rect 6018 15934 6020 15986
rect 5404 15932 6020 15934
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 3500 14590 3502 14642
rect 3554 14590 3556 14642
rect 3500 14578 3556 14590
rect 2940 13694 2942 13746
rect 2994 13694 2996 13746
rect 2940 13682 2996 13694
rect 3612 14196 3668 14206
rect 3612 13074 3668 14140
rect 5404 13970 5460 15932
rect 5964 15922 6020 15932
rect 5740 15092 5796 15102
rect 5740 14998 5796 15036
rect 6076 14418 6132 16604
rect 6188 16100 6244 16828
rect 6188 15988 6244 16044
rect 6300 15988 6356 15998
rect 6188 15986 6356 15988
rect 6188 15934 6302 15986
rect 6354 15934 6356 15986
rect 6188 15932 6356 15934
rect 6300 15204 6356 15932
rect 6860 15204 6916 21532
rect 7644 20914 7700 23662
rect 7980 23042 8036 23054
rect 7980 22990 7982 23042
rect 8034 22990 8036 23042
rect 7980 22932 8036 22990
rect 7980 22866 8036 22876
rect 9212 22594 9268 23772
rect 11340 23826 11396 23838
rect 11340 23774 11342 23826
rect 11394 23774 11396 23826
rect 9436 23268 9492 23278
rect 9436 23174 9492 23212
rect 10220 23266 10276 23278
rect 10220 23214 10222 23266
rect 10274 23214 10276 23266
rect 9212 22542 9214 22594
rect 9266 22542 9268 22594
rect 9212 22530 9268 22542
rect 9884 23044 9940 23054
rect 8540 22484 8596 22494
rect 7644 20862 7646 20914
rect 7698 20862 7700 20914
rect 7644 20850 7700 20862
rect 8428 21586 8484 21598
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 7980 20804 8036 20814
rect 7420 20692 7476 20702
rect 7420 20598 7476 20636
rect 7196 20244 7252 20254
rect 6972 19348 7028 19358
rect 6972 19254 7028 19292
rect 7196 19234 7252 20188
rect 7980 20244 8036 20748
rect 7980 20178 8036 20188
rect 7980 19906 8036 19918
rect 7980 19854 7982 19906
rect 8034 19854 8036 19906
rect 7196 19182 7198 19234
rect 7250 19182 7252 19234
rect 7196 19170 7252 19182
rect 7532 19794 7588 19806
rect 7532 19742 7534 19794
rect 7586 19742 7588 19794
rect 6972 18564 7028 18574
rect 7532 18564 7588 19742
rect 7980 19348 8036 19854
rect 8316 19908 8372 19918
rect 8316 19814 8372 19852
rect 7980 19282 8036 19292
rect 7756 19236 7812 19246
rect 7756 19142 7812 19180
rect 8428 19124 8484 21534
rect 8540 20802 8596 22428
rect 9324 22372 9380 22382
rect 9100 22370 9380 22372
rect 9100 22318 9326 22370
rect 9378 22318 9380 22370
rect 9100 22316 9380 22318
rect 8540 20750 8542 20802
rect 8594 20750 8596 20802
rect 8540 20738 8596 20750
rect 8652 22146 8708 22158
rect 8652 22094 8654 22146
rect 8706 22094 8708 22146
rect 8652 20130 8708 22094
rect 9100 21586 9156 22316
rect 9324 22306 9380 22316
rect 9884 22370 9940 22988
rect 9884 22318 9886 22370
rect 9938 22318 9940 22370
rect 9884 22306 9940 22318
rect 10220 21812 10276 23214
rect 11340 22036 11396 23774
rect 11340 21970 11396 21980
rect 10220 21746 10276 21756
rect 9100 21534 9102 21586
rect 9154 21534 9156 21586
rect 9100 20804 9156 21534
rect 8652 20078 8654 20130
rect 8706 20078 8708 20130
rect 8652 20066 8708 20078
rect 8988 20692 9044 20702
rect 8988 20130 9044 20636
rect 9100 20188 9156 20748
rect 9996 21700 10052 21710
rect 9996 21586 10052 21644
rect 9996 21534 9998 21586
rect 10050 21534 10052 21586
rect 9996 20804 10052 21534
rect 11004 21698 11060 21710
rect 11004 21646 11006 21698
rect 11058 21646 11060 21698
rect 10220 21476 10276 21486
rect 10220 21474 10948 21476
rect 10220 21422 10222 21474
rect 10274 21422 10948 21474
rect 10220 21420 10948 21422
rect 10220 21410 10276 21420
rect 9996 20738 10052 20748
rect 10892 20690 10948 21420
rect 11004 21028 11060 21646
rect 11788 21700 11844 24108
rect 11900 24070 11956 24108
rect 12572 24052 12628 24062
rect 12012 23156 12068 23166
rect 12460 23156 12516 23166
rect 11788 21634 11844 21644
rect 11900 21812 11956 21822
rect 11004 20962 11060 20972
rect 11900 20914 11956 21756
rect 12012 21474 12068 23100
rect 12236 23154 12516 23156
rect 12236 23102 12462 23154
rect 12514 23102 12516 23154
rect 12236 23100 12516 23102
rect 12012 21422 12014 21474
rect 12066 21422 12068 21474
rect 12012 21410 12068 21422
rect 12124 21700 12180 21710
rect 11900 20862 11902 20914
rect 11954 20862 11956 20914
rect 11900 20850 11956 20862
rect 12124 20916 12180 21644
rect 12124 20802 12180 20860
rect 12124 20750 12126 20802
rect 12178 20750 12180 20802
rect 12124 20738 12180 20750
rect 10892 20638 10894 20690
rect 10946 20638 10948 20690
rect 10892 20626 10948 20638
rect 9996 20580 10052 20590
rect 9100 20132 9828 20188
rect 8988 20078 8990 20130
rect 9042 20078 9044 20130
rect 8988 20066 9044 20078
rect 9772 20130 9828 20132
rect 9772 20078 9774 20130
rect 9826 20078 9828 20130
rect 9772 20066 9828 20078
rect 6972 18562 7588 18564
rect 6972 18510 6974 18562
rect 7026 18510 7588 18562
rect 6972 18508 7588 18510
rect 7980 19068 8484 19124
rect 6972 18498 7028 18508
rect 7980 18338 8036 19068
rect 9996 18562 10052 20524
rect 11676 20580 11732 20590
rect 11676 20486 11732 20524
rect 10108 19908 10164 19918
rect 10108 19122 10164 19852
rect 10108 19070 10110 19122
rect 10162 19070 10164 19122
rect 10108 19058 10164 19070
rect 11228 19236 11284 19246
rect 9996 18510 9998 18562
rect 10050 18510 10052 18562
rect 9996 18498 10052 18510
rect 10892 19010 10948 19022
rect 10892 18958 10894 19010
rect 10946 18958 10948 19010
rect 7980 18286 7982 18338
rect 8034 18286 8036 18338
rect 7980 18274 8036 18286
rect 8540 17666 8596 17678
rect 8540 17614 8542 17666
rect 8594 17614 8596 17666
rect 7196 16996 7252 17006
rect 6972 15204 7028 15214
rect 6860 15202 7028 15204
rect 6860 15150 6974 15202
rect 7026 15150 7028 15202
rect 6860 15148 7028 15150
rect 6300 15138 6356 15148
rect 6972 15138 7028 15148
rect 6076 14366 6078 14418
rect 6130 14366 6132 14418
rect 6076 14354 6132 14366
rect 5404 13918 5406 13970
rect 5458 13918 5460 13970
rect 5404 13906 5460 13918
rect 7196 13634 7252 16940
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 8428 16212 8484 16830
rect 8428 16146 8484 16156
rect 7420 16100 7476 16110
rect 7420 14642 7476 16044
rect 8540 16100 8596 17614
rect 9212 17668 9268 17678
rect 9436 17668 9492 17678
rect 9212 17666 9492 17668
rect 9212 17614 9214 17666
rect 9266 17614 9438 17666
rect 9490 17614 9492 17666
rect 9212 17612 9492 17614
rect 9212 17602 9268 17612
rect 8876 16884 8932 16894
rect 8876 16790 8932 16828
rect 9436 16884 9492 17612
rect 9436 16790 9492 16828
rect 9884 17666 9940 17678
rect 9884 17614 9886 17666
rect 9938 17614 9940 17666
rect 8540 16034 8596 16044
rect 9884 15988 9940 17614
rect 10892 16996 10948 18958
rect 11228 18338 11284 19180
rect 12236 19236 12292 23100
rect 12460 23090 12516 23100
rect 12348 22146 12404 22158
rect 12348 22094 12350 22146
rect 12402 22094 12404 22146
rect 12348 20916 12404 22094
rect 12572 21810 12628 23996
rect 12908 23826 12964 23838
rect 12908 23774 12910 23826
rect 12962 23774 12964 23826
rect 12908 23044 12964 23774
rect 13132 23156 13188 23166
rect 13356 23156 13412 25452
rect 13580 25396 13636 25406
rect 13580 25302 13636 25340
rect 13468 24948 13524 24958
rect 13468 24050 13524 24892
rect 14028 24946 14084 25676
rect 14924 25620 14980 25630
rect 14924 25526 14980 25564
rect 14028 24894 14030 24946
rect 14082 24894 14084 24946
rect 14028 24882 14084 24894
rect 15484 25284 15540 26126
rect 15820 26180 15876 26190
rect 15820 25284 15876 26124
rect 16156 26178 16212 26190
rect 16156 26126 16158 26178
rect 16210 26126 16212 26178
rect 15932 25284 15988 25294
rect 15484 25282 15988 25284
rect 15484 25230 15486 25282
rect 15538 25230 15934 25282
rect 15986 25230 15988 25282
rect 15484 25228 15988 25230
rect 13468 23998 13470 24050
rect 13522 23998 13524 24050
rect 13468 23986 13524 23998
rect 13692 24052 13748 24062
rect 13692 23938 13748 23996
rect 15484 24052 15540 25228
rect 15932 25218 15988 25228
rect 15484 23986 15540 23996
rect 15932 24050 15988 24062
rect 15932 23998 15934 24050
rect 15986 23998 15988 24050
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 13692 23874 13748 23886
rect 14924 23826 14980 23838
rect 14924 23774 14926 23826
rect 14978 23774 14980 23826
rect 13132 23154 13412 23156
rect 13132 23102 13134 23154
rect 13186 23102 13358 23154
rect 13410 23102 13412 23154
rect 13132 23100 13412 23102
rect 13132 23090 13188 23100
rect 13020 23044 13076 23054
rect 12908 22988 13020 23044
rect 13020 22372 13076 22988
rect 13020 22316 13300 22372
rect 13020 22146 13076 22158
rect 13020 22094 13022 22146
rect 13074 22094 13076 22146
rect 13020 21924 13076 22094
rect 13020 21858 13076 21868
rect 12572 21758 12574 21810
rect 12626 21758 12628 21810
rect 12572 21746 12628 21758
rect 12572 20916 12628 20926
rect 12348 20914 12628 20916
rect 12348 20862 12574 20914
rect 12626 20862 12628 20914
rect 12348 20860 12628 20862
rect 12572 20850 12628 20860
rect 12796 20916 12852 20926
rect 12796 20802 12852 20860
rect 12796 20750 12798 20802
rect 12850 20750 12852 20802
rect 12796 20738 12852 20750
rect 12460 20020 12516 20030
rect 12460 19458 12516 19964
rect 13244 20020 13300 22316
rect 13356 21586 13412 23100
rect 13804 23156 13860 23166
rect 13804 23062 13860 23100
rect 13580 23044 13636 23054
rect 13580 22482 13636 22988
rect 13580 22430 13582 22482
rect 13634 22430 13636 22482
rect 13580 22418 13636 22430
rect 13804 22932 13860 22942
rect 13356 21534 13358 21586
rect 13410 21534 13412 21586
rect 13356 21522 13412 21534
rect 13804 21586 13860 22876
rect 14924 22596 14980 23774
rect 14924 22530 14980 22540
rect 15820 23044 15876 23054
rect 15372 22482 15428 22494
rect 15372 22430 15374 22482
rect 15426 22430 15428 22482
rect 14364 22260 14420 22270
rect 14364 22166 14420 22204
rect 13804 21534 13806 21586
rect 13858 21534 13860 21586
rect 13804 21522 13860 21534
rect 13916 22036 13972 22046
rect 13356 21028 13412 21038
rect 13356 20934 13412 20972
rect 13916 20578 13972 21980
rect 13916 20526 13918 20578
rect 13970 20526 13972 20578
rect 13916 20514 13972 20526
rect 14364 21924 14420 21934
rect 13244 19954 13300 19964
rect 12460 19406 12462 19458
rect 12514 19406 12516 19458
rect 12460 19394 12516 19406
rect 12236 19170 12292 19180
rect 11228 18286 11230 18338
rect 11282 18286 11284 18338
rect 11228 18274 11284 18286
rect 11452 19124 11508 19134
rect 10892 16930 10948 16940
rect 11116 17444 11172 17454
rect 10108 16882 10164 16894
rect 10108 16830 10110 16882
rect 10162 16830 10164 16882
rect 9884 15932 10052 15988
rect 7644 15876 7700 15886
rect 8428 15876 8484 15886
rect 7644 15874 8036 15876
rect 7644 15822 7646 15874
rect 7698 15822 8036 15874
rect 7644 15820 8036 15822
rect 7644 15810 7700 15820
rect 7980 15426 8036 15820
rect 8428 15874 9940 15876
rect 8428 15822 8430 15874
rect 8482 15822 9940 15874
rect 8428 15820 9940 15822
rect 8428 15810 8484 15820
rect 7980 15374 7982 15426
rect 8034 15374 8036 15426
rect 7980 15362 8036 15374
rect 9884 15426 9940 15820
rect 9884 15374 9886 15426
rect 9938 15374 9940 15426
rect 9884 15362 9940 15374
rect 9996 15316 10052 15932
rect 9996 15250 10052 15260
rect 7420 14590 7422 14642
rect 7474 14590 7476 14642
rect 7420 14578 7476 14590
rect 8428 15092 8484 15102
rect 8428 13858 8484 15036
rect 8428 13806 8430 13858
rect 8482 13806 8484 13858
rect 8428 13794 8484 13806
rect 7196 13582 7198 13634
rect 7250 13582 7252 13634
rect 7196 13570 7252 13582
rect 4956 13524 5012 13534
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 3612 13022 3614 13074
rect 3666 13022 3668 13074
rect 3612 13010 3668 13022
rect 4956 12850 5012 13468
rect 5964 13524 6020 13534
rect 5964 13430 6020 13468
rect 10108 13076 10164 16830
rect 10668 16212 10724 16222
rect 10220 15428 10276 15438
rect 10220 15334 10276 15372
rect 10668 13636 10724 16156
rect 10780 16098 10836 16110
rect 10780 16046 10782 16098
rect 10834 16046 10836 16098
rect 10780 14644 10836 16046
rect 11116 15426 11172 17388
rect 11340 16884 11396 16894
rect 11340 16098 11396 16828
rect 11340 16046 11342 16098
rect 11394 16046 11396 16098
rect 11340 16034 11396 16046
rect 11452 16100 11508 19068
rect 12572 19124 12628 19134
rect 12460 17442 12516 17454
rect 12460 17390 12462 17442
rect 12514 17390 12516 17442
rect 12348 16996 12404 17006
rect 11564 16100 11620 16110
rect 11452 16098 11620 16100
rect 11452 16046 11566 16098
rect 11618 16046 11620 16098
rect 11452 16044 11620 16046
rect 11564 16034 11620 16044
rect 11116 15374 11118 15426
rect 11170 15374 11172 15426
rect 11116 15362 11172 15374
rect 11452 15876 11508 15886
rect 11452 15428 11508 15820
rect 12124 15876 12180 15886
rect 12124 15782 12180 15820
rect 11452 15334 11508 15372
rect 11564 15316 11620 15326
rect 11452 14644 11508 14654
rect 10780 14642 11508 14644
rect 10780 14590 11454 14642
rect 11506 14590 11508 14642
rect 10780 14588 11508 14590
rect 11452 14578 11508 14588
rect 11452 13636 11508 13646
rect 10668 13634 11508 13636
rect 10668 13582 11454 13634
rect 11506 13582 11508 13634
rect 10668 13580 11508 13582
rect 11452 13570 11508 13580
rect 10108 13010 10164 13020
rect 11564 13074 11620 15260
rect 11676 15090 11732 15102
rect 11676 15038 11678 15090
rect 11730 15038 11732 15090
rect 11676 13636 11732 15038
rect 12348 14420 12404 16940
rect 12460 15764 12516 17390
rect 12572 17106 12628 19068
rect 13468 19124 13524 19134
rect 13468 19030 13524 19068
rect 13804 19124 13860 19134
rect 13804 19030 13860 19068
rect 12572 17054 12574 17106
rect 12626 17054 12628 17106
rect 12572 17042 12628 17054
rect 12684 18450 12740 18462
rect 13020 18452 13076 18462
rect 12684 18398 12686 18450
rect 12738 18398 12740 18450
rect 12684 16884 12740 18398
rect 12684 16818 12740 16828
rect 12908 18450 13076 18452
rect 12908 18398 13022 18450
rect 13074 18398 13076 18450
rect 12908 18396 13076 18398
rect 12908 16100 12964 18396
rect 13020 18386 13076 18396
rect 14140 18340 14196 18350
rect 14140 17554 14196 18284
rect 14140 17502 14142 17554
rect 14194 17502 14196 17554
rect 14140 17490 14196 17502
rect 12908 16034 12964 16044
rect 13020 17442 13076 17454
rect 13020 17390 13022 17442
rect 13074 17390 13076 17442
rect 13020 15876 13076 17390
rect 13356 17442 13412 17454
rect 13356 17390 13358 17442
rect 13410 17390 13412 17442
rect 13244 16884 13300 16894
rect 13244 16790 13300 16828
rect 13132 16660 13188 16670
rect 13132 16566 13188 16604
rect 13020 15810 13076 15820
rect 12460 15698 12516 15708
rect 13356 15652 13412 17390
rect 13916 16996 13972 17006
rect 13916 16882 13972 16940
rect 13916 16830 13918 16882
rect 13970 16830 13972 16882
rect 13916 16818 13972 16830
rect 12796 15596 13412 15652
rect 14140 16660 14196 16670
rect 12460 15426 12516 15438
rect 12460 15374 12462 15426
rect 12514 15374 12516 15426
rect 12460 14644 12516 15374
rect 12460 14578 12516 14588
rect 12460 14420 12516 14430
rect 12348 14418 12516 14420
rect 12348 14366 12462 14418
rect 12514 14366 12516 14418
rect 12348 14364 12516 14366
rect 12460 14354 12516 14364
rect 12796 13858 12852 15596
rect 14028 14644 14084 14654
rect 14028 14550 14084 14588
rect 12796 13806 12798 13858
rect 12850 13806 12852 13858
rect 12796 13794 12852 13806
rect 11676 13570 11732 13580
rect 12460 13636 12516 13646
rect 11564 13022 11566 13074
rect 11618 13022 11620 13074
rect 11564 13010 11620 13022
rect 4956 12798 4958 12850
rect 5010 12798 5012 12850
rect 4956 12786 5012 12798
rect 12460 12850 12516 13580
rect 12460 12798 12462 12850
rect 12514 12798 12516 12850
rect 12460 12786 12516 12798
rect 14140 12292 14196 16604
rect 14252 16100 14308 16110
rect 14252 13634 14308 16044
rect 14364 15986 14420 21868
rect 15372 21588 15428 22430
rect 15820 22482 15876 22988
rect 15820 22430 15822 22482
rect 15874 22430 15876 22482
rect 15820 22418 15876 22430
rect 15932 22484 15988 23998
rect 16156 23378 16212 26126
rect 16268 25506 16324 26348
rect 16268 25454 16270 25506
rect 16322 25454 16324 25506
rect 16268 25284 16324 25454
rect 16268 25218 16324 25228
rect 16268 24724 16324 24734
rect 16380 24724 16436 26852
rect 16716 26290 16772 26302
rect 16716 26238 16718 26290
rect 16770 26238 16772 26290
rect 16492 26178 16548 26190
rect 16492 26126 16494 26178
rect 16546 26126 16548 26178
rect 16492 25732 16548 26126
rect 16716 26180 16772 26238
rect 16716 26114 16772 26124
rect 16492 25666 16548 25676
rect 17052 25620 17108 28366
rect 17052 25554 17108 25564
rect 16828 25508 16884 25518
rect 16828 25414 16884 25452
rect 16268 24722 16436 24724
rect 16268 24670 16270 24722
rect 16322 24670 16436 24722
rect 16268 24668 16436 24670
rect 16940 25284 16996 25294
rect 16940 24724 16996 25228
rect 16268 24658 16324 24668
rect 16940 24630 16996 24668
rect 17164 24164 17220 24174
rect 17276 24164 17332 31052
rect 17948 30100 18004 30110
rect 17948 30006 18004 30044
rect 17500 29428 17556 29438
rect 17500 29334 17556 29372
rect 17948 29428 18004 29438
rect 18060 29428 18116 31836
rect 18508 31826 18564 31836
rect 20300 31892 20356 31902
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19628 30994 19684 31006
rect 19628 30942 19630 30994
rect 19682 30942 19684 30994
rect 17948 29426 18116 29428
rect 17948 29374 17950 29426
rect 18002 29374 18116 29426
rect 17948 29372 18116 29374
rect 19180 30322 19236 30334
rect 19180 30270 19182 30322
rect 19234 30270 19236 30322
rect 17948 29362 18004 29372
rect 19180 28532 19236 30270
rect 19628 29428 19684 30942
rect 20300 30994 20356 31836
rect 22316 31892 22372 31902
rect 22316 31798 22372 31836
rect 42924 31780 42980 31790
rect 42700 31778 42980 31780
rect 42700 31726 42926 31778
rect 42978 31726 42980 31778
rect 42700 31724 42980 31726
rect 21532 31668 21588 31678
rect 20300 30942 20302 30994
rect 20354 30942 20356 30994
rect 20300 30930 20356 30942
rect 21420 31612 21532 31668
rect 20300 30436 20356 30446
rect 20188 30100 20244 30110
rect 20188 30006 20244 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20300 29428 20356 30380
rect 21308 30100 21364 30110
rect 20412 30098 21364 30100
rect 20412 30046 21310 30098
rect 21362 30046 21364 30098
rect 20412 30044 21364 30046
rect 20412 29650 20468 30044
rect 21308 30034 21364 30044
rect 20412 29598 20414 29650
rect 20466 29598 20468 29650
rect 20412 29586 20468 29598
rect 20972 29652 21028 29662
rect 21420 29652 21476 31612
rect 21532 31602 21588 31612
rect 23548 31668 23604 31678
rect 23548 31574 23604 31612
rect 42700 31218 42756 31724
rect 42924 31714 42980 31724
rect 44044 31668 44100 31678
rect 44044 31574 44100 31612
rect 42700 31166 42702 31218
rect 42754 31166 42756 31218
rect 42700 31154 42756 31166
rect 22540 31106 22596 31118
rect 28028 31108 28084 31118
rect 22540 31054 22542 31106
rect 22594 31054 22596 31106
rect 22540 30436 22596 31054
rect 27916 31052 28028 31108
rect 27020 30884 27076 30894
rect 22540 30370 22596 30380
rect 23324 30770 23380 30782
rect 23324 30718 23326 30770
rect 23378 30718 23380 30770
rect 21756 30324 21812 30334
rect 20972 29650 21476 29652
rect 20972 29598 20974 29650
rect 21026 29598 21476 29650
rect 20972 29596 21476 29598
rect 21644 30098 21700 30110
rect 21644 30046 21646 30098
rect 21698 30046 21700 30098
rect 20972 29586 21028 29596
rect 21644 29540 21700 30046
rect 20300 29372 20692 29428
rect 19404 28644 19460 28654
rect 19628 28644 19684 29372
rect 20636 28754 20692 29372
rect 20636 28702 20638 28754
rect 20690 28702 20692 28754
rect 20636 28690 20692 28702
rect 21308 29426 21364 29438
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 19740 28644 19796 28654
rect 19404 28550 19460 28588
rect 19516 28642 19796 28644
rect 19516 28590 19742 28642
rect 19794 28590 19796 28642
rect 19516 28588 19796 28590
rect 19180 28466 19236 28476
rect 18844 27970 18900 27982
rect 18844 27918 18846 27970
rect 18898 27918 18900 27970
rect 17724 27748 17780 27758
rect 17724 27076 17780 27692
rect 18060 27748 18116 27758
rect 18060 27746 18676 27748
rect 18060 27694 18062 27746
rect 18114 27694 18676 27746
rect 18060 27692 18676 27694
rect 18060 27682 18116 27692
rect 17724 27010 17780 27020
rect 18620 26962 18676 27692
rect 18620 26910 18622 26962
rect 18674 26910 18676 26962
rect 18620 26898 18676 26910
rect 18844 26404 18900 27918
rect 19404 27188 19460 27198
rect 19404 27094 19460 27132
rect 18844 26338 18900 26348
rect 19068 26964 19124 26974
rect 19068 25394 19124 26908
rect 19180 26852 19236 26862
rect 19180 26180 19236 26796
rect 19516 26852 19572 28588
rect 19740 28578 19796 28588
rect 20524 28642 20580 28654
rect 20524 28590 20526 28642
rect 20578 28590 20580 28642
rect 20524 28420 20580 28590
rect 21308 28532 21364 29374
rect 20580 28364 20692 28420
rect 20524 28354 20580 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19852 27748 19908 27758
rect 19852 27746 20132 27748
rect 19852 27694 19854 27746
rect 19906 27694 20132 27746
rect 19852 27692 20132 27694
rect 19852 27682 19908 27692
rect 19852 27076 19908 27086
rect 19852 26982 19908 27020
rect 19628 26964 19684 26974
rect 19628 26870 19684 26908
rect 20076 26908 20132 27692
rect 20636 27076 20692 28364
rect 21308 27858 21364 28476
rect 21644 28420 21700 29484
rect 21756 29426 21812 30268
rect 23100 30324 23156 30334
rect 23100 30230 23156 30268
rect 23324 30100 23380 30718
rect 24668 30324 24724 30334
rect 23324 30034 23380 30044
rect 24108 30100 24164 30110
rect 24108 30006 24164 30044
rect 24220 29652 24276 29662
rect 24220 29558 24276 29596
rect 21756 29374 21758 29426
rect 21810 29374 21812 29426
rect 21756 29362 21812 29374
rect 22316 28756 22372 28766
rect 22316 28662 22372 28700
rect 23996 28642 24052 28654
rect 23996 28590 23998 28642
rect 24050 28590 24052 28642
rect 23548 28530 23604 28542
rect 23996 28532 24052 28590
rect 24668 28642 24724 30268
rect 25900 30324 25956 30334
rect 25900 30230 25956 30268
rect 24780 30100 24836 30110
rect 24780 29650 24836 30044
rect 26908 30100 26964 30110
rect 26908 30006 26964 30044
rect 24780 29598 24782 29650
rect 24834 29598 24836 29650
rect 24780 29586 24836 29598
rect 25340 29652 25396 29662
rect 25340 29558 25396 29596
rect 25228 29540 25284 29550
rect 25228 29446 25284 29484
rect 26236 29426 26292 29438
rect 26236 29374 26238 29426
rect 26290 29374 26292 29426
rect 24668 28590 24670 28642
rect 24722 28590 24724 28642
rect 24668 28578 24724 28590
rect 25788 29316 25844 29326
rect 23548 28478 23550 28530
rect 23602 28478 23604 28530
rect 21700 28364 22148 28420
rect 21644 28354 21700 28364
rect 21308 27806 21310 27858
rect 21362 27806 21364 27858
rect 21308 27794 21364 27806
rect 21756 27858 21812 27870
rect 21756 27806 21758 27858
rect 21810 27806 21812 27858
rect 20412 26962 20468 26974
rect 20412 26910 20414 26962
rect 20466 26910 20468 26962
rect 20076 26852 20244 26908
rect 19516 26786 19572 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26404 19684 26414
rect 19684 26348 19908 26404
rect 19628 26338 19684 26348
rect 19180 26114 19236 26124
rect 19628 26180 19684 26190
rect 19068 25342 19070 25394
rect 19122 25342 19124 25394
rect 19068 25330 19124 25342
rect 17948 25284 18004 25294
rect 17164 24162 17332 24164
rect 17164 24110 17166 24162
rect 17218 24110 17332 24162
rect 17164 24108 17332 24110
rect 17612 24498 17668 24510
rect 17612 24446 17614 24498
rect 17666 24446 17668 24498
rect 17164 24098 17220 24108
rect 16380 24052 16436 24062
rect 16380 23958 16436 23996
rect 17612 24052 17668 24446
rect 17612 23986 17668 23996
rect 17948 23826 18004 25228
rect 17948 23774 17950 23826
rect 18002 23774 18004 23826
rect 17948 23762 18004 23774
rect 18396 24722 18452 24734
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24500 18452 24670
rect 19628 24724 19684 26124
rect 19852 25730 19908 26348
rect 19852 25678 19854 25730
rect 19906 25678 19908 25730
rect 19852 25666 19908 25678
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 25060 20244 26852
rect 20300 25620 20356 25630
rect 20300 25526 20356 25564
rect 20412 25284 20468 26910
rect 20524 25620 20580 25630
rect 20636 25620 20692 27020
rect 20972 27746 21028 27758
rect 20972 27694 20974 27746
rect 21026 27694 21028 27746
rect 20972 26964 21028 27694
rect 21532 26964 21588 26974
rect 20972 26962 21588 26964
rect 20972 26910 21534 26962
rect 21586 26910 21588 26962
rect 20972 26908 21588 26910
rect 20524 25618 20692 25620
rect 20524 25566 20526 25618
rect 20578 25566 20692 25618
rect 20524 25564 20692 25566
rect 20524 25554 20580 25564
rect 20412 25218 20468 25228
rect 20188 25004 20468 25060
rect 19852 24724 19908 24734
rect 19684 24722 19908 24724
rect 19684 24670 19854 24722
rect 19906 24670 19908 24722
rect 19684 24668 19908 24670
rect 19628 24630 19684 24668
rect 16940 23716 16996 23726
rect 16828 23660 16940 23716
rect 16156 23326 16158 23378
rect 16210 23326 16212 23378
rect 16156 23314 16212 23326
rect 16380 23492 16436 23502
rect 15932 22418 15988 22428
rect 16380 21810 16436 23436
rect 16828 23044 16884 23660
rect 16940 23622 16996 23660
rect 18396 23716 18452 24444
rect 18396 23650 18452 23660
rect 19068 24610 19124 24622
rect 19068 24558 19070 24610
rect 19122 24558 19124 24610
rect 19068 23492 19124 24558
rect 19404 24612 19460 24622
rect 19404 24518 19460 24556
rect 19852 23716 19908 24668
rect 20300 24724 20356 24734
rect 20300 24630 20356 24668
rect 20188 23940 20244 23950
rect 20412 23940 20468 25004
rect 21532 24500 21588 26908
rect 21756 25620 21812 27806
rect 22092 27298 22148 28364
rect 22092 27246 22094 27298
rect 22146 27246 22148 27298
rect 22092 26852 22148 27246
rect 23436 27972 23492 27982
rect 23436 27186 23492 27916
rect 23436 27134 23438 27186
rect 23490 27134 23492 27186
rect 23436 27122 23492 27134
rect 23548 27188 23604 28478
rect 23548 27122 23604 27132
rect 23884 28476 23996 28532
rect 23884 27860 23940 28476
rect 23996 28466 24052 28476
rect 23996 27972 24052 27982
rect 23996 27878 24052 27916
rect 23884 27074 23940 27804
rect 25116 27860 25172 27870
rect 25116 27766 25172 27804
rect 25788 27858 25844 29260
rect 25788 27806 25790 27858
rect 25842 27806 25844 27858
rect 25788 27794 25844 27806
rect 26236 27860 26292 29374
rect 26908 29428 26964 29438
rect 27020 29428 27076 30828
rect 27804 30882 27860 30894
rect 27804 30830 27806 30882
rect 27858 30830 27860 30882
rect 27692 30100 27748 30110
rect 26908 29426 27076 29428
rect 26908 29374 26910 29426
rect 26962 29374 27076 29426
rect 26908 29372 27076 29374
rect 27132 30098 27748 30100
rect 27132 30046 27694 30098
rect 27746 30046 27748 30098
rect 27132 30044 27748 30046
rect 26908 29362 26964 29372
rect 27132 28418 27188 30044
rect 27692 30034 27748 30044
rect 27804 29316 27860 30830
rect 27804 29250 27860 29260
rect 27132 28366 27134 28418
rect 27186 28366 27188 28418
rect 27132 28354 27188 28366
rect 27356 28980 27412 28990
rect 26236 27794 26292 27804
rect 24780 27634 24836 27646
rect 24780 27582 24782 27634
rect 24834 27582 24836 27634
rect 23884 27022 23886 27074
rect 23938 27022 23940 27074
rect 23884 27010 23940 27022
rect 24332 27074 24388 27086
rect 24332 27022 24334 27074
rect 24386 27022 24388 27074
rect 23100 26962 23156 26974
rect 23100 26910 23102 26962
rect 23154 26910 23156 26962
rect 23100 26908 23156 26910
rect 23100 26852 23268 26908
rect 22092 26786 22148 26796
rect 21868 26292 21924 26302
rect 21868 26198 21924 26236
rect 23212 26290 23268 26796
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 23212 26226 23268 26238
rect 22988 26180 23044 26190
rect 21756 25554 21812 25564
rect 22764 26178 23044 26180
rect 22764 26126 22990 26178
rect 23042 26126 23044 26178
rect 22764 26124 23044 26126
rect 22764 24946 22820 26124
rect 22988 26114 23044 26124
rect 23772 26180 23828 26190
rect 22876 25620 22932 25630
rect 22876 25526 22932 25564
rect 22764 24894 22766 24946
rect 22818 24894 22820 24946
rect 22764 24882 22820 24894
rect 23324 25396 23380 25406
rect 23324 24946 23380 25340
rect 23324 24894 23326 24946
rect 23378 24894 23380 24946
rect 23324 24882 23380 24894
rect 23548 24612 23604 24622
rect 21532 24434 21588 24444
rect 23436 24610 23604 24612
rect 23436 24558 23550 24610
rect 23602 24558 23604 24610
rect 23436 24556 23604 24558
rect 23324 24052 23380 24062
rect 23324 23958 23380 23996
rect 20188 23938 20468 23940
rect 20188 23886 20190 23938
rect 20242 23886 20468 23938
rect 20188 23884 20468 23886
rect 20860 23940 20916 23950
rect 20188 23874 20244 23884
rect 20860 23846 20916 23884
rect 22316 23826 22372 23838
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 19852 23660 20356 23716
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19068 23426 19124 23436
rect 16940 23380 16996 23390
rect 16940 23286 16996 23324
rect 16828 22978 16884 22988
rect 18060 23266 18116 23278
rect 18060 23214 18062 23266
rect 18114 23214 18116 23266
rect 16940 22596 16996 22606
rect 16604 22260 16660 22270
rect 16604 22166 16660 22204
rect 16380 21758 16382 21810
rect 16434 21758 16436 21810
rect 16380 21746 16436 21758
rect 16940 21810 16996 22540
rect 17724 22484 17780 22494
rect 17388 22148 17444 22158
rect 17388 22146 17556 22148
rect 17388 22094 17390 22146
rect 17442 22094 17556 22146
rect 17388 22092 17556 22094
rect 17388 22082 17444 22092
rect 16940 21758 16942 21810
rect 16994 21758 16996 21810
rect 16940 21746 16996 21758
rect 15372 21522 15428 21532
rect 16380 20804 16436 20814
rect 15484 20802 16436 20804
rect 15484 20750 16382 20802
rect 16434 20750 16436 20802
rect 15484 20748 16436 20750
rect 14812 20018 14868 20030
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19236 14868 19966
rect 15036 19236 15092 19246
rect 14812 19234 15092 19236
rect 14812 19182 15038 19234
rect 15090 19182 15092 19234
rect 14812 19180 15092 19182
rect 15036 19012 15092 19180
rect 15036 18946 15092 18956
rect 14364 15934 14366 15986
rect 14418 15934 14420 15986
rect 14364 15922 14420 15934
rect 15372 16884 15428 16894
rect 15260 15876 15316 15886
rect 14700 15764 14756 15774
rect 14364 15204 14420 15214
rect 14364 14642 14420 15148
rect 14364 14590 14366 14642
rect 14418 14590 14420 14642
rect 14364 14578 14420 14590
rect 14700 14642 14756 15708
rect 14700 14590 14702 14642
rect 14754 14590 14756 14642
rect 14700 14578 14756 14590
rect 14812 15314 14868 15326
rect 14812 15262 14814 15314
rect 14866 15262 14868 15314
rect 14252 13582 14254 13634
rect 14306 13582 14308 13634
rect 14252 13570 14308 13582
rect 14812 13636 14868 15262
rect 15036 15204 15092 15214
rect 15036 14642 15092 15148
rect 15036 14590 15038 14642
rect 15090 14590 15092 14642
rect 15036 14578 15092 14590
rect 15260 13858 15316 15820
rect 15372 15314 15428 16828
rect 15484 16210 15540 20748
rect 16380 20738 16436 20748
rect 17052 20804 17108 20814
rect 17388 20804 17444 20814
rect 17052 20802 17444 20804
rect 17052 20750 17054 20802
rect 17106 20750 17390 20802
rect 17442 20750 17444 20802
rect 17052 20748 17444 20750
rect 17052 20738 17108 20748
rect 16156 20020 16212 20030
rect 17388 20020 17444 20748
rect 17500 20244 17556 22092
rect 17724 20802 17780 22428
rect 18060 21812 18116 23214
rect 19068 23156 19124 23166
rect 19068 23042 19124 23100
rect 19068 22990 19070 23042
rect 19122 22990 19124 23042
rect 19068 22978 19124 22990
rect 20300 23154 20356 23660
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 19740 22370 19796 22382
rect 19740 22318 19742 22370
rect 19794 22318 19796 22370
rect 19740 22260 19796 22318
rect 20300 22370 20356 23102
rect 20860 23156 20916 23166
rect 20860 23062 20916 23100
rect 20300 22318 20302 22370
rect 20354 22318 20356 22370
rect 20300 22306 20356 22318
rect 21420 22370 21476 22382
rect 21420 22318 21422 22370
rect 21474 22318 21476 22370
rect 19740 22194 19796 22204
rect 20860 22148 20916 22158
rect 20860 22054 20916 22092
rect 21420 22148 21476 22318
rect 21420 22082 21476 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 18060 21746 18116 21756
rect 21308 21810 21364 21822
rect 21308 21758 21310 21810
rect 21362 21758 21364 21810
rect 17724 20750 17726 20802
rect 17778 20750 17780 20802
rect 17724 20738 17780 20750
rect 18396 21586 18452 21598
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 17500 20178 17556 20188
rect 17500 20020 17556 20030
rect 17388 20018 17556 20020
rect 17388 19966 17502 20018
rect 17554 19966 17556 20018
rect 17388 19964 17556 19966
rect 16156 19926 16212 19964
rect 16828 19906 16884 19918
rect 16828 19854 16830 19906
rect 16882 19854 16884 19906
rect 15820 19794 15876 19806
rect 15820 19742 15822 19794
rect 15874 19742 15876 19794
rect 15820 19124 15876 19742
rect 15820 19058 15876 19068
rect 16716 19124 16772 19134
rect 15484 16158 15486 16210
rect 15538 16158 15540 16210
rect 15484 16146 15540 16158
rect 15596 18674 15652 18686
rect 15596 18622 15598 18674
rect 15650 18622 15652 18674
rect 15596 15426 15652 18622
rect 16492 18340 16548 18350
rect 16716 18340 16772 19068
rect 16828 19012 16884 19854
rect 16828 18946 16884 18956
rect 17052 18452 17108 18462
rect 17500 18452 17556 19964
rect 17948 20018 18004 20030
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17612 18452 17668 18462
rect 17500 18396 17612 18452
rect 16828 18340 16884 18350
rect 16716 18338 16884 18340
rect 16716 18286 16830 18338
rect 16882 18286 16884 18338
rect 16716 18284 16884 18286
rect 16492 18246 16548 18284
rect 16156 18228 16212 18238
rect 15596 15374 15598 15426
rect 15650 15374 15652 15426
rect 15596 15362 15652 15374
rect 16044 18226 16212 18228
rect 16044 18174 16158 18226
rect 16210 18174 16212 18226
rect 16044 18172 16212 18174
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 15372 15250 15428 15262
rect 15932 15204 15988 15242
rect 15932 15138 15988 15148
rect 15932 14420 15988 14430
rect 16044 14420 16100 18172
rect 16156 18162 16212 18172
rect 16492 17668 16548 17678
rect 16492 17666 16772 17668
rect 16492 17614 16494 17666
rect 16546 17614 16772 17666
rect 16492 17612 16772 17614
rect 16492 17602 16548 17612
rect 16380 17106 16436 17118
rect 16380 17054 16382 17106
rect 16434 17054 16436 17106
rect 16380 15540 16436 17054
rect 16716 16436 16772 17612
rect 16828 16772 16884 18284
rect 17052 17666 17108 18396
rect 17612 18358 17668 18396
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 17052 16884 17108 17614
rect 17948 17668 18004 19966
rect 18396 19122 18452 21534
rect 18844 21588 18900 21598
rect 18844 21494 18900 21532
rect 20300 20578 20356 20590
rect 20300 20526 20302 20578
rect 20354 20526 20356 20578
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20244 20020 20254
rect 19964 19346 20020 20188
rect 20188 20132 20244 20142
rect 20188 20038 20244 20076
rect 20300 19460 20356 20526
rect 20300 19394 20356 19404
rect 20860 20578 20916 20590
rect 20860 20526 20862 20578
rect 20914 20526 20916 20578
rect 19964 19294 19966 19346
rect 20018 19294 20020 19346
rect 19964 19282 20020 19294
rect 20300 19236 20356 19246
rect 20300 19142 20356 19180
rect 18396 19070 18398 19122
rect 18450 19070 18452 19122
rect 18060 18452 18116 18462
rect 18396 18452 18452 19070
rect 20748 19012 20804 19022
rect 20748 18918 20804 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18060 18450 18228 18452
rect 18060 18398 18062 18450
rect 18114 18398 18228 18450
rect 18060 18396 18228 18398
rect 18060 18386 18116 18396
rect 17948 17612 18116 17668
rect 17052 16818 17108 16828
rect 17164 17442 17220 17454
rect 17164 17390 17166 17442
rect 17218 17390 17220 17442
rect 16828 16706 16884 16716
rect 16940 16658 16996 16670
rect 16940 16606 16942 16658
rect 16994 16606 16996 16658
rect 16716 16380 16884 16436
rect 16380 15474 16436 15484
rect 16716 15874 16772 15886
rect 16716 15822 16718 15874
rect 16770 15822 16772 15874
rect 15932 14418 16100 14420
rect 15932 14366 15934 14418
rect 15986 14366 16100 14418
rect 15932 14364 16100 14366
rect 16604 14756 16660 14766
rect 15932 14354 15988 14364
rect 15260 13806 15262 13858
rect 15314 13806 15316 13858
rect 15260 13794 15316 13806
rect 14812 13580 15204 13636
rect 14252 12292 14308 12302
rect 14140 12290 14308 12292
rect 14140 12238 14254 12290
rect 14306 12238 14308 12290
rect 14140 12236 14308 12238
rect 14252 12226 14308 12236
rect 15148 12068 15204 13580
rect 15260 13076 15316 13086
rect 15260 12982 15316 13020
rect 16604 12850 16660 14700
rect 16716 14420 16772 15822
rect 16828 14642 16884 16380
rect 16828 14590 16830 14642
rect 16882 14590 16884 14642
rect 16828 14578 16884 14590
rect 16716 14354 16772 14364
rect 16604 12798 16606 12850
rect 16658 12798 16660 12850
rect 16604 12786 16660 12798
rect 16940 12292 16996 16606
rect 17164 12852 17220 17390
rect 17724 17442 17780 17454
rect 17724 17390 17726 17442
rect 17778 17390 17780 17442
rect 17500 16770 17556 16782
rect 17500 16718 17502 16770
rect 17554 16718 17556 16770
rect 17500 15986 17556 16718
rect 17724 16324 17780 17390
rect 18060 17108 18116 17612
rect 18060 17042 18116 17052
rect 17724 16258 17780 16268
rect 17836 16772 17892 16782
rect 17500 15934 17502 15986
rect 17554 15934 17556 15986
rect 17500 15922 17556 15934
rect 17724 15540 17780 15550
rect 17724 15426 17780 15484
rect 17724 15374 17726 15426
rect 17778 15374 17780 15426
rect 17724 15362 17780 15374
rect 17836 15204 17892 16716
rect 18060 16660 18116 16670
rect 17836 15138 17892 15148
rect 17948 16658 18116 16660
rect 17948 16606 18062 16658
rect 18114 16606 18116 16658
rect 17948 16604 18116 16606
rect 17948 14756 18004 16604
rect 18060 16594 18116 16604
rect 18172 15876 18228 18396
rect 18396 17444 18452 18396
rect 20524 18674 20580 18686
rect 20524 18622 20526 18674
rect 20578 18622 20580 18674
rect 20524 17780 20580 18622
rect 20860 18004 20916 20526
rect 20524 17714 20580 17724
rect 20748 17948 20916 18004
rect 20972 19794 21028 19806
rect 20972 19742 20974 19794
rect 21026 19742 21028 19794
rect 20188 17668 20244 17678
rect 20188 17666 20356 17668
rect 20188 17614 20190 17666
rect 20242 17614 20356 17666
rect 20188 17612 20356 17614
rect 20188 17602 20244 17612
rect 18396 17378 18452 17388
rect 20188 17444 20244 17454
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 18844 16994 18900 17006
rect 18844 16942 18846 16994
rect 18898 16942 18900 16994
rect 18844 16436 18900 16942
rect 18844 16370 18900 16380
rect 19516 16996 19572 17006
rect 18172 15810 18228 15820
rect 18844 16100 18900 16110
rect 18060 15204 18116 15242
rect 18844 15148 18900 16044
rect 18060 15138 18116 15148
rect 17948 14690 18004 14700
rect 18732 15092 18900 15148
rect 19068 15876 19124 15886
rect 18508 14420 18564 14430
rect 18508 14326 18564 14364
rect 17836 12852 17892 12862
rect 17164 12850 17892 12852
rect 17164 12798 17838 12850
rect 17890 12798 17892 12850
rect 17164 12796 17892 12798
rect 17836 12786 17892 12796
rect 17500 12292 17556 12302
rect 16940 12290 17556 12292
rect 16940 12238 17502 12290
rect 17554 12238 17556 12290
rect 16940 12236 17556 12238
rect 17500 12226 17556 12236
rect 15372 12068 15428 12078
rect 15148 12066 15428 12068
rect 15148 12014 15374 12066
rect 15426 12014 15428 12066
rect 15148 12012 15428 12014
rect 15372 12002 15428 12012
rect 18732 12066 18788 15092
rect 19068 13074 19124 15820
rect 19516 13636 19572 16940
rect 19740 16100 19796 16110
rect 19740 16006 19796 16044
rect 19852 15876 19908 17052
rect 20188 16098 20244 17388
rect 20188 16046 20190 16098
rect 20242 16046 20244 16098
rect 20188 16034 20244 16046
rect 19628 15820 19908 15876
rect 19628 15202 19684 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15150 19630 15202
rect 19682 15150 19684 15202
rect 19628 15138 19684 15150
rect 20300 15148 20356 17612
rect 20748 15426 20804 17948
rect 20860 17666 20916 17678
rect 20860 17614 20862 17666
rect 20914 17614 20916 17666
rect 20860 16884 20916 17614
rect 20972 17444 21028 19742
rect 21084 19794 21140 19806
rect 21084 19742 21086 19794
rect 21138 19742 21140 19794
rect 21084 18452 21140 19742
rect 21308 19346 21364 21758
rect 21980 21812 22036 21822
rect 21980 21718 22036 21756
rect 22092 21588 22148 21598
rect 21868 20914 21924 20926
rect 22092 20916 22148 21532
rect 22316 21026 22372 23774
rect 23436 23378 23492 24556
rect 23548 24546 23604 24556
rect 23436 23326 23438 23378
rect 23490 23326 23492 23378
rect 23436 23314 23492 23326
rect 23100 23044 23156 23054
rect 22652 22932 22708 22942
rect 22652 21698 22708 22876
rect 22652 21646 22654 21698
rect 22706 21646 22708 21698
rect 22652 21634 22708 21646
rect 22316 20974 22318 21026
rect 22370 20974 22372 21026
rect 22316 20962 22372 20974
rect 21868 20862 21870 20914
rect 21922 20862 21924 20914
rect 21868 20242 21924 20862
rect 21868 20190 21870 20242
rect 21922 20190 21924 20242
rect 21868 20178 21924 20190
rect 21980 20914 22148 20916
rect 21980 20862 22094 20914
rect 22146 20862 22148 20914
rect 21980 20860 22148 20862
rect 21308 19294 21310 19346
rect 21362 19294 21364 19346
rect 21308 19282 21364 19294
rect 21420 19460 21476 19470
rect 21980 19460 22036 20860
rect 22092 20850 22148 20860
rect 23100 20690 23156 22988
rect 23100 20638 23102 20690
rect 23154 20638 23156 20690
rect 23100 20626 23156 20638
rect 23212 22260 23268 22270
rect 21084 18386 21140 18396
rect 21420 18338 21476 19404
rect 21644 19404 22036 19460
rect 22092 20132 22148 20142
rect 21644 19346 21700 19404
rect 21644 19294 21646 19346
rect 21698 19294 21700 19346
rect 21644 19236 21700 19294
rect 22092 19346 22148 20076
rect 22092 19294 22094 19346
rect 22146 19294 22148 19346
rect 22092 19282 22148 19294
rect 21644 18562 21700 19180
rect 22428 19236 22484 19246
rect 22428 19142 22484 19180
rect 21644 18510 21646 18562
rect 21698 18510 21700 18562
rect 21644 18498 21700 18510
rect 22540 18452 22596 18462
rect 21420 18286 21422 18338
rect 21474 18286 21476 18338
rect 21420 18274 21476 18286
rect 22092 18338 22148 18350
rect 22092 18286 22094 18338
rect 22146 18286 22148 18338
rect 21084 18228 21140 18238
rect 21084 18134 21140 18172
rect 21420 17780 21476 17790
rect 21420 17686 21476 17724
rect 21644 17554 21700 17566
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 20972 17388 21588 17444
rect 20860 16818 20916 16828
rect 21196 16882 21252 16894
rect 21196 16830 21198 16882
rect 21250 16830 21252 16882
rect 20748 15374 20750 15426
rect 20802 15374 20804 15426
rect 20748 15362 20804 15374
rect 20972 16660 21028 16670
rect 19740 15092 20356 15148
rect 19740 14642 19796 15092
rect 19740 14590 19742 14642
rect 19794 14590 19796 14642
rect 19740 14578 19796 14590
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20972 13858 21028 16604
rect 21196 15988 21252 16830
rect 21196 15922 21252 15932
rect 21308 16884 21364 16894
rect 21308 15540 21364 16828
rect 21308 15314 21364 15484
rect 21308 15262 21310 15314
rect 21362 15262 21364 15314
rect 21308 15250 21364 15262
rect 21420 16324 21476 16334
rect 21420 14642 21476 16268
rect 21420 14590 21422 14642
rect 21474 14590 21476 14642
rect 21420 14578 21476 14590
rect 20972 13806 20974 13858
rect 21026 13806 21028 13858
rect 20972 13794 21028 13806
rect 21532 13860 21588 17388
rect 21644 15988 21700 17502
rect 22092 17444 22148 18286
rect 22316 17666 22372 17678
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 17444 22372 17614
rect 22092 17442 22372 17444
rect 22092 17390 22094 17442
rect 22146 17390 22372 17442
rect 22092 17388 22372 17390
rect 21756 16884 21812 16894
rect 22092 16884 22148 17388
rect 22540 16994 22596 18396
rect 23212 18338 23268 22204
rect 23548 22260 23604 22270
rect 23772 22260 23828 26124
rect 24332 25620 24388 27022
rect 24332 25554 24388 25564
rect 23884 25396 23940 25406
rect 23884 25302 23940 25340
rect 24780 25396 24836 27582
rect 27356 27298 27412 28924
rect 27692 28868 27748 28878
rect 27916 28868 27972 31052
rect 28028 31042 28084 31052
rect 28700 31106 28756 31118
rect 28700 31054 28702 31106
rect 28754 31054 28756 31106
rect 27692 28866 27972 28868
rect 27692 28814 27694 28866
rect 27746 28814 27972 28866
rect 27692 28812 27972 28814
rect 28028 30100 28084 30110
rect 27692 28802 27748 28812
rect 28028 28644 28084 30044
rect 28700 28980 28756 31054
rect 31500 31108 31556 31118
rect 31500 31014 31556 31052
rect 32732 31108 32788 31118
rect 30492 30884 30548 30894
rect 30492 30790 30548 30828
rect 31052 30322 31108 30334
rect 31052 30270 31054 30322
rect 31106 30270 31108 30322
rect 29484 30100 29540 30110
rect 29484 30006 29540 30044
rect 29372 29986 29428 29998
rect 29372 29934 29374 29986
rect 29426 29934 29428 29986
rect 29372 29650 29428 29934
rect 29372 29598 29374 29650
rect 29426 29598 29428 29650
rect 29372 29586 29428 29598
rect 29708 29316 29764 29326
rect 29596 29092 29652 29102
rect 28700 28914 28756 28924
rect 29484 29036 29596 29092
rect 27356 27246 27358 27298
rect 27410 27246 27412 27298
rect 27356 27234 27412 27246
rect 27916 28588 28084 28644
rect 29036 28642 29092 28654
rect 29036 28590 29038 28642
rect 29090 28590 29092 28642
rect 27916 28530 27972 28588
rect 27916 28478 27918 28530
rect 27970 28478 27972 28530
rect 26572 26964 26628 26974
rect 26572 26870 26628 26908
rect 27580 26964 27636 26974
rect 27580 26870 27636 26908
rect 27916 26964 27972 28478
rect 28028 28418 28084 28430
rect 28028 28366 28030 28418
rect 28082 28366 28084 28418
rect 28028 28082 28084 28366
rect 28028 28030 28030 28082
rect 28082 28030 28084 28082
rect 28028 28018 28084 28030
rect 27916 26870 27972 26908
rect 28588 27860 28644 27870
rect 28588 26402 28644 27804
rect 29036 27860 29092 28590
rect 29036 27766 29092 27804
rect 29484 27858 29540 29036
rect 29596 29026 29652 29036
rect 29708 28642 29764 29260
rect 29932 29204 29988 29214
rect 29932 29110 29988 29148
rect 31052 29092 31108 30270
rect 32060 30098 32116 30110
rect 32060 30046 32062 30098
rect 32114 30046 32116 30098
rect 31500 29316 31556 29326
rect 31052 29026 31108 29036
rect 31388 29314 31556 29316
rect 31388 29262 31502 29314
rect 31554 29262 31556 29314
rect 31388 29260 31556 29262
rect 29708 28590 29710 28642
rect 29762 28590 29764 28642
rect 29708 28578 29764 28590
rect 31164 28756 31220 28766
rect 29484 27806 29486 27858
rect 29538 27806 29540 27858
rect 29484 27794 29540 27806
rect 28588 26350 28590 26402
rect 28642 26350 28644 26402
rect 26796 26180 26852 26190
rect 26796 26086 26852 26124
rect 25676 25620 25732 25630
rect 25676 25526 25732 25564
rect 24780 25330 24836 25340
rect 26908 25396 26964 25406
rect 26908 25302 26964 25340
rect 27020 25172 27076 25182
rect 26460 24724 26516 24734
rect 23884 24612 23940 24622
rect 23884 24518 23940 24556
rect 24444 24612 24500 24622
rect 24332 24500 24388 24510
rect 24332 24050 24388 24444
rect 24332 23998 24334 24050
rect 24386 23998 24388 24050
rect 24332 23986 24388 23998
rect 24444 23156 24500 24556
rect 26236 24500 26292 24510
rect 25228 24052 25284 24062
rect 24556 23940 24612 23950
rect 24556 23846 24612 23884
rect 25228 23938 25284 23996
rect 25228 23886 25230 23938
rect 25282 23886 25284 23938
rect 25228 23874 25284 23886
rect 25788 23940 25844 23950
rect 24556 23156 24612 23166
rect 24444 23100 24556 23156
rect 24556 23062 24612 23100
rect 25452 23156 25508 23166
rect 24332 23044 24388 23054
rect 25452 23044 25508 23100
rect 24332 22950 24388 22988
rect 25340 23042 25508 23044
rect 25340 22990 25454 23042
rect 25506 22990 25508 23042
rect 25340 22988 25508 22990
rect 23996 22932 24052 22942
rect 23996 22838 24052 22876
rect 23548 22258 23828 22260
rect 23548 22206 23550 22258
rect 23602 22206 23828 22258
rect 23548 22204 23828 22206
rect 23548 19012 23604 22204
rect 25340 21588 25396 22988
rect 25452 22978 25508 22988
rect 25396 21532 25508 21588
rect 25340 21494 25396 21532
rect 23660 21474 23716 21486
rect 23660 21422 23662 21474
rect 23714 21422 23716 21474
rect 23660 20804 23716 21422
rect 23660 20738 23716 20748
rect 25340 20804 25396 20814
rect 25340 20710 25396 20748
rect 24108 20018 24164 20030
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 23548 18946 23604 18956
rect 23884 19234 23940 19246
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 23884 19012 23940 19182
rect 23884 18946 23940 18956
rect 23212 18286 23214 18338
rect 23266 18286 23268 18338
rect 23212 18274 23268 18286
rect 23548 18228 23604 18238
rect 22540 16942 22542 16994
rect 22594 16942 22596 16994
rect 22540 16930 22596 16942
rect 22988 17666 23044 17678
rect 22988 17614 22990 17666
rect 23042 17614 23044 17666
rect 21812 16828 22148 16884
rect 21756 16790 21812 16828
rect 22988 16772 23044 17614
rect 23436 16772 23492 16782
rect 22988 16770 23492 16772
rect 22988 16718 23438 16770
rect 23490 16718 23492 16770
rect 22988 16716 23492 16718
rect 23436 16706 23492 16716
rect 22092 16436 22148 16446
rect 21980 15988 22036 15998
rect 21644 15986 22036 15988
rect 21644 15934 21982 15986
rect 22034 15934 22036 15986
rect 21644 15932 22036 15934
rect 21756 15314 21812 15326
rect 21756 15262 21758 15314
rect 21810 15262 21812 15314
rect 21756 14868 21812 15262
rect 21980 15204 22036 15932
rect 22092 15874 22148 16380
rect 22764 16098 22820 16110
rect 22764 16046 22766 16098
rect 22818 16046 22820 16098
rect 22092 15822 22094 15874
rect 22146 15822 22148 15874
rect 22092 15810 22148 15822
rect 22316 15988 22372 15998
rect 21756 14812 21924 14868
rect 21644 14532 21700 14542
rect 21868 14532 21924 14812
rect 21644 14418 21700 14476
rect 21644 14366 21646 14418
rect 21698 14366 21700 14418
rect 21644 14354 21700 14366
rect 21756 14476 21924 14532
rect 21980 14532 22036 15148
rect 21644 13860 21700 13870
rect 21532 13858 21700 13860
rect 21532 13806 21646 13858
rect 21698 13806 21700 13858
rect 21532 13804 21700 13806
rect 21644 13794 21700 13804
rect 19740 13636 19796 13646
rect 19516 13634 19796 13636
rect 19516 13582 19742 13634
rect 19794 13582 19796 13634
rect 19516 13580 19796 13582
rect 19740 13570 19796 13580
rect 19068 13022 19070 13074
rect 19122 13022 19124 13074
rect 19068 13010 19124 13022
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 18732 12014 18734 12066
rect 18786 12014 18788 12066
rect 18732 12002 18788 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 21756 11508 21812 14476
rect 21980 14466 22036 14476
rect 22316 12066 22372 15932
rect 22764 15540 22820 16046
rect 22764 15474 22820 15484
rect 23324 16098 23380 16110
rect 23324 16046 23326 16098
rect 23378 16046 23380 16098
rect 23324 14084 23380 16046
rect 23436 15540 23492 15550
rect 23436 14530 23492 15484
rect 23436 14478 23438 14530
rect 23490 14478 23492 14530
rect 23436 14466 23492 14478
rect 23324 14018 23380 14028
rect 22988 13636 23044 13646
rect 22988 13542 23044 13580
rect 23324 13412 23380 13422
rect 23324 12850 23380 13356
rect 23324 12798 23326 12850
rect 23378 12798 23380 12850
rect 23324 12786 23380 12798
rect 22540 12740 22596 12750
rect 22540 12738 23044 12740
rect 22540 12686 22542 12738
rect 22594 12686 23044 12738
rect 22540 12684 23044 12686
rect 22540 12674 22596 12684
rect 22316 12014 22318 12066
rect 22370 12014 22372 12066
rect 22316 12002 22372 12014
rect 21756 11442 21812 11452
rect 22988 11282 23044 12684
rect 23548 12290 23604 18172
rect 23548 12238 23550 12290
rect 23602 12238 23604 12290
rect 23548 12226 23604 12238
rect 23884 14530 23940 14542
rect 23884 14478 23886 14530
rect 23938 14478 23940 14530
rect 23884 11508 23940 14478
rect 24108 13636 24164 19966
rect 24556 20018 24612 20030
rect 24556 19966 24558 20018
rect 24610 19966 24612 20018
rect 24332 19908 24388 19918
rect 24332 19234 24388 19852
rect 24332 19182 24334 19234
rect 24386 19182 24388 19234
rect 24332 19170 24388 19182
rect 24556 19012 24612 19966
rect 25452 20018 25508 21532
rect 25788 21586 25844 23884
rect 26236 23828 26292 24444
rect 26460 23940 26516 24668
rect 27020 24722 27076 25116
rect 27020 24670 27022 24722
rect 27074 24670 27076 24722
rect 27020 24658 27076 24670
rect 27132 24724 27188 24734
rect 26460 23874 26516 23884
rect 26236 23154 26292 23772
rect 26236 23102 26238 23154
rect 26290 23102 26292 23154
rect 26236 23090 26292 23102
rect 27132 23154 27188 24668
rect 28588 24724 28644 26350
rect 28812 27634 28868 27646
rect 28812 27582 28814 27634
rect 28866 27582 28868 27634
rect 28812 25396 28868 27582
rect 30492 27076 30548 27086
rect 30268 27074 30548 27076
rect 30268 27022 30494 27074
rect 30546 27022 30548 27074
rect 30268 27020 30548 27022
rect 29260 26964 29316 26974
rect 29260 26870 29316 26908
rect 28812 25330 28868 25340
rect 29372 26850 29428 26862
rect 29372 26798 29374 26850
rect 29426 26798 29428 26850
rect 29372 24946 29428 26798
rect 30156 25620 30212 25630
rect 29932 25618 30212 25620
rect 29932 25566 30158 25618
rect 30210 25566 30212 25618
rect 29932 25564 30212 25566
rect 29932 25060 29988 25564
rect 30156 25554 30212 25564
rect 30268 25396 30324 27020
rect 30492 27010 30548 27020
rect 31164 27074 31220 28700
rect 31164 27022 31166 27074
rect 31218 27022 31220 27074
rect 31164 27010 31220 27022
rect 30156 25340 30324 25396
rect 31388 26964 31444 29260
rect 31500 29250 31556 29260
rect 31836 29314 31892 29326
rect 31836 29262 31838 29314
rect 31890 29262 31892 29314
rect 31836 28532 31892 29262
rect 31948 28532 32004 28542
rect 31836 28530 32004 28532
rect 31836 28478 31950 28530
rect 32002 28478 32004 28530
rect 31836 28476 32004 28478
rect 31948 28466 32004 28476
rect 31836 27970 31892 27982
rect 31836 27918 31838 27970
rect 31890 27918 31892 27970
rect 31388 26068 31444 26908
rect 30156 25060 30212 25340
rect 29932 24994 29988 25004
rect 30044 25004 30212 25060
rect 29372 24894 29374 24946
rect 29426 24894 29428 24946
rect 29372 24882 29428 24894
rect 28588 24658 28644 24668
rect 29036 24724 29092 24734
rect 29036 23938 29092 24668
rect 29036 23886 29038 23938
rect 29090 23886 29092 23938
rect 29036 23874 29092 23886
rect 29708 23938 29764 23950
rect 29708 23886 29710 23938
rect 29762 23886 29764 23938
rect 27692 23716 27748 23726
rect 28252 23716 28308 23726
rect 27692 23714 28196 23716
rect 27692 23662 27694 23714
rect 27746 23662 28196 23714
rect 27692 23660 28196 23662
rect 27692 23650 27748 23660
rect 27132 23102 27134 23154
rect 27186 23102 27188 23154
rect 27132 23090 27188 23102
rect 27580 23154 27636 23166
rect 27580 23102 27582 23154
rect 27634 23102 27636 23154
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25564 21476 25620 21486
rect 25564 21474 25732 21476
rect 25564 21422 25566 21474
rect 25618 21422 25732 21474
rect 25564 21420 25732 21422
rect 25564 21410 25620 21420
rect 25676 20244 25732 21420
rect 25788 20802 25844 21534
rect 26460 21588 26516 21598
rect 26460 21494 26516 21532
rect 27580 20916 27636 23102
rect 27916 22484 27972 22494
rect 27916 22390 27972 22428
rect 28140 22482 28196 23660
rect 28252 23622 28308 23660
rect 28924 23044 28980 23054
rect 28476 22484 28532 22494
rect 28140 22430 28142 22482
rect 28194 22430 28196 22482
rect 28140 22418 28196 22430
rect 28364 22428 28476 22484
rect 27580 20850 27636 20860
rect 25788 20750 25790 20802
rect 25842 20750 25844 20802
rect 25788 20738 25844 20750
rect 27020 20804 27076 20814
rect 25676 20188 26628 20244
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 25452 19954 25508 19966
rect 26012 20018 26068 20030
rect 26460 20020 26516 20030
rect 26012 19966 26014 20018
rect 26066 19966 26068 20018
rect 24556 18946 24612 18956
rect 25228 19906 25284 19918
rect 25228 19854 25230 19906
rect 25282 19854 25284 19906
rect 24556 18788 24612 18798
rect 24556 18562 24612 18732
rect 24556 18510 24558 18562
rect 24610 18510 24612 18562
rect 24556 18498 24612 18510
rect 25228 17554 25284 19854
rect 26012 19012 26068 19966
rect 25228 17502 25230 17554
rect 25282 17502 25284 17554
rect 25228 17490 25284 17502
rect 25340 18340 25396 18350
rect 25116 16660 25172 16670
rect 25116 16566 25172 16604
rect 24220 15538 24276 15550
rect 24220 15486 24222 15538
rect 24274 15486 24276 15538
rect 24220 15428 24276 15486
rect 25340 15540 25396 18284
rect 26012 18340 26068 18956
rect 26012 18246 26068 18284
rect 26348 20018 26516 20020
rect 26348 19966 26462 20018
rect 26514 19966 26516 20018
rect 26348 19964 26516 19966
rect 26012 17892 26068 17902
rect 26012 17798 26068 17836
rect 25900 16994 25956 17006
rect 25900 16942 25902 16994
rect 25954 16942 25956 16994
rect 25900 16212 25956 16942
rect 26348 16996 26404 19964
rect 26460 19954 26516 19964
rect 26572 19122 26628 20188
rect 27020 20188 27076 20748
rect 28364 20802 28420 22428
rect 28476 22390 28532 22428
rect 28924 21810 28980 22988
rect 28924 21758 28926 21810
rect 28978 21758 28980 21810
rect 28924 21746 28980 21758
rect 29372 22932 29428 22942
rect 29372 22484 29428 22876
rect 29708 22596 29764 23886
rect 30044 23940 30100 25004
rect 31388 24834 31444 26012
rect 31500 27636 31556 27646
rect 31500 25394 31556 27580
rect 31500 25342 31502 25394
rect 31554 25342 31556 25394
rect 31500 25330 31556 25342
rect 31388 24782 31390 24834
rect 31442 24782 31444 24834
rect 31388 24770 31444 24782
rect 31724 24836 31780 24846
rect 31836 24836 31892 27918
rect 31724 24834 31892 24836
rect 31724 24782 31726 24834
rect 31778 24782 31892 24834
rect 31724 24780 31892 24782
rect 31724 24770 31780 24780
rect 31052 24724 31108 24734
rect 31052 24630 31108 24668
rect 31612 24724 31668 24734
rect 30156 24612 30212 24622
rect 30156 24518 30212 24556
rect 29932 23378 29988 23390
rect 29932 23326 29934 23378
rect 29986 23326 29988 23378
rect 29932 23268 29988 23326
rect 29932 23202 29988 23212
rect 29708 22530 29764 22540
rect 29820 22932 29876 22942
rect 29372 22370 29428 22428
rect 29372 22318 29374 22370
rect 29426 22318 29428 22370
rect 29372 20914 29428 22318
rect 29596 22258 29652 22270
rect 29596 22206 29598 22258
rect 29650 22206 29652 22258
rect 29484 21364 29540 21374
rect 29484 21270 29540 21308
rect 29372 20862 29374 20914
rect 29426 20862 29428 20914
rect 29372 20850 29428 20862
rect 28364 20750 28366 20802
rect 28418 20750 28420 20802
rect 28364 20738 28420 20750
rect 28364 20578 28420 20590
rect 28364 20526 28366 20578
rect 28418 20526 28420 20578
rect 28364 20188 28420 20526
rect 29596 20188 29652 22206
rect 29820 21810 29876 22876
rect 30044 22370 30100 23884
rect 31500 23268 31556 23278
rect 31500 23174 31556 23212
rect 31612 23156 31668 24668
rect 32060 24612 32116 30046
rect 32620 30100 32676 30110
rect 32620 28082 32676 30044
rect 32732 28866 32788 31052
rect 34636 31108 34692 31118
rect 34636 31014 34692 31052
rect 42476 31108 42532 31118
rect 42476 30994 42532 31052
rect 43820 31108 43876 31118
rect 43820 31014 43876 31052
rect 42476 30942 42478 30994
rect 42530 30942 42532 30994
rect 42476 30930 42532 30942
rect 43596 30996 43652 31006
rect 43596 30902 43652 30940
rect 44156 30996 44212 31006
rect 44156 30902 44212 30940
rect 35980 30882 36036 30894
rect 35980 30830 35982 30882
rect 36034 30830 36036 30882
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 33852 30322 33908 30334
rect 33852 30270 33854 30322
rect 33906 30270 33908 30322
rect 32732 28814 32734 28866
rect 32786 28814 32788 28866
rect 32732 28802 32788 28814
rect 33516 28868 33572 28878
rect 32620 28030 32622 28082
rect 32674 28030 32676 28082
rect 32620 28018 32676 28030
rect 33068 28642 33124 28654
rect 33068 28590 33070 28642
rect 33122 28590 33124 28642
rect 32956 27636 33012 27646
rect 32956 27542 33012 27580
rect 33068 26964 33124 28590
rect 33516 28642 33572 28812
rect 33852 28756 33908 30270
rect 34860 30100 34916 30110
rect 34860 30006 34916 30044
rect 35644 30098 35700 30110
rect 35644 30046 35646 30098
rect 35698 30046 35700 30098
rect 34188 29540 34244 29550
rect 34076 29316 34132 29326
rect 34076 29222 34132 29260
rect 33852 28690 33908 28700
rect 33516 28590 33518 28642
rect 33570 28590 33572 28642
rect 33516 28578 33572 28590
rect 33740 27972 33796 27982
rect 33740 27970 33908 27972
rect 33740 27918 33742 27970
rect 33794 27918 33908 27970
rect 33740 27916 33908 27918
rect 33740 27906 33796 27916
rect 33068 26898 33124 26908
rect 33404 26850 33460 26862
rect 33404 26798 33406 26850
rect 33458 26798 33460 26850
rect 33404 26514 33460 26798
rect 33404 26462 33406 26514
rect 33458 26462 33460 26514
rect 33404 26450 33460 26462
rect 32172 26290 32228 26302
rect 32172 26238 32174 26290
rect 32226 26238 32228 26290
rect 32172 26180 32228 26238
rect 33404 26292 33460 26302
rect 33404 26198 33460 26236
rect 32172 25284 32228 26124
rect 32956 25618 33012 25630
rect 32956 25566 32958 25618
rect 33010 25566 33012 25618
rect 32732 25284 32788 25294
rect 32172 25190 32228 25228
rect 32284 25282 32788 25284
rect 32284 25230 32734 25282
rect 32786 25230 32788 25282
rect 32284 25228 32788 25230
rect 32284 24724 32340 25228
rect 32732 25218 32788 25228
rect 32956 25172 33012 25566
rect 32956 25106 33012 25116
rect 33628 25284 33684 25294
rect 32284 24630 32340 24668
rect 33516 25060 33572 25070
rect 32060 24546 32116 24556
rect 32508 24610 32564 24622
rect 32508 24558 32510 24610
rect 32562 24558 32564 24610
rect 31948 23716 32004 23726
rect 31724 23156 31780 23166
rect 31612 23154 31780 23156
rect 31612 23102 31726 23154
rect 31778 23102 31780 23154
rect 31612 23100 31780 23102
rect 30828 23044 30884 23054
rect 30828 22950 30884 22988
rect 31164 23044 31220 23054
rect 31164 22950 31220 22988
rect 31612 23044 31668 23100
rect 31724 23090 31780 23100
rect 31612 22978 31668 22988
rect 30604 22930 30660 22942
rect 30604 22878 30606 22930
rect 30658 22878 30660 22930
rect 30044 22318 30046 22370
rect 30098 22318 30100 22370
rect 30044 22306 30100 22318
rect 30492 22372 30548 22382
rect 30492 22278 30548 22316
rect 29820 21758 29822 21810
rect 29874 21758 29876 21810
rect 29820 21746 29876 21758
rect 30156 20916 30212 20926
rect 30156 20822 30212 20860
rect 30604 20692 30660 22878
rect 31948 21698 32004 23660
rect 32172 23714 32228 23726
rect 32172 23662 32174 23714
rect 32226 23662 32228 23714
rect 32172 23266 32228 23662
rect 32508 23380 32564 24558
rect 32844 23940 32900 23950
rect 32844 23846 32900 23884
rect 33516 23938 33572 25004
rect 33628 24722 33684 25228
rect 33852 25284 33908 27916
rect 34188 27298 34244 29484
rect 35308 29538 35364 29550
rect 35308 29486 35310 29538
rect 35362 29486 35364 29538
rect 35308 29204 35364 29486
rect 35308 29138 35364 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34188 27246 34190 27298
rect 34242 27246 34244 27298
rect 34188 27234 34244 27246
rect 35532 27186 35588 27198
rect 35532 27134 35534 27186
rect 35586 27134 35588 27186
rect 34860 27074 34916 27086
rect 34860 27022 34862 27074
rect 34914 27022 34916 27074
rect 34076 26964 34132 26974
rect 34076 26290 34132 26908
rect 34860 26964 34916 27022
rect 34076 26238 34078 26290
rect 34130 26238 34132 26290
rect 33964 25396 34020 25406
rect 33964 25302 34020 25340
rect 33852 25218 33908 25228
rect 33628 24670 33630 24722
rect 33682 24670 33684 24722
rect 33628 24658 33684 24670
rect 33516 23886 33518 23938
rect 33570 23886 33572 23938
rect 33516 23874 33572 23886
rect 34076 23940 34132 26238
rect 34524 26852 34580 26862
rect 34524 26290 34580 26796
rect 34524 26238 34526 26290
rect 34578 26238 34580 26290
rect 34524 26226 34580 26238
rect 34076 23874 34132 23884
rect 34860 25506 34916 26908
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34860 25454 34862 25506
rect 34914 25454 34916 25506
rect 32508 23314 32564 23324
rect 32732 23714 32788 23726
rect 32732 23662 32734 23714
rect 32786 23662 32788 23714
rect 32172 23214 32174 23266
rect 32226 23214 32228 23266
rect 32172 23202 32228 23214
rect 31948 21646 31950 21698
rect 32002 21646 32004 21698
rect 31948 21634 32004 21646
rect 32508 23044 32564 23054
rect 32508 21588 32564 22988
rect 32732 22260 32788 23662
rect 32956 23492 33012 23502
rect 32956 23378 33012 23436
rect 32956 23326 32958 23378
rect 33010 23326 33012 23378
rect 32956 23314 33012 23326
rect 33516 23380 33572 23390
rect 33516 23286 33572 23324
rect 32732 22194 32788 22204
rect 33180 22596 33236 22606
rect 32956 22148 33012 22158
rect 32956 22146 33124 22148
rect 32956 22094 32958 22146
rect 33010 22094 33124 22146
rect 32956 22092 33124 22094
rect 32956 22082 33012 22092
rect 33068 21698 33124 22092
rect 33068 21646 33070 21698
rect 33122 21646 33124 21698
rect 33068 21634 33124 21646
rect 32508 21522 32564 21532
rect 30716 21476 30772 21486
rect 30716 21382 30772 21420
rect 30604 20626 30660 20636
rect 31164 21364 31220 21374
rect 31164 20690 31220 21308
rect 33180 20914 33236 22540
rect 33516 22596 33572 22606
rect 33516 22502 33572 22540
rect 34748 22484 34804 22494
rect 34748 22390 34804 22428
rect 34860 22260 34916 25454
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 24052 35588 27134
rect 35644 26292 35700 30046
rect 35756 29986 35812 29998
rect 35756 29934 35758 29986
rect 35810 29934 35812 29986
rect 35756 28530 35812 29934
rect 35756 28478 35758 28530
rect 35810 28478 35812 28530
rect 35756 28466 35812 28478
rect 35980 27858 36036 30830
rect 37996 30322 38052 30334
rect 37996 30270 37998 30322
rect 38050 30270 38052 30322
rect 36540 30100 36596 30110
rect 36540 28866 36596 30044
rect 37884 29540 37940 29550
rect 37884 29446 37940 29484
rect 36540 28814 36542 28866
rect 36594 28814 36596 28866
rect 36540 28802 36596 28814
rect 36876 29314 36932 29326
rect 36876 29262 36878 29314
rect 36930 29262 36932 29314
rect 36876 28868 36932 29262
rect 36876 28802 36932 28812
rect 37548 28756 37604 28766
rect 36988 28642 37044 28654
rect 36988 28590 36990 28642
rect 37042 28590 37044 28642
rect 35980 27806 35982 27858
rect 36034 27806 36036 27858
rect 35980 27794 36036 27806
rect 36652 27860 36708 27870
rect 36988 27860 37044 28590
rect 37548 28642 37604 28700
rect 37548 28590 37550 28642
rect 37602 28590 37604 28642
rect 37548 28578 37604 28590
rect 36652 27858 37156 27860
rect 36652 27806 36654 27858
rect 36706 27806 36990 27858
rect 37042 27806 37156 27858
rect 36652 27804 37156 27806
rect 36652 27794 36708 27804
rect 36988 27794 37044 27804
rect 37100 27074 37156 27804
rect 37100 27022 37102 27074
rect 37154 27022 37156 27074
rect 36316 26964 36372 26974
rect 36372 26908 36484 26964
rect 36316 26870 36372 26908
rect 35644 25620 35700 26236
rect 35644 25526 35700 25564
rect 36428 25618 36484 26908
rect 36428 25566 36430 25618
rect 36482 25566 36484 25618
rect 36428 25554 36484 25566
rect 36876 26514 36932 26526
rect 36876 26462 36878 26514
rect 36930 26462 36932 26514
rect 35532 23986 35588 23996
rect 35644 24610 35700 24622
rect 35644 24558 35646 24610
rect 35698 24558 35700 24610
rect 35644 23940 35700 24558
rect 36876 24052 36932 26462
rect 36988 25620 37044 25630
rect 36988 25526 37044 25564
rect 37100 25508 37156 27022
rect 37436 27858 37492 27870
rect 37436 27806 37438 27858
rect 37490 27806 37492 27858
rect 37436 26180 37492 27806
rect 37548 27748 37604 27758
rect 37548 27074 37604 27692
rect 37548 27022 37550 27074
rect 37602 27022 37604 27074
rect 37548 27010 37604 27022
rect 37996 26852 38052 30270
rect 39004 30100 39060 30110
rect 39004 30006 39060 30044
rect 41804 28756 41860 28766
rect 41804 28662 41860 28700
rect 40796 28532 40852 28542
rect 40684 28476 40796 28532
rect 40012 28420 40068 28430
rect 40012 28418 40180 28420
rect 40012 28366 40014 28418
rect 40066 28366 40180 28418
rect 40012 28364 40180 28366
rect 40012 28354 40068 28364
rect 39676 27972 39732 27982
rect 39340 27970 39732 27972
rect 39340 27918 39678 27970
rect 39730 27918 39732 27970
rect 39340 27916 39732 27918
rect 37996 26786 38052 26796
rect 38220 27188 38276 27198
rect 37548 26404 37604 26414
rect 37548 26310 37604 26348
rect 37436 26114 37492 26124
rect 37548 25508 37604 25518
rect 37100 25506 37604 25508
rect 37100 25454 37550 25506
rect 37602 25454 37604 25506
rect 37100 25452 37604 25454
rect 37100 25284 37156 25294
rect 37100 25190 37156 25228
rect 37436 24612 37492 24622
rect 36988 24052 37044 24062
rect 36876 24050 37044 24052
rect 36876 23998 36990 24050
rect 37042 23998 37044 24050
rect 36876 23996 37044 23998
rect 36988 23986 37044 23996
rect 37212 24052 37268 24062
rect 35644 23874 35700 23884
rect 36428 23940 36484 23950
rect 35980 23714 36036 23726
rect 35980 23662 35982 23714
rect 36034 23662 36036 23714
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34748 22204 34916 22260
rect 35756 22260 35812 22270
rect 33852 22146 33908 22158
rect 33852 22094 33854 22146
rect 33906 22094 33908 22146
rect 33404 21588 33460 21598
rect 33404 21494 33460 21532
rect 33852 21588 33908 22094
rect 34300 22146 34356 22158
rect 34300 22094 34302 22146
rect 34354 22094 34356 22146
rect 33852 21494 33908 21532
rect 34188 21586 34244 21598
rect 34188 21534 34190 21586
rect 34242 21534 34244 21586
rect 33180 20862 33182 20914
rect 33234 20862 33236 20914
rect 33180 20850 33236 20862
rect 31164 20638 31166 20690
rect 31218 20638 31220 20690
rect 31164 20626 31220 20638
rect 33628 20804 33684 20814
rect 27020 20132 27300 20188
rect 28364 20132 28868 20188
rect 29596 20132 29764 20188
rect 26572 19070 26574 19122
rect 26626 19070 26628 19122
rect 26572 19058 26628 19070
rect 26460 18900 26516 18910
rect 26460 18452 26516 18844
rect 26460 18358 26516 18396
rect 27244 17668 27300 20132
rect 28812 20130 28868 20132
rect 28812 20078 28814 20130
rect 28866 20078 28868 20130
rect 28812 20066 28868 20078
rect 29596 19796 29652 19806
rect 29596 19702 29652 19740
rect 28252 19124 28308 19134
rect 28140 19122 28308 19124
rect 28140 19070 28254 19122
rect 28306 19070 28308 19122
rect 28140 19068 28308 19070
rect 27356 19010 27412 19022
rect 27356 18958 27358 19010
rect 27410 18958 27412 19010
rect 27356 18004 27412 18958
rect 27692 19012 27748 19022
rect 27692 18918 27748 18956
rect 27356 17938 27412 17948
rect 27356 17668 27412 17678
rect 27020 17666 27412 17668
rect 27020 17614 27358 17666
rect 27410 17614 27412 17666
rect 27020 17612 27412 17614
rect 26348 16930 26404 16940
rect 26572 17554 26628 17566
rect 26572 17502 26574 17554
rect 26626 17502 26628 17554
rect 25900 16146 25956 16156
rect 25788 15876 25844 15886
rect 26348 15876 26404 15886
rect 25788 15874 26292 15876
rect 25788 15822 25790 15874
rect 25842 15822 26292 15874
rect 25788 15820 26292 15822
rect 25788 15810 25844 15820
rect 25340 15446 25396 15484
rect 24220 15362 24276 15372
rect 25788 15428 25844 15438
rect 25788 15334 25844 15372
rect 26124 15428 26180 15438
rect 26236 15428 26292 15820
rect 26348 15782 26404 15820
rect 26460 15428 26516 15438
rect 26236 15426 26516 15428
rect 26236 15374 26462 15426
rect 26514 15374 26516 15426
rect 26236 15372 26516 15374
rect 26124 15334 26180 15372
rect 26460 15362 26516 15372
rect 26348 15204 26404 15214
rect 24108 13570 24164 13580
rect 24780 15090 24836 15102
rect 24780 15038 24782 15090
rect 24834 15038 24836 15090
rect 24780 13636 24836 15038
rect 26348 14306 26404 15148
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 14242 26404 14254
rect 24780 13570 24836 13580
rect 26124 14084 26180 14094
rect 25676 12962 25732 12974
rect 25676 12910 25678 12962
rect 25730 12910 25732 12962
rect 25676 12068 25732 12910
rect 26124 12068 26180 14028
rect 26572 13412 26628 17502
rect 26908 17554 26964 17566
rect 26908 17502 26910 17554
rect 26962 17502 26964 17554
rect 26908 16436 26964 17502
rect 26684 16380 26964 16436
rect 26684 15988 26740 16380
rect 26908 16212 26964 16222
rect 27020 16212 27076 17612
rect 27356 17602 27412 17612
rect 28140 17554 28196 19068
rect 28252 19058 28308 19068
rect 28140 17502 28142 17554
rect 28194 17502 28196 17554
rect 26908 16210 27076 16212
rect 26908 16158 26910 16210
rect 26962 16158 27076 16210
rect 26908 16156 27076 16158
rect 27804 16212 27860 16222
rect 26908 16146 26964 16156
rect 27804 16118 27860 16156
rect 26684 15428 26740 15932
rect 27468 15988 27524 15998
rect 27468 15894 27524 15932
rect 28140 15988 28196 17502
rect 28364 19010 28420 19022
rect 28364 18958 28366 19010
rect 28418 18958 28420 19010
rect 28364 17556 28420 18958
rect 28364 17490 28420 17500
rect 28588 19012 28644 19022
rect 28364 16996 28420 17006
rect 28252 16884 28308 16894
rect 28252 16790 28308 16828
rect 28140 15894 28196 15932
rect 27356 15874 27412 15886
rect 27356 15822 27358 15874
rect 27410 15822 27412 15874
rect 26684 15314 26740 15372
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15250 26740 15262
rect 27132 15540 27188 15550
rect 27132 15314 27188 15484
rect 27132 15262 27134 15314
rect 27186 15262 27188 15314
rect 27132 14644 27188 15262
rect 27356 15204 27412 15822
rect 27356 15138 27412 15148
rect 27804 15314 27860 15326
rect 27804 15262 27806 15314
rect 27858 15262 27860 15314
rect 27244 14644 27300 14654
rect 27580 14644 27636 14654
rect 27692 14644 27748 14654
rect 26572 13346 26628 13356
rect 26684 14642 27748 14644
rect 26684 14590 27246 14642
rect 27298 14590 27582 14642
rect 27634 14590 27694 14642
rect 27746 14590 27748 14642
rect 26684 14588 27748 14590
rect 26684 13076 26740 14588
rect 27244 14578 27300 14588
rect 27580 14550 27636 14588
rect 27692 14578 27748 14588
rect 26236 13074 26740 13076
rect 26236 13022 26686 13074
rect 26738 13022 26740 13074
rect 26236 13020 26740 13022
rect 26236 12962 26292 13020
rect 26684 13010 26740 13020
rect 26908 14306 26964 14318
rect 26908 14254 26910 14306
rect 26962 14254 26964 14306
rect 26236 12910 26238 12962
rect 26290 12910 26292 12962
rect 26236 12898 26292 12910
rect 26908 12852 26964 14254
rect 26908 12786 26964 12796
rect 27244 13636 27300 13646
rect 27244 12290 27300 13580
rect 27244 12238 27246 12290
rect 27298 12238 27300 12290
rect 27244 12226 27300 12238
rect 26236 12068 26292 12078
rect 26124 12066 26292 12068
rect 26124 12014 26238 12066
rect 26290 12014 26292 12066
rect 26124 12012 26292 12014
rect 25676 12002 25732 12012
rect 26236 12002 26292 12012
rect 24108 11508 24164 11518
rect 23884 11506 24164 11508
rect 23884 11454 24110 11506
rect 24162 11454 24164 11506
rect 23884 11452 24164 11454
rect 24108 11442 24164 11452
rect 26684 11508 26740 11518
rect 26684 11414 26740 11452
rect 27804 11508 27860 15262
rect 28140 14754 28196 14766
rect 28140 14702 28142 14754
rect 28194 14702 28196 14754
rect 28140 14642 28196 14702
rect 28140 14590 28142 14642
rect 28194 14590 28196 14642
rect 28140 14578 28196 14590
rect 28364 13634 28420 16940
rect 28588 16884 28644 18956
rect 29036 19010 29092 19022
rect 29036 18958 29038 19010
rect 29090 18958 29092 19010
rect 29036 18788 29092 18958
rect 29708 19010 29764 20132
rect 31948 20130 32004 20142
rect 31948 20078 31950 20130
rect 32002 20078 32004 20130
rect 29708 18958 29710 19010
rect 29762 18958 29764 19010
rect 29708 18946 29764 18958
rect 30044 19908 30100 19918
rect 30492 19908 30548 19918
rect 30044 19906 30548 19908
rect 30044 19854 30046 19906
rect 30098 19854 30494 19906
rect 30546 19854 30548 19906
rect 30044 19852 30548 19854
rect 30044 19012 30100 19852
rect 30492 19842 30548 19852
rect 30828 19908 30884 19918
rect 30828 19814 30884 19852
rect 29036 18722 29092 18732
rect 30044 18562 30100 18956
rect 30044 18510 30046 18562
rect 30098 18510 30100 18562
rect 30044 18498 30100 18510
rect 29148 18004 29204 18014
rect 29204 17948 29316 18004
rect 29148 17938 29204 17948
rect 29036 17444 29092 17454
rect 29036 17442 29204 17444
rect 29036 17390 29038 17442
rect 29090 17390 29204 17442
rect 29036 17388 29204 17390
rect 29036 17378 29092 17388
rect 28924 16884 28980 16894
rect 28588 16882 29092 16884
rect 28588 16830 28590 16882
rect 28642 16830 28926 16882
rect 28978 16830 29092 16882
rect 28588 16828 29092 16830
rect 28588 16210 28644 16828
rect 28924 16818 28980 16828
rect 28588 16158 28590 16210
rect 28642 16158 28644 16210
rect 28588 16146 28644 16158
rect 29036 16772 29092 16828
rect 29036 16098 29092 16716
rect 29036 16046 29038 16098
rect 29090 16046 29092 16098
rect 29036 16034 29092 16046
rect 29148 15652 29204 17388
rect 29148 15586 29204 15596
rect 28588 14754 28644 14766
rect 28588 14702 28590 14754
rect 28642 14702 28644 14754
rect 28588 14642 28644 14702
rect 28588 14590 28590 14642
rect 28642 14590 28644 14642
rect 28588 14578 28644 14590
rect 29260 13858 29316 17948
rect 31948 17892 32004 20078
rect 33516 20020 33572 20030
rect 33516 19926 33572 19964
rect 32172 19908 32228 19918
rect 32172 19234 32228 19852
rect 32172 19182 32174 19234
rect 32226 19182 32228 19234
rect 32172 19170 32228 19182
rect 32732 19236 32788 19246
rect 32732 19142 32788 19180
rect 33628 19122 33684 20748
rect 33964 20692 34020 20702
rect 33964 20598 34020 20636
rect 33628 19070 33630 19122
rect 33682 19070 33684 19122
rect 33628 19058 33684 19070
rect 33964 20018 34020 20030
rect 33964 19966 33966 20018
rect 34018 19966 34020 20018
rect 33964 19124 34020 19966
rect 34188 20020 34244 21534
rect 34300 21588 34356 22094
rect 34300 21522 34356 21532
rect 34748 20916 34804 22204
rect 35756 22166 35812 22204
rect 35980 22148 36036 23662
rect 36092 23154 36148 23166
rect 36092 23102 36094 23154
rect 36146 23102 36148 23154
rect 36092 23044 36148 23102
rect 36428 23156 36484 23884
rect 37212 23938 37268 23996
rect 37212 23886 37214 23938
rect 37266 23886 37268 23938
rect 37212 23874 37268 23886
rect 36540 23716 36596 23726
rect 36540 23622 36596 23660
rect 36764 23156 36820 23166
rect 36428 23154 36932 23156
rect 36428 23102 36430 23154
rect 36482 23102 36766 23154
rect 36818 23102 36932 23154
rect 36428 23100 36932 23102
rect 36428 23090 36484 23100
rect 36764 23090 36820 23100
rect 36092 22978 36148 22988
rect 36876 22370 36932 23100
rect 37436 23154 37492 24556
rect 37548 23940 37604 25452
rect 38220 25506 38276 27132
rect 38892 26178 38948 26190
rect 38892 26126 38894 26178
rect 38946 26126 38948 26178
rect 38220 25454 38222 25506
rect 38274 25454 38276 25506
rect 38220 25442 38276 25454
rect 38780 25620 38836 25630
rect 38444 24052 38500 24062
rect 37548 23874 37604 23884
rect 38108 23940 38164 23950
rect 38108 23846 38164 23884
rect 37436 23102 37438 23154
rect 37490 23102 37492 23154
rect 37436 23090 37492 23102
rect 36876 22318 36878 22370
rect 36930 22318 36932 22370
rect 36876 22306 36932 22318
rect 37548 22370 37604 22382
rect 37548 22318 37550 22370
rect 37602 22318 37604 22370
rect 35980 22082 36036 22092
rect 36988 22148 37044 22158
rect 34860 21812 34916 21822
rect 34860 21586 34916 21756
rect 34860 21534 34862 21586
rect 34914 21534 34916 21586
rect 34860 21522 34916 21534
rect 35756 21588 35812 21598
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35756 21026 35812 21532
rect 35756 20974 35758 21026
rect 35810 20974 35812 21026
rect 35756 20962 35812 20974
rect 34748 20802 34804 20860
rect 36428 20916 36484 20926
rect 36428 20822 36484 20860
rect 36988 20914 37044 22092
rect 37324 21812 37380 21822
rect 37324 21810 37492 21812
rect 37324 21758 37326 21810
rect 37378 21758 37492 21810
rect 37324 21756 37492 21758
rect 37324 21746 37380 21756
rect 37212 21700 37268 21710
rect 37212 21588 37268 21644
rect 37212 21532 37380 21588
rect 36988 20862 36990 20914
rect 37042 20862 37044 20914
rect 36988 20850 37044 20862
rect 37212 20916 37268 20926
rect 34748 20750 34750 20802
rect 34802 20750 34804 20802
rect 34748 20738 34804 20750
rect 34188 19236 34244 19964
rect 36204 20130 36260 20142
rect 36204 20078 36206 20130
rect 36258 20078 36260 20130
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35980 19572 36036 19582
rect 34188 19170 34244 19180
rect 35980 19234 36036 19516
rect 35980 19182 35982 19234
rect 36034 19182 36036 19234
rect 35980 19170 36036 19182
rect 33964 19058 34020 19068
rect 32844 19012 32900 19022
rect 32844 18918 32900 18956
rect 35644 19012 35700 19022
rect 36092 19012 36148 19022
rect 35700 18956 35812 19012
rect 35644 18946 35700 18956
rect 32060 18452 32116 18462
rect 32060 18358 32116 18396
rect 32508 18452 32564 18462
rect 33068 18452 33124 18462
rect 32564 18450 33124 18452
rect 32564 18398 33070 18450
rect 33122 18398 33124 18450
rect 32564 18396 33124 18398
rect 32508 18358 32564 18396
rect 33068 18386 33124 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 31948 17826 32004 17836
rect 32172 17666 32228 17678
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 29596 17556 29652 17566
rect 29596 17442 29652 17500
rect 29596 17390 29598 17442
rect 29650 17390 29652 17442
rect 29596 17378 29652 17390
rect 32172 17108 32228 17614
rect 32172 17042 32228 17052
rect 32508 17666 32564 17678
rect 32508 17614 32510 17666
rect 32562 17614 32564 17666
rect 31836 16994 31892 17006
rect 31836 16942 31838 16994
rect 31890 16942 31892 16994
rect 29596 16882 29652 16894
rect 29596 16830 29598 16882
rect 29650 16830 29652 16882
rect 29596 16324 29652 16830
rect 29596 16258 29652 16268
rect 30044 16884 30100 16894
rect 29708 16098 29764 16110
rect 29708 16046 29710 16098
rect 29762 16046 29764 16098
rect 29708 14644 29764 16046
rect 29708 14578 29764 14588
rect 29260 13806 29262 13858
rect 29314 13806 29316 13858
rect 29260 13794 29316 13806
rect 29372 14306 29428 14318
rect 29372 14254 29374 14306
rect 29426 14254 29428 14306
rect 28364 13582 28366 13634
rect 28418 13582 28420 13634
rect 28364 13570 28420 13582
rect 27804 11442 27860 11452
rect 28028 12740 28084 12750
rect 22988 11230 22990 11282
rect 23042 11230 23044 11282
rect 22988 11218 23044 11230
rect 28028 11282 28084 12684
rect 29372 12740 29428 14254
rect 30044 13076 30100 16828
rect 30940 16324 30996 16334
rect 30268 15876 30324 15886
rect 30324 15820 30436 15876
rect 30268 15810 30324 15820
rect 30268 15538 30324 15550
rect 30268 15486 30270 15538
rect 30322 15486 30324 15538
rect 30268 15428 30324 15486
rect 30268 15362 30324 15372
rect 30156 15204 30212 15214
rect 30156 14418 30212 15148
rect 30156 14366 30158 14418
rect 30210 14366 30212 14418
rect 30156 14354 30212 14366
rect 30156 13076 30212 13086
rect 30044 13074 30212 13076
rect 30044 13022 30158 13074
rect 30210 13022 30212 13074
rect 30044 13020 30212 13022
rect 30156 13010 30212 13020
rect 29372 12674 29428 12684
rect 30380 12290 30436 15820
rect 30828 15090 30884 15102
rect 30828 15038 30830 15090
rect 30882 15038 30884 15090
rect 30828 14532 30884 15038
rect 30828 14466 30884 14476
rect 30940 13634 30996 16268
rect 31388 15988 31444 15998
rect 31052 15428 31108 15438
rect 31052 15334 31108 15372
rect 31388 15428 31444 15932
rect 31836 15540 31892 16942
rect 32508 16772 32564 17614
rect 32620 17556 32676 17566
rect 32620 17106 32676 17500
rect 32844 17444 32900 17454
rect 32844 17350 32900 17388
rect 33628 17444 33684 17454
rect 35532 17444 35588 17454
rect 33628 17442 34468 17444
rect 33628 17390 33630 17442
rect 33682 17390 34468 17442
rect 33628 17388 34468 17390
rect 33628 17378 33684 17388
rect 32620 17054 32622 17106
rect 32674 17054 32676 17106
rect 32620 17042 32676 17054
rect 32060 15874 32116 15886
rect 32060 15822 32062 15874
rect 32114 15822 32116 15874
rect 31836 15474 31892 15484
rect 31948 15652 32004 15662
rect 31724 15428 31780 15438
rect 31388 15426 31724 15428
rect 31388 15374 31390 15426
rect 31442 15374 31724 15426
rect 31388 15372 31724 15374
rect 31388 15362 31444 15372
rect 31724 15334 31780 15372
rect 31948 13858 32004 15596
rect 32060 15426 32116 15822
rect 32508 15538 32564 16716
rect 33180 16882 33236 16894
rect 33180 16830 33182 16882
rect 33234 16830 33236 16882
rect 33180 16772 33236 16830
rect 33068 16100 33124 16110
rect 33180 16100 33236 16716
rect 33628 16882 33684 16894
rect 33628 16830 33630 16882
rect 33682 16830 33684 16882
rect 33068 16098 33236 16100
rect 33068 16046 33070 16098
rect 33122 16046 33236 16098
rect 33068 16044 33236 16046
rect 33068 16034 33124 16044
rect 32508 15486 32510 15538
rect 32562 15486 32564 15538
rect 32508 15474 32564 15486
rect 32732 15874 32788 15886
rect 32732 15822 32734 15874
rect 32786 15822 32788 15874
rect 32060 15374 32062 15426
rect 32114 15374 32116 15426
rect 32060 15362 32116 15374
rect 31948 13806 31950 13858
rect 32002 13806 32004 13858
rect 31948 13794 32004 13806
rect 32508 14530 32564 14542
rect 32508 14478 32510 14530
rect 32562 14478 32564 14530
rect 30940 13582 30942 13634
rect 30994 13582 30996 13634
rect 30940 13570 30996 13582
rect 31164 12852 31220 12862
rect 31164 12758 31220 12796
rect 30380 12238 30382 12290
rect 30434 12238 30436 12290
rect 30380 12226 30436 12238
rect 29036 12068 29092 12078
rect 29036 11974 29092 12012
rect 32508 12068 32564 14478
rect 32732 13524 32788 15822
rect 33068 15428 33124 15438
rect 33068 15334 33124 15372
rect 33068 14532 33124 14542
rect 33180 14532 33236 16044
rect 33516 16098 33572 16110
rect 33516 16046 33518 16098
rect 33570 16046 33572 16098
rect 33292 15316 33348 15326
rect 33292 15222 33348 15260
rect 33068 14530 33236 14532
rect 33068 14478 33070 14530
rect 33122 14478 33236 14530
rect 33068 14476 33236 14478
rect 33068 14466 33124 14476
rect 33516 14308 33572 16046
rect 33628 14980 33684 16830
rect 34412 15426 34468 17388
rect 34412 15374 34414 15426
rect 34466 15374 34468 15426
rect 34412 15362 34468 15374
rect 34972 16772 35028 16782
rect 33740 15316 33796 15326
rect 33740 15222 33796 15260
rect 34972 15314 35028 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34972 15250 35028 15262
rect 33964 15204 34020 15214
rect 33964 15110 34020 15148
rect 34748 15204 34804 15214
rect 34748 15110 34804 15148
rect 33628 14924 34468 14980
rect 34300 14644 34356 14654
rect 34300 14550 34356 14588
rect 33516 14242 33572 14252
rect 34300 14308 34356 14318
rect 32732 13458 32788 13468
rect 34300 13074 34356 14252
rect 34412 13634 34468 14924
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35308 14420 35364 14430
rect 35308 14326 35364 14364
rect 35532 13972 35588 17388
rect 35644 15314 35700 15326
rect 35644 15262 35646 15314
rect 35698 15262 35700 15314
rect 35644 14196 35700 15262
rect 35644 14130 35700 14140
rect 35532 13916 35700 13972
rect 34412 13582 34414 13634
rect 34466 13582 34468 13634
rect 34412 13570 34468 13582
rect 35420 13524 35476 13534
rect 35476 13468 35588 13524
rect 35420 13458 35476 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34300 13022 34302 13074
rect 34354 13022 34356 13074
rect 34300 13010 34356 13022
rect 34860 12740 34916 12750
rect 32508 12002 32564 12012
rect 34076 12068 34132 12078
rect 34076 11974 34132 12012
rect 33516 11508 33572 11518
rect 33516 11414 33572 11452
rect 28028 11230 28030 11282
rect 28082 11230 28084 11282
rect 28028 11218 28084 11230
rect 34860 11282 34916 12684
rect 35420 12292 35476 12302
rect 35532 12292 35588 13468
rect 35644 12850 35700 13916
rect 35756 13858 35812 18956
rect 35980 17780 36036 17790
rect 35980 17666 36036 17724
rect 35980 17614 35982 17666
rect 36034 17614 36036 17666
rect 35980 17602 36036 17614
rect 36092 17106 36148 18956
rect 36204 18452 36260 20078
rect 37212 19908 37268 20860
rect 37324 20914 37380 21532
rect 37436 21252 37492 21756
rect 37548 21476 37604 22318
rect 38444 21700 38500 23996
rect 38780 23938 38836 25564
rect 38892 25060 38948 26126
rect 38892 24994 38948 25004
rect 39340 24834 39396 27916
rect 39676 27906 39732 27916
rect 40012 26850 40068 26862
rect 40012 26798 40014 26850
rect 40066 26798 40068 26850
rect 39340 24782 39342 24834
rect 39394 24782 39396 24834
rect 39340 24770 39396 24782
rect 39788 26402 39844 26414
rect 39788 26350 39790 26402
rect 39842 26350 39844 26402
rect 39004 24724 39060 24734
rect 39004 24610 39060 24668
rect 39676 24724 39732 24734
rect 39676 24630 39732 24668
rect 39004 24558 39006 24610
rect 39058 24558 39060 24610
rect 39004 24052 39060 24558
rect 39004 23986 39060 23996
rect 38780 23886 38782 23938
rect 38834 23886 38836 23938
rect 38780 23874 38836 23886
rect 39788 23492 39844 26350
rect 40012 24834 40068 26798
rect 40124 26516 40180 28364
rect 40572 28418 40628 28430
rect 40572 28366 40574 28418
rect 40626 28366 40628 28418
rect 40460 27972 40516 27982
rect 40460 27878 40516 27916
rect 40572 27636 40628 28366
rect 40572 27570 40628 27580
rect 40572 27300 40628 27310
rect 40684 27300 40740 28476
rect 40796 28466 40852 28476
rect 42812 28532 42868 28542
rect 42812 28438 42868 28476
rect 42924 27972 42980 27982
rect 42924 27878 42980 27916
rect 41916 27748 41972 27758
rect 41916 27654 41972 27692
rect 40572 27298 40740 27300
rect 40572 27246 40574 27298
rect 40626 27246 40740 27298
rect 40572 27244 40740 27246
rect 42812 27636 42868 27646
rect 40572 27234 40628 27244
rect 41804 27188 41860 27198
rect 41804 27094 41860 27132
rect 40124 26450 40180 26460
rect 40684 26964 40740 26974
rect 40684 25282 40740 26908
rect 42812 26962 42868 27580
rect 42812 26910 42814 26962
rect 42866 26910 42868 26962
rect 42812 26898 42868 26910
rect 43596 26962 43652 26974
rect 43596 26910 43598 26962
rect 43650 26910 43652 26962
rect 42924 26404 42980 26414
rect 42924 26310 42980 26348
rect 41916 26180 41972 26190
rect 41916 26086 41972 26124
rect 43596 26180 43652 26910
rect 43932 26964 43988 26974
rect 43932 26870 43988 26908
rect 43820 26516 43876 26526
rect 43820 26422 43876 26460
rect 43708 26180 43764 26190
rect 43596 26178 43764 26180
rect 43596 26126 43710 26178
rect 43762 26126 43764 26178
rect 43596 26124 43764 26126
rect 42476 25620 42532 25630
rect 42476 25526 42532 25564
rect 41244 25396 41300 25406
rect 41244 25302 41300 25340
rect 40684 25230 40686 25282
rect 40738 25230 40740 25282
rect 40684 25218 40740 25230
rect 40012 24782 40014 24834
rect 40066 24782 40068 24834
rect 40012 24770 40068 24782
rect 43148 24834 43204 24846
rect 43148 24782 43150 24834
rect 43202 24782 43204 24834
rect 41916 24612 41972 24622
rect 41916 24518 41972 24556
rect 42252 24052 42308 24062
rect 42252 23938 42308 23996
rect 42252 23886 42254 23938
rect 42306 23886 42308 23938
rect 42252 23874 42308 23886
rect 41244 23828 41300 23838
rect 41244 23714 41300 23772
rect 42028 23828 42084 23838
rect 42028 23734 42084 23772
rect 41804 23716 41860 23726
rect 41244 23662 41246 23714
rect 41298 23662 41300 23714
rect 41244 23650 41300 23662
rect 41580 23714 41860 23716
rect 41580 23662 41806 23714
rect 41858 23662 41860 23714
rect 41580 23660 41860 23662
rect 39788 23426 39844 23436
rect 39676 23266 39732 23278
rect 39676 23214 39678 23266
rect 39730 23214 39732 23266
rect 38444 21606 38500 21644
rect 39452 21700 39508 21710
rect 39452 21606 39508 21644
rect 38108 21588 38164 21598
rect 37548 21410 37604 21420
rect 37772 21586 38164 21588
rect 37772 21534 38110 21586
rect 38162 21534 38164 21586
rect 37772 21532 38164 21534
rect 37772 21252 37828 21532
rect 38108 21522 38164 21532
rect 38780 21474 38836 21486
rect 38780 21422 38782 21474
rect 38834 21422 38836 21474
rect 37884 21364 37940 21374
rect 37884 21270 37940 21308
rect 37436 21196 37828 21252
rect 37324 20862 37326 20914
rect 37378 20862 37380 20914
rect 37324 20850 37380 20862
rect 38444 20916 38500 20926
rect 37772 20802 37828 20814
rect 37772 20750 37774 20802
rect 37826 20750 37828 20802
rect 37324 19908 37380 19918
rect 37212 19906 37380 19908
rect 37212 19854 37326 19906
rect 37378 19854 37380 19906
rect 37212 19852 37380 19854
rect 36988 19796 37044 19806
rect 36988 19794 37156 19796
rect 36988 19742 36990 19794
rect 37042 19742 37156 19794
rect 36988 19740 37156 19742
rect 36988 19730 37044 19740
rect 36204 18386 36260 18396
rect 36540 19236 36596 19246
rect 36540 18338 36596 19180
rect 36540 18286 36542 18338
rect 36594 18286 36596 18338
rect 36540 17668 36596 18286
rect 36988 17668 37044 17678
rect 36540 17666 37044 17668
rect 36540 17614 36542 17666
rect 36594 17614 36990 17666
rect 37042 17614 37044 17666
rect 36540 17612 37044 17614
rect 36540 17602 36596 17612
rect 36092 17054 36094 17106
rect 36146 17054 36148 17106
rect 36092 17042 36148 17054
rect 36652 17444 36708 17454
rect 36652 17106 36708 17388
rect 36652 17054 36654 17106
rect 36706 17054 36708 17106
rect 36652 17042 36708 17054
rect 36988 16884 37044 17612
rect 37100 16996 37156 19740
rect 37212 19234 37268 19852
rect 37324 19842 37380 19852
rect 37212 19182 37214 19234
rect 37266 19182 37268 19234
rect 37212 19170 37268 19182
rect 37772 19236 37828 20750
rect 38444 20802 38500 20860
rect 38444 20750 38446 20802
rect 38498 20750 38500 20802
rect 38444 20738 38500 20750
rect 38780 20804 38836 21422
rect 38780 20738 38836 20748
rect 39116 21474 39172 21486
rect 39116 21422 39118 21474
rect 39170 21422 39172 21474
rect 39116 20188 39172 21422
rect 39676 21474 39732 23214
rect 40460 22930 40516 22942
rect 40460 22878 40462 22930
rect 40514 22878 40516 22930
rect 40012 22260 40068 22270
rect 40012 22146 40068 22204
rect 40012 22094 40014 22146
rect 40066 22094 40068 22146
rect 40012 22082 40068 22094
rect 40460 21700 40516 22878
rect 40460 21634 40516 21644
rect 40572 22146 40628 22158
rect 40572 22094 40574 22146
rect 40626 22094 40628 22146
rect 39676 21422 39678 21474
rect 39730 21422 39732 21474
rect 39676 21410 39732 21422
rect 40572 20692 40628 22094
rect 40572 20626 40628 20636
rect 40908 22148 40964 22158
rect 40908 20578 40964 22092
rect 41468 22146 41524 22158
rect 41468 22094 41470 22146
rect 41522 22094 41524 22146
rect 41468 21588 41524 22094
rect 41468 21522 41524 21532
rect 40908 20526 40910 20578
rect 40962 20526 40964 20578
rect 40908 20514 40964 20526
rect 41468 20578 41524 20590
rect 41468 20526 41470 20578
rect 41522 20526 41524 20578
rect 38892 20132 39172 20188
rect 38220 19908 38276 19918
rect 38220 19814 38276 19852
rect 37884 19348 37940 19358
rect 37884 19254 37940 19292
rect 38892 19348 38948 20132
rect 39228 20130 39284 20142
rect 39228 20078 39230 20130
rect 39282 20078 39284 20130
rect 39228 19796 39284 20078
rect 39228 19730 39284 19740
rect 37772 19170 37828 19180
rect 38892 19122 38948 19292
rect 39116 19236 39172 19246
rect 39116 19142 39172 19180
rect 39788 19234 39844 19246
rect 39788 19182 39790 19234
rect 39842 19182 39844 19234
rect 38892 19070 38894 19122
rect 38946 19070 38948 19122
rect 38780 19012 38836 19022
rect 38780 18918 38836 18956
rect 38780 18452 38836 18462
rect 38892 18452 38948 19070
rect 39788 18564 39844 19182
rect 39788 18498 39844 18508
rect 38780 18450 38948 18452
rect 38780 18398 38782 18450
rect 38834 18398 38948 18450
rect 38780 18396 38948 18398
rect 39340 18452 39396 18462
rect 38780 18340 38836 18396
rect 39340 18358 39396 18396
rect 39564 18450 39620 18462
rect 39564 18398 39566 18450
rect 39618 18398 39620 18450
rect 37548 17666 37604 17678
rect 37548 17614 37550 17666
rect 37602 17614 37604 17666
rect 37100 16930 37156 16940
rect 37212 17108 37268 17118
rect 36988 16790 37044 16828
rect 35980 15874 36036 15886
rect 35980 15822 35982 15874
rect 36034 15822 36036 15874
rect 35980 14644 36036 15822
rect 36540 15874 36596 15886
rect 36540 15822 36542 15874
rect 36594 15822 36596 15874
rect 36316 15204 36372 15214
rect 36092 14644 36148 14654
rect 35980 14642 36148 14644
rect 35980 14590 36094 14642
rect 36146 14590 36148 14642
rect 35980 14588 36148 14590
rect 36092 14578 36148 14588
rect 36316 14530 36372 15148
rect 36316 14478 36318 14530
rect 36370 14478 36372 14530
rect 36316 14466 36372 14478
rect 36540 14308 36596 15822
rect 36876 15874 36932 15886
rect 36876 15822 36878 15874
rect 36930 15822 36932 15874
rect 36876 14868 36932 15822
rect 36876 14802 36932 14812
rect 36540 14242 36596 14252
rect 36876 14306 36932 14318
rect 36876 14254 36878 14306
rect 36930 14254 36932 14306
rect 35756 13806 35758 13858
rect 35810 13806 35812 13858
rect 35756 13794 35812 13806
rect 35644 12798 35646 12850
rect 35698 12798 35700 12850
rect 35644 12786 35700 12798
rect 36876 12740 36932 14254
rect 37212 13634 37268 17052
rect 37436 16882 37492 16894
rect 37436 16830 37438 16882
rect 37490 16830 37492 16882
rect 37436 16212 37492 16830
rect 37548 16772 37604 17614
rect 37548 16706 37604 16716
rect 37436 16146 37492 16156
rect 37660 16660 37716 16670
rect 37660 15986 37716 16604
rect 37660 15934 37662 15986
rect 37714 15934 37716 15986
rect 37660 15922 37716 15934
rect 38108 15538 38164 15550
rect 38108 15486 38110 15538
rect 38162 15486 38164 15538
rect 38108 15428 38164 15486
rect 38108 15362 38164 15372
rect 38780 15204 38836 18284
rect 39004 18340 39060 18350
rect 39564 18340 39620 18398
rect 40236 18450 40292 18462
rect 40236 18398 40238 18450
rect 40290 18398 40292 18450
rect 39004 18338 39284 18340
rect 39004 18286 39006 18338
rect 39058 18286 39284 18338
rect 39004 18284 39284 18286
rect 39004 18274 39060 18284
rect 39228 17892 39284 18284
rect 39564 18274 39620 18284
rect 40012 18338 40068 18350
rect 40012 18286 40014 18338
rect 40066 18286 40068 18338
rect 39228 17836 39844 17892
rect 39788 17554 39844 17836
rect 39788 17502 39790 17554
rect 39842 17502 39844 17554
rect 39788 17490 39844 17502
rect 39900 17108 39956 17118
rect 40012 17108 40068 18286
rect 40236 18340 40292 18398
rect 40236 18274 40292 18284
rect 39900 17106 40068 17108
rect 39900 17054 39902 17106
rect 39954 17054 40068 17106
rect 39900 17052 40068 17054
rect 40572 17442 40628 17454
rect 40572 17390 40574 17442
rect 40626 17390 40628 17442
rect 39900 17042 39956 17052
rect 40348 16884 40404 16894
rect 40012 16098 40068 16110
rect 40012 16046 40014 16098
rect 40066 16046 40068 16098
rect 38892 15428 38948 15438
rect 38892 15334 38948 15372
rect 38780 15138 38836 15148
rect 39116 15314 39172 15326
rect 39116 15262 39118 15314
rect 39170 15262 39172 15314
rect 39116 15204 39172 15262
rect 39116 15138 39172 15148
rect 38668 15090 38724 15102
rect 38668 15038 38670 15090
rect 38722 15038 38724 15090
rect 38220 14868 38276 14878
rect 37660 14420 37716 14430
rect 37660 14326 37716 14364
rect 37212 13582 37214 13634
rect 37266 13582 37268 13634
rect 37212 13570 37268 13582
rect 37996 14196 38052 14206
rect 37996 13074 38052 14140
rect 38220 13858 38276 14812
rect 38668 13972 38724 15038
rect 40012 15092 40068 16046
rect 40012 15026 40068 15036
rect 40348 16098 40404 16828
rect 40348 16046 40350 16098
rect 40402 16046 40404 16098
rect 40012 14530 40068 14542
rect 40012 14478 40014 14530
rect 40066 14478 40068 14530
rect 38668 13906 38724 13916
rect 39004 14308 39060 14318
rect 38220 13806 38222 13858
rect 38274 13806 38276 13858
rect 38220 13794 38276 13806
rect 37996 13022 37998 13074
rect 38050 13022 38052 13074
rect 37996 13010 38052 13022
rect 39004 12850 39060 14252
rect 40012 13076 40068 14478
rect 40348 14530 40404 16046
rect 40460 16658 40516 16670
rect 40460 16606 40462 16658
rect 40514 16606 40516 16658
rect 40460 15204 40516 16606
rect 40572 15988 40628 17390
rect 40572 15922 40628 15932
rect 41468 15428 41524 20526
rect 41580 20132 41636 23660
rect 41804 23650 41860 23660
rect 42812 23716 42868 23726
rect 41916 23044 41972 23054
rect 41916 22950 41972 22988
rect 41804 22482 41860 22494
rect 41804 22430 41806 22482
rect 41858 22430 41860 22482
rect 41804 21812 41860 22430
rect 42812 22258 42868 23660
rect 42924 23716 42980 23726
rect 42924 23714 43092 23716
rect 42924 23662 42926 23714
rect 42978 23662 43092 23714
rect 42924 23660 43092 23662
rect 42924 23650 42980 23660
rect 42924 23266 42980 23278
rect 42924 23214 42926 23266
rect 42978 23214 42980 23266
rect 42924 22596 42980 23214
rect 42924 22530 42980 22540
rect 42812 22206 42814 22258
rect 42866 22206 42868 22258
rect 42812 22194 42868 22206
rect 43036 21924 43092 23660
rect 41804 21746 41860 21756
rect 42812 21868 43092 21924
rect 42476 21588 42532 21598
rect 41916 21476 41972 21486
rect 41916 21382 41972 21420
rect 42252 21476 42308 21486
rect 41580 20066 41636 20076
rect 41916 19906 41972 19918
rect 41916 19854 41918 19906
rect 41970 19854 41972 19906
rect 41916 19572 41972 19854
rect 41916 19506 41972 19516
rect 41916 19124 41972 19134
rect 41692 18564 41748 18574
rect 41692 16548 41748 18508
rect 41916 18338 41972 19068
rect 42252 19010 42308 21420
rect 42476 20914 42532 21532
rect 42476 20862 42478 20914
rect 42530 20862 42532 20914
rect 42476 20850 42532 20862
rect 42700 20916 42756 20926
rect 42700 20822 42756 20860
rect 42812 19458 42868 21868
rect 42924 21700 42980 21710
rect 42924 21606 42980 21644
rect 43148 21364 43204 24782
rect 43484 24050 43540 24062
rect 43484 23998 43486 24050
rect 43538 23998 43540 24050
rect 43484 22372 43540 23998
rect 43596 24052 43652 26124
rect 43708 26114 43764 26124
rect 43708 25396 43764 25406
rect 43708 25302 43764 25340
rect 43596 23548 43652 23996
rect 43596 23492 43764 23548
rect 43708 23266 43764 23492
rect 43708 23214 43710 23266
rect 43762 23214 43764 23266
rect 43708 23202 43764 23214
rect 43484 22306 43540 22316
rect 43932 23042 43988 23054
rect 43932 22990 43934 23042
rect 43986 22990 43988 23042
rect 43596 22258 43652 22270
rect 43596 22206 43598 22258
rect 43650 22206 43652 22258
rect 43596 21588 43652 22206
rect 43932 22260 43988 22990
rect 43932 22194 43988 22204
rect 43708 22148 43764 22158
rect 43708 22054 43764 22092
rect 43708 21588 43764 21598
rect 43652 21586 43764 21588
rect 43652 21534 43710 21586
rect 43762 21534 43764 21586
rect 43652 21532 43764 21534
rect 43596 21494 43652 21532
rect 43708 21522 43764 21532
rect 43932 21476 43988 21486
rect 43932 21382 43988 21420
rect 43148 21298 43204 21308
rect 43708 20692 43764 20702
rect 43708 20598 43764 20636
rect 42924 20132 42980 20142
rect 42924 20038 42980 20076
rect 42812 19406 42814 19458
rect 42866 19406 42868 19458
rect 42812 19394 42868 19406
rect 42252 18958 42254 19010
rect 42306 18958 42308 19010
rect 42252 18946 42308 18958
rect 41916 18286 41918 18338
rect 41970 18286 41972 18338
rect 41916 18274 41972 18286
rect 42924 18562 42980 18574
rect 42924 18510 42926 18562
rect 42978 18510 42980 18562
rect 41804 17780 41860 17790
rect 41804 17686 41860 17724
rect 42812 17556 42868 17566
rect 42812 17462 42868 17500
rect 42924 17444 42980 18510
rect 43596 18340 43652 18350
rect 43596 17780 43652 18284
rect 43596 17778 43764 17780
rect 43596 17726 43598 17778
rect 43650 17726 43764 17778
rect 43596 17724 43764 17726
rect 43596 17686 43652 17724
rect 42924 17378 42980 17388
rect 42924 16996 42980 17006
rect 42924 16902 42980 16940
rect 43708 16994 43764 17724
rect 43708 16942 43710 16994
rect 43762 16942 43764 16994
rect 43708 16930 43764 16942
rect 43932 17554 43988 17566
rect 43932 17502 43934 17554
rect 43986 17502 43988 17554
rect 41916 16772 41972 16782
rect 41916 16678 41972 16716
rect 43932 16660 43988 17502
rect 43932 16594 43988 16604
rect 44044 16770 44100 16782
rect 44044 16718 44046 16770
rect 44098 16718 44100 16770
rect 41692 16492 41972 16548
rect 41804 16212 41860 16222
rect 41804 16118 41860 16156
rect 41468 15362 41524 15372
rect 40460 15138 40516 15148
rect 41916 15202 41972 16492
rect 42812 15988 42868 15998
rect 42812 15894 42868 15932
rect 42924 15428 42980 15438
rect 42924 15334 42980 15372
rect 41916 15150 41918 15202
rect 41970 15150 41972 15202
rect 41916 15138 41972 15150
rect 42924 15204 42980 15214
rect 41804 15092 41860 15102
rect 41804 14642 41860 15036
rect 41804 14590 41806 14642
rect 41858 14590 41860 14642
rect 41804 14578 41860 14590
rect 40348 14478 40350 14530
rect 40402 14478 40404 14530
rect 40348 14466 40404 14478
rect 42924 14418 42980 15148
rect 42924 14366 42926 14418
rect 42978 14366 42980 14418
rect 42924 14354 42980 14366
rect 44044 14420 44100 16718
rect 44044 14354 44100 14364
rect 42028 13972 42084 13982
rect 40012 13010 40068 13020
rect 40796 13076 40852 13086
rect 40796 12982 40852 13020
rect 39004 12798 39006 12850
rect 39058 12798 39060 12850
rect 39004 12786 39060 12798
rect 42028 12850 42084 13916
rect 42028 12798 42030 12850
rect 42082 12798 42084 12850
rect 42028 12786 42084 12798
rect 36876 12674 36932 12684
rect 35420 12290 35588 12292
rect 35420 12238 35422 12290
rect 35474 12238 35588 12290
rect 35420 12236 35588 12238
rect 35420 12226 35476 12236
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34860 11230 34862 11282
rect 34914 11230 34916 11282
rect 34860 11218 34916 11230
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20076 9154 20132 9166
rect 20076 9102 20078 9154
rect 20130 9102 20132 9154
rect 19740 9042 19796 9054
rect 19740 8990 19742 9042
rect 19794 8990 19796 9042
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 19740 8428 19796 8990
rect 19628 8372 19796 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19628 4564 19684 8372
rect 20076 8036 20132 9102
rect 20860 9154 20916 9166
rect 20860 9102 20862 9154
rect 20914 9102 20916 9154
rect 20636 9042 20692 9054
rect 20636 8990 20638 9042
rect 20690 8990 20692 9042
rect 20636 8428 20692 8990
rect 20860 8428 20916 9102
rect 43820 9154 43876 9166
rect 43820 9102 43822 9154
rect 43874 9102 43876 9154
rect 43596 8932 43652 8942
rect 43596 8838 43652 8876
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 20636 8372 20804 8428
rect 20860 8372 21140 8428
rect 20076 7980 20244 8036
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20188 7700 20244 7980
rect 20076 7644 20244 7700
rect 20076 6468 20132 7644
rect 20076 6412 20244 6468
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6412
rect 20076 6076 20244 6132
rect 20076 4900 20132 6076
rect 20076 4844 20244 4900
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20076 4564 20132 4574
rect 19628 4562 20132 4564
rect 19628 4510 20078 4562
rect 20130 4510 20132 4562
rect 19628 4508 20132 4510
rect 20076 4498 20132 4508
rect 19068 4452 19124 4462
rect 19068 4450 19796 4452
rect 19068 4398 19070 4450
rect 19122 4398 19796 4450
rect 19068 4396 19796 4398
rect 19068 4386 19124 4396
rect 19740 4338 19796 4396
rect 20188 4340 20244 4844
rect 20748 4562 20804 8372
rect 20748 4510 20750 4562
rect 20802 4510 20804 4562
rect 20748 4498 20804 4510
rect 19740 4286 19742 4338
rect 19794 4286 19796 4338
rect 19516 4228 19572 4238
rect 19516 4134 19572 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 19404 3332 19460 3342
rect 19740 3332 19796 4286
rect 20076 4284 20244 4340
rect 20412 4338 20468 4350
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20076 3554 20132 4284
rect 20076 3502 20078 3554
rect 20130 3502 20132 3554
rect 20076 3490 20132 3502
rect 20188 4116 20244 4126
rect 20412 4116 20468 4286
rect 20244 4060 20468 4116
rect 18844 3330 19460 3332
rect 18844 3278 19406 3330
rect 19458 3278 19460 3330
rect 18844 3276 19460 3278
rect 18844 800 18900 3276
rect 19404 3266 19460 3276
rect 19516 3276 19796 3332
rect 19516 800 19572 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 4060
rect 21084 3554 21140 8372
rect 27020 8260 27076 8270
rect 42924 8260 42980 8270
rect 27020 8258 27188 8260
rect 27020 8206 27022 8258
rect 27074 8206 27188 8258
rect 27020 8204 27188 8206
rect 27020 8194 27076 8204
rect 24444 6580 24500 6590
rect 23996 6578 24500 6580
rect 23996 6526 24446 6578
rect 24498 6526 24500 6578
rect 23996 6524 24500 6526
rect 21532 3668 21588 3678
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 21196 3666 21588 3668
rect 21196 3614 21534 3666
rect 21586 3614 21588 3666
rect 21196 3612 21588 3614
rect 21196 1764 21252 3612
rect 21532 3602 21588 3612
rect 23772 3554 23828 3566
rect 23772 3502 23774 3554
rect 23826 3502 23828 3554
rect 20860 1708 21252 1764
rect 21532 3332 21588 3342
rect 20860 800 20916 1708
rect 21532 800 21588 3276
rect 22652 3332 22708 3342
rect 23660 3332 23716 3342
rect 22652 3238 22708 3276
rect 23548 3276 23660 3332
rect 23548 800 23604 3276
rect 23660 3266 23716 3276
rect 23772 2548 23828 3502
rect 23996 3442 24052 6524
rect 24444 6514 24500 6524
rect 24780 6468 24836 6478
rect 24780 6466 25060 6468
rect 24780 6414 24782 6466
rect 24834 6414 25060 6466
rect 24780 6412 25060 6414
rect 24780 6402 24836 6412
rect 25004 4452 25060 6412
rect 25116 5122 25172 5134
rect 25116 5070 25118 5122
rect 25170 5070 25172 5122
rect 25116 4564 25172 5070
rect 25340 4900 25396 4910
rect 25340 4898 26180 4900
rect 25340 4846 25342 4898
rect 25394 4846 26180 4898
rect 25340 4844 26180 4846
rect 25340 4834 25396 4844
rect 25228 4564 25284 4574
rect 25116 4562 25284 4564
rect 25116 4510 25230 4562
rect 25282 4510 25284 4562
rect 25116 4508 25284 4510
rect 25228 4498 25284 4508
rect 25004 4396 25172 4452
rect 24892 4340 24948 4350
rect 25116 4340 25172 4396
rect 25564 4340 25620 4350
rect 25116 4284 25284 4340
rect 23996 3390 23998 3442
rect 24050 3390 24052 3442
rect 23996 3378 24052 3390
rect 24220 4226 24276 4238
rect 24220 4174 24222 4226
rect 24274 4174 24276 4226
rect 24220 2548 24276 4174
rect 24780 4228 24836 4238
rect 24892 4228 24948 4284
rect 24780 4226 24948 4228
rect 24780 4174 24782 4226
rect 24834 4174 24948 4226
rect 24780 4172 24948 4174
rect 24780 4162 24836 4172
rect 24556 3332 24612 3342
rect 24556 3238 24612 3276
rect 23772 2492 24276 2548
rect 24220 800 24276 2492
rect 24892 800 24948 4172
rect 25228 3554 25284 4284
rect 25564 4246 25620 4284
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3490 25284 3502
rect 25564 3668 25620 3678
rect 25564 800 25620 3612
rect 26124 3554 26180 4844
rect 27132 4562 27188 8204
rect 42476 8258 42980 8260
rect 42476 8206 42926 8258
rect 42978 8206 42980 8258
rect 42476 8204 42980 8206
rect 27244 8036 27300 8046
rect 27244 8034 28420 8036
rect 27244 7982 27246 8034
rect 27298 7982 28420 8034
rect 27244 7980 28420 7982
rect 27244 7970 27300 7980
rect 27132 4510 27134 4562
rect 27186 4510 27188 4562
rect 27132 4498 27188 4510
rect 26460 4450 26516 4462
rect 26460 4398 26462 4450
rect 26514 4398 26516 4450
rect 26236 4228 26292 4238
rect 26236 4134 26292 4172
rect 26124 3502 26126 3554
rect 26178 3502 26180 3554
rect 26124 3490 26180 3502
rect 26460 1092 26516 4398
rect 27356 4338 27412 4350
rect 27356 4286 27358 4338
rect 27410 4286 27412 4338
rect 27356 4228 27412 4286
rect 26572 3668 26628 3678
rect 26572 3574 26628 3612
rect 27356 3388 27412 4172
rect 26236 1036 26516 1092
rect 26908 3332 27412 3388
rect 27580 3668 27636 3678
rect 26236 800 26292 1036
rect 26908 800 26964 3332
rect 27580 800 27636 3612
rect 28364 3554 28420 7980
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 41804 5908 41860 5918
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35756 5236 35812 5246
rect 33404 5124 33460 5134
rect 33404 5122 33572 5124
rect 33404 5070 33406 5122
rect 33458 5070 33572 5122
rect 33404 5068 33572 5070
rect 33404 5058 33460 5068
rect 31836 5012 31892 5022
rect 31500 5010 31892 5012
rect 31500 4958 31838 5010
rect 31890 4958 31892 5010
rect 31500 4956 31892 4958
rect 28812 3668 28868 3678
rect 28812 3574 28868 3612
rect 28364 3502 28366 3554
rect 28418 3502 28420 3554
rect 28364 3490 28420 3502
rect 30940 3444 30996 3454
rect 31164 3444 31220 3454
rect 30940 3442 31220 3444
rect 30940 3390 30942 3442
rect 30994 3390 31166 3442
rect 31218 3390 31220 3442
rect 30940 3388 31220 3390
rect 30940 800 30996 3388
rect 31164 3378 31220 3388
rect 31500 3442 31556 4956
rect 31836 4946 31892 4956
rect 32172 4900 32228 4910
rect 32060 4898 32228 4900
rect 32060 4846 32174 4898
rect 32226 4846 32228 4898
rect 32060 4844 32228 4846
rect 31500 3390 31502 3442
rect 31554 3390 31556 3442
rect 31500 3378 31556 3390
rect 31612 3668 31668 3678
rect 31612 800 31668 3612
rect 32060 3556 32116 4844
rect 32172 4834 32228 4844
rect 33516 4562 33572 5068
rect 33628 4900 33684 4910
rect 33628 4898 33908 4900
rect 33628 4846 33630 4898
rect 33682 4846 33908 4898
rect 33628 4844 33908 4846
rect 33628 4834 33684 4844
rect 33516 4510 33518 4562
rect 33570 4510 33572 4562
rect 33516 4498 33572 4510
rect 32396 4452 32452 4462
rect 32284 4450 32452 4452
rect 32284 4398 32398 4450
rect 32450 4398 32452 4450
rect 32284 4396 32452 4398
rect 32172 4228 32228 4238
rect 32172 4134 32228 4172
rect 32172 3556 32228 3566
rect 32060 3554 32228 3556
rect 32060 3502 32174 3554
rect 32226 3502 32228 3554
rect 32060 3500 32228 3502
rect 32172 3490 32228 3500
rect 32284 800 32340 4396
rect 32396 4386 32452 4396
rect 33180 4338 33236 4350
rect 33180 4286 33182 4338
rect 33234 4286 33236 4338
rect 32956 4228 33012 4238
rect 32956 3892 33012 4172
rect 33180 3892 33236 4286
rect 32956 3836 33236 3892
rect 32620 3668 32676 3678
rect 32620 3574 32676 3612
rect 32956 800 33012 3836
rect 33852 3554 33908 4844
rect 35756 4562 35812 5180
rect 37884 5236 37940 5246
rect 36428 5124 36484 5134
rect 37436 5124 37492 5134
rect 35756 4510 35758 4562
rect 35810 4510 35812 4562
rect 35756 4498 35812 4510
rect 35868 4898 35924 4910
rect 35868 4846 35870 4898
rect 35922 4846 35924 4898
rect 35868 4340 35924 4846
rect 36428 4562 36484 5068
rect 37100 5122 37492 5124
rect 37100 5070 37438 5122
rect 37490 5070 37492 5122
rect 37100 5068 37492 5070
rect 36428 4510 36430 4562
rect 36482 4510 36484 4562
rect 36428 4498 36484 4510
rect 36540 4898 36596 4910
rect 36540 4846 36542 4898
rect 36594 4846 36596 4898
rect 36092 4340 36148 4350
rect 35868 4338 36148 4340
rect 35868 4286 36094 4338
rect 36146 4286 36148 4338
rect 35868 4284 36148 4286
rect 36540 4340 36596 4846
rect 37100 4562 37156 5068
rect 37436 5058 37492 5068
rect 37884 5010 37940 5180
rect 38108 5124 38164 5134
rect 38108 5030 38164 5068
rect 38668 5124 38724 5134
rect 38668 5122 38836 5124
rect 38668 5070 38670 5122
rect 38722 5070 38836 5122
rect 38668 5068 38836 5070
rect 38668 5058 38724 5068
rect 37884 4958 37886 5010
rect 37938 4958 37940 5010
rect 37884 4946 37940 4958
rect 37100 4510 37102 4562
rect 37154 4510 37156 4562
rect 37100 4498 37156 4510
rect 37212 4898 37268 4910
rect 37212 4846 37214 4898
rect 37266 4846 37268 4898
rect 36764 4340 36820 4350
rect 36540 4338 36820 4340
rect 36540 4286 36766 4338
rect 36818 4286 36820 4338
rect 36540 4284 36820 4286
rect 34972 4116 35028 4126
rect 34748 4114 35028 4116
rect 34748 4062 34974 4114
rect 35026 4062 35028 4114
rect 34748 4060 35028 4062
rect 34300 3668 34356 3678
rect 33852 3502 33854 3554
rect 33906 3502 33908 3554
rect 33852 3490 33908 3502
rect 34076 3666 34356 3668
rect 34076 3614 34302 3666
rect 34354 3614 34356 3666
rect 34076 3612 34356 3614
rect 34076 3388 34132 3612
rect 34300 3602 34356 3612
rect 34748 3388 34804 4060
rect 34972 4050 35028 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 33852 3332 34132 3388
rect 34300 3332 34804 3388
rect 34972 3556 35028 3566
rect 33852 980 33908 3332
rect 33628 924 33908 980
rect 33628 800 33684 924
rect 34300 800 34356 3332
rect 34972 800 35028 3500
rect 36092 3556 36148 4284
rect 36092 3490 36148 3500
rect 36764 3388 36820 4284
rect 37212 3554 37268 4846
rect 38780 4564 38836 5068
rect 39228 5012 39284 5022
rect 39228 4918 39284 4956
rect 40908 5012 40964 5022
rect 38892 4900 38948 4910
rect 38892 4898 39172 4900
rect 38892 4846 38894 4898
rect 38946 4846 39172 4898
rect 38892 4844 39172 4846
rect 38892 4834 38948 4844
rect 38892 4564 38948 4574
rect 38780 4562 38948 4564
rect 38780 4510 38894 4562
rect 38946 4510 38948 4562
rect 38780 4508 38948 4510
rect 38892 4498 38948 4508
rect 37996 4452 38052 4462
rect 37996 4338 38052 4396
rect 37996 4286 37998 4338
rect 38050 4286 38052 4338
rect 37996 4274 38052 4286
rect 38220 4450 38276 4462
rect 38220 4398 38222 4450
rect 38274 4398 38276 4450
rect 37212 3502 37214 3554
rect 37266 3502 37268 3554
rect 37212 3490 37268 3502
rect 37660 4228 37716 4238
rect 36428 3330 36484 3342
rect 36428 3278 36430 3330
rect 36482 3278 36484 3330
rect 36428 1652 36484 3278
rect 35644 1596 36484 1652
rect 36540 3332 36820 3388
rect 37548 3332 37604 3342
rect 35644 800 35700 1596
rect 36540 980 36596 3332
rect 36316 924 36596 980
rect 36988 3330 37604 3332
rect 36988 3278 37550 3330
rect 37602 3278 37604 3330
rect 36988 3276 37604 3278
rect 36316 800 36372 924
rect 36988 800 37044 3276
rect 37548 3266 37604 3276
rect 37660 800 37716 4172
rect 38220 3556 38276 4398
rect 38556 4338 38612 4350
rect 38556 4286 38558 4338
rect 38610 4286 38612 4338
rect 38556 4228 38612 4286
rect 38556 4162 38612 4172
rect 38220 3490 38276 3500
rect 39004 3668 39060 3678
rect 38444 3332 38500 3342
rect 38332 3330 38500 3332
rect 38332 3278 38446 3330
rect 38498 3278 38500 3330
rect 38332 3276 38500 3278
rect 38332 800 38388 3276
rect 38444 3266 38500 3276
rect 39004 800 39060 3612
rect 39116 3554 39172 4844
rect 39116 3502 39118 3554
rect 39170 3502 39172 3554
rect 39116 3490 39172 3502
rect 39564 4898 39620 4910
rect 39564 4846 39566 4898
rect 39618 4846 39620 4898
rect 39564 3444 39620 4846
rect 40684 4898 40740 4910
rect 40684 4846 40686 4898
rect 40738 4846 40740 4898
rect 39900 4452 39956 4462
rect 39564 3378 39620 3388
rect 39676 4450 39956 4452
rect 39676 4398 39902 4450
rect 39954 4398 39956 4450
rect 39676 4396 39956 4398
rect 39676 800 39732 4396
rect 39900 4386 39956 4396
rect 40236 3668 40292 3678
rect 40236 3574 40292 3612
rect 39788 3556 39844 3566
rect 39788 3462 39844 3500
rect 40684 3108 40740 4846
rect 40908 4562 40964 4956
rect 40908 4510 40910 4562
rect 40962 4510 40964 4562
rect 40908 4498 40964 4510
rect 41468 5010 41524 5022
rect 41468 4958 41470 5010
rect 41522 4958 41524 5010
rect 41468 4564 41524 4958
rect 41804 5010 41860 5852
rect 42252 5794 42308 5806
rect 42252 5742 42254 5794
rect 42306 5742 42308 5794
rect 41804 4958 41806 5010
rect 41858 4958 41860 5010
rect 41804 4946 41860 4958
rect 42140 5010 42196 5022
rect 42140 4958 42142 5010
rect 42194 4958 42196 5010
rect 41468 4498 41524 4508
rect 41580 4452 41636 4462
rect 41580 4358 41636 4396
rect 41132 4338 41188 4350
rect 41132 4286 41134 4338
rect 41186 4286 41188 4338
rect 41132 3444 41188 4286
rect 41804 4338 41860 4350
rect 41804 4286 41806 4338
rect 41858 4286 41860 4338
rect 41804 3780 41860 4286
rect 42140 4228 42196 4958
rect 42252 4900 42308 5742
rect 42476 5010 42532 8204
rect 42924 8194 42980 8204
rect 42588 7586 42644 7598
rect 42588 7534 42590 7586
rect 42642 7534 42644 7586
rect 42588 6804 42644 7534
rect 42924 7476 42980 7486
rect 42588 6738 42644 6748
rect 42812 7474 42980 7476
rect 42812 7422 42926 7474
rect 42978 7422 42980 7474
rect 42812 7420 42980 7422
rect 42476 4958 42478 5010
rect 42530 4958 42532 5010
rect 42476 4946 42532 4958
rect 42700 5794 42756 5806
rect 42700 5742 42702 5794
rect 42754 5742 42756 5794
rect 42252 4834 42308 4844
rect 42140 4162 42196 4172
rect 42364 4450 42420 4462
rect 42364 4398 42366 4450
rect 42418 4398 42420 4450
rect 42364 4116 42420 4398
rect 42700 4340 42756 5742
rect 42812 5010 42868 7420
rect 42924 7410 42980 7420
rect 43148 6692 43204 6702
rect 43148 6690 43540 6692
rect 43148 6638 43150 6690
rect 43202 6638 43540 6690
rect 43148 6636 43540 6638
rect 43148 6626 43204 6636
rect 42924 5908 42980 5918
rect 42924 5814 42980 5852
rect 42812 4958 42814 5010
rect 42866 4958 42868 5010
rect 42812 4946 42868 4958
rect 43148 5010 43204 5022
rect 43148 4958 43150 5010
rect 43202 4958 43204 5010
rect 43036 4788 43092 4798
rect 42924 4732 43036 4788
rect 42812 4564 42868 4574
rect 42924 4564 42980 4732
rect 43036 4722 43092 4732
rect 43148 4676 43204 4958
rect 43484 5010 43540 6636
rect 43820 5122 43876 9102
rect 44156 9042 44212 9054
rect 44156 8990 44158 9042
rect 44210 8990 44212 9042
rect 44156 8820 44212 8990
rect 44156 8754 44212 8764
rect 44044 8148 44100 8158
rect 44044 8054 44100 8092
rect 44044 7476 44100 7486
rect 44044 7382 44100 7420
rect 44044 6578 44100 6590
rect 44044 6526 44046 6578
rect 44098 6526 44100 6578
rect 44044 6132 44100 6526
rect 44044 6066 44100 6076
rect 44044 5794 44100 5806
rect 44044 5742 44046 5794
rect 44098 5742 44100 5794
rect 44044 5460 44100 5742
rect 44044 5394 44100 5404
rect 43820 5070 43822 5122
rect 43874 5070 43876 5122
rect 43820 5058 43876 5070
rect 43484 4958 43486 5010
rect 43538 4958 43540 5010
rect 43484 4946 43540 4958
rect 44156 4900 44212 4910
rect 43148 4610 43204 4620
rect 43820 4676 43876 4686
rect 42812 4562 42980 4564
rect 42812 4510 42814 4562
rect 42866 4510 42980 4562
rect 42812 4508 42980 4510
rect 43036 4564 43092 4574
rect 42812 4498 42868 4508
rect 43036 4452 43092 4508
rect 43820 4562 43876 4620
rect 43820 4510 43822 4562
rect 43874 4510 43876 4562
rect 43820 4498 43876 4510
rect 43148 4452 43204 4462
rect 43036 4450 43204 4452
rect 43036 4398 43150 4450
rect 43202 4398 43204 4450
rect 43036 4396 43204 4398
rect 43148 4386 43204 4396
rect 42700 4274 42756 4284
rect 43372 4338 43428 4350
rect 43372 4286 43374 4338
rect 43426 4286 43428 4338
rect 42364 4050 42420 4060
rect 41580 3724 41860 3780
rect 40908 3388 41188 3444
rect 41244 3444 41300 3454
rect 41580 3444 41636 3724
rect 42252 3668 42308 3678
rect 41244 3442 41636 3444
rect 41244 3390 41246 3442
rect 41298 3390 41636 3442
rect 41244 3388 41636 3390
rect 41692 3666 42308 3668
rect 41692 3614 42254 3666
rect 42306 3614 42308 3666
rect 41692 3612 42308 3614
rect 40908 3108 40964 3388
rect 41244 3332 41300 3388
rect 40348 3052 40964 3108
rect 41020 3276 41300 3332
rect 40348 800 40404 3052
rect 41020 800 41076 3276
rect 41692 800 41748 3612
rect 42252 3602 42308 3612
rect 41804 3444 41860 3454
rect 41804 3350 41860 3388
rect 43148 3444 43204 3454
rect 43372 3444 43428 4286
rect 44044 4340 44100 4350
rect 44044 4246 44100 4284
rect 43148 3442 43428 3444
rect 43148 3390 43150 3442
rect 43202 3390 43428 3442
rect 43148 3388 43428 3390
rect 43820 4228 43876 4238
rect 43820 3442 43876 4172
rect 43820 3390 43822 3442
rect 43874 3390 43876 3442
rect 43148 2772 43204 3388
rect 43820 3378 43876 3390
rect 44156 3444 44212 4844
rect 44156 3350 44212 3388
rect 44380 4340 44436 4350
rect 43148 2706 43204 2716
rect 44380 2100 44436 4284
rect 44380 2034 44436 2044
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
rect 40320 0 40432 800
rect 40992 0 41104 800
rect 41664 0 41776 800
rect 42336 0 42448 800
rect 43008 0 43120 800
rect 43680 0 43792 800
rect 44352 0 44464 800
rect 45024 0 45136 800
rect 45696 0 45808 800
<< via2 >>
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 14588 41970 14644 41972
rect 14588 41918 14590 41970
rect 14590 41918 14642 41970
rect 14642 41918 14644 41970
rect 14588 41916 14644 41918
rect 14476 40460 14532 40516
rect 15260 41970 15316 41972
rect 15260 41918 15262 41970
rect 15262 41918 15314 41970
rect 15314 41918 15316 41970
rect 15260 41916 15316 41918
rect 15148 41132 15204 41188
rect 16380 41916 16436 41972
rect 16940 41132 16996 41188
rect 17388 41916 17444 41972
rect 18172 41356 18228 41412
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19292 41356 19348 41412
rect 18844 41132 18900 41188
rect 15484 40514 15540 40516
rect 15484 40462 15486 40514
rect 15486 40462 15538 40514
rect 15538 40462 15540 40514
rect 15484 40460 15540 40462
rect 20188 41020 20244 41076
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 21644 35922 21700 35924
rect 21644 35870 21646 35922
rect 21646 35870 21698 35922
rect 21698 35870 21700 35922
rect 21644 35868 21700 35870
rect 41916 45724 41972 45780
rect 22428 35868 22484 35924
rect 24892 41298 24948 41300
rect 24892 41246 24894 41298
rect 24894 41246 24946 41298
rect 24946 41246 24948 41298
rect 24892 41244 24948 41246
rect 26236 41916 26292 41972
rect 26012 41244 26068 41300
rect 26908 41916 26964 41972
rect 27916 41970 27972 41972
rect 27916 41918 27918 41970
rect 27918 41918 27970 41970
rect 27970 41918 27972 41970
rect 27916 41916 27972 41918
rect 26236 38556 26292 38612
rect 26460 35922 26516 35924
rect 26460 35870 26462 35922
rect 26462 35870 26514 35922
rect 26514 35870 26516 35922
rect 26460 35868 26516 35870
rect 28588 41970 28644 41972
rect 28588 41918 28590 41970
rect 28590 41918 28642 41970
rect 28642 41918 28644 41970
rect 28588 41916 28644 41918
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 36316 40460 36372 40516
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 39004 41916 39060 41972
rect 38220 40962 38276 40964
rect 38220 40910 38222 40962
rect 38222 40910 38274 40962
rect 38274 40910 38276 40962
rect 38220 40908 38276 40910
rect 39564 40572 39620 40628
rect 38780 40514 38836 40516
rect 38780 40462 38782 40514
rect 38782 40462 38834 40514
rect 38834 40462 38836 40514
rect 38780 40460 38836 40462
rect 40348 41916 40404 41972
rect 39788 40908 39844 40964
rect 40124 40796 40180 40852
rect 37548 39564 37604 39620
rect 39116 39618 39172 39620
rect 39116 39566 39118 39618
rect 39118 39566 39170 39618
rect 39170 39566 39172 39618
rect 39116 39564 39172 39566
rect 39900 39618 39956 39620
rect 39900 39566 39902 39618
rect 39902 39566 39954 39618
rect 39954 39566 39956 39618
rect 39900 39564 39956 39566
rect 40348 39676 40404 39732
rect 40908 39564 40964 39620
rect 41692 40908 41748 40964
rect 44268 45052 44324 45108
rect 43932 44380 43988 44436
rect 43708 43708 43764 43764
rect 43484 42364 43540 42420
rect 43148 41858 43204 41860
rect 43148 41806 43150 41858
rect 43150 41806 43202 41858
rect 43202 41806 43204 41858
rect 43148 41804 43204 41806
rect 41804 40796 41860 40852
rect 41692 40402 41748 40404
rect 41692 40350 41694 40402
rect 41694 40350 41746 40402
rect 41746 40350 41748 40402
rect 41692 40348 41748 40350
rect 41916 40514 41972 40516
rect 41916 40462 41918 40514
rect 41918 40462 41970 40514
rect 41970 40462 41972 40514
rect 41916 40460 41972 40462
rect 42252 39340 42308 39396
rect 42924 40514 42980 40516
rect 42924 40462 42926 40514
rect 42926 40462 42978 40514
rect 42978 40462 42980 40514
rect 42924 40460 42980 40462
rect 43820 40572 43876 40628
rect 44156 41804 44212 41860
rect 44044 41692 44100 41748
rect 43484 40348 43540 40404
rect 42812 39506 42868 39508
rect 42812 39454 42814 39506
rect 42814 39454 42866 39506
rect 42866 39454 42868 39506
rect 42812 39452 42868 39454
rect 43372 39394 43428 39396
rect 43372 39342 43374 39394
rect 43374 39342 43426 39394
rect 43426 39342 43428 39394
rect 43372 39340 43428 39342
rect 42364 39058 42420 39060
rect 42364 39006 42366 39058
rect 42366 39006 42418 39058
rect 42418 39006 42420 39058
rect 42364 39004 42420 39006
rect 28364 38556 28420 38612
rect 42812 38556 42868 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 43148 38162 43204 38164
rect 43148 38110 43150 38162
rect 43150 38110 43202 38162
rect 43202 38110 43204 38162
rect 43148 38108 43204 38110
rect 43484 37826 43540 37828
rect 43484 37774 43486 37826
rect 43486 37774 43538 37826
rect 43538 37774 43540 37826
rect 43484 37772 43540 37774
rect 43820 39452 43876 39508
rect 44380 43036 44436 43092
rect 44044 38108 44100 38164
rect 44492 41804 44548 41860
rect 44492 41020 44548 41076
rect 44380 38108 44436 38164
rect 44156 36988 44212 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 43708 36370 43764 36372
rect 43708 36318 43710 36370
rect 43710 36318 43762 36370
rect 43762 36318 43764 36370
rect 43708 36316 43764 36318
rect 27132 35868 27188 35924
rect 44156 35810 44212 35812
rect 44156 35758 44158 35810
rect 44158 35758 44210 35810
rect 44210 35758 44212 35810
rect 44156 35756 44212 35758
rect 44268 35644 44324 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1820 28588 1876 28644
rect 3612 28924 3668 28980
rect 3052 28700 3108 28756
rect 3052 27692 3108 27748
rect 1708 27580 1764 27636
rect 2828 26124 2884 26180
rect 3052 23826 3108 23828
rect 3052 23774 3054 23826
rect 3054 23774 3106 23826
rect 3106 23774 3108 23826
rect 3052 23772 3108 23774
rect 3052 22258 3108 22260
rect 3052 22206 3054 22258
rect 3054 22206 3106 22258
rect 3106 22206 3108 22258
rect 3052 22204 3108 22206
rect 3948 28476 4004 28532
rect 3836 27804 3892 27860
rect 3724 26178 3780 26180
rect 3724 26126 3726 26178
rect 3726 26126 3778 26178
rect 3778 26126 3780 26178
rect 3724 26124 3780 26126
rect 3724 25564 3780 25620
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4956 28754 5012 28756
rect 4956 28702 4958 28754
rect 4958 28702 5010 28754
rect 5010 28702 5012 28754
rect 4956 28700 5012 28702
rect 4844 28642 4900 28644
rect 4844 28590 4846 28642
rect 4846 28590 4898 28642
rect 4898 28590 4900 28642
rect 4844 28588 4900 28590
rect 4284 27692 4340 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3948 27020 4004 27076
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4508 25618 4564 25620
rect 4508 25566 4510 25618
rect 4510 25566 4562 25618
rect 4562 25566 4564 25618
rect 4508 25564 4564 25566
rect 11228 30322 11284 30324
rect 11228 30270 11230 30322
rect 11230 30270 11282 30322
rect 11282 30270 11284 30322
rect 11228 30268 11284 30270
rect 5292 30044 5348 30100
rect 7644 30098 7700 30100
rect 7644 30046 7646 30098
rect 7646 30046 7698 30098
rect 7698 30046 7700 30098
rect 7644 30044 7700 30046
rect 6188 29260 6244 29316
rect 5740 28642 5796 28644
rect 5740 28590 5742 28642
rect 5742 28590 5794 28642
rect 5794 28590 5796 28642
rect 5740 28588 5796 28590
rect 5516 27916 5572 27972
rect 5292 27858 5348 27860
rect 5292 27806 5294 27858
rect 5294 27806 5346 27858
rect 5346 27806 5348 27858
rect 5292 27804 5348 27806
rect 5740 27858 5796 27860
rect 5740 27806 5742 27858
rect 5742 27806 5794 27858
rect 5794 27806 5796 27858
rect 5740 27804 5796 27806
rect 5516 27074 5572 27076
rect 5516 27022 5518 27074
rect 5518 27022 5570 27074
rect 5570 27022 5572 27074
rect 5516 27020 5572 27022
rect 7532 29314 7588 29316
rect 7532 29262 7534 29314
rect 7534 29262 7586 29314
rect 7586 29262 7588 29314
rect 7532 29260 7588 29262
rect 6748 28642 6804 28644
rect 6748 28590 6750 28642
rect 6750 28590 6802 28642
rect 6802 28590 6804 28642
rect 6748 28588 6804 28590
rect 7420 28642 7476 28644
rect 7420 28590 7422 28642
rect 7422 28590 7474 28642
rect 7474 28590 7476 28642
rect 7420 28588 7476 28590
rect 6636 27970 6692 27972
rect 6636 27918 6638 27970
rect 6638 27918 6690 27970
rect 6690 27918 6692 27970
rect 6636 27916 6692 27918
rect 6300 27020 6356 27076
rect 7868 27804 7924 27860
rect 7644 27692 7700 27748
rect 8540 27692 8596 27748
rect 9996 29372 10052 29428
rect 9324 27804 9380 27860
rect 9884 27746 9940 27748
rect 9884 27694 9886 27746
rect 9886 27694 9938 27746
rect 9938 27694 9940 27746
rect 9884 27692 9940 27694
rect 9548 27356 9604 27412
rect 7420 26012 7476 26068
rect 8876 26124 8932 26180
rect 8316 26012 8372 26068
rect 8652 26012 8708 26068
rect 7420 25564 7476 25620
rect 11452 29372 11508 29428
rect 11564 31612 11620 31668
rect 12460 31666 12516 31668
rect 12460 31614 12462 31666
rect 12462 31614 12514 31666
rect 12514 31614 12516 31666
rect 12460 31612 12516 31614
rect 16604 31612 16660 31668
rect 14140 31106 14196 31108
rect 14140 31054 14142 31106
rect 14142 31054 14194 31106
rect 14194 31054 14196 31106
rect 14140 31052 14196 31054
rect 12124 30268 12180 30324
rect 10780 27692 10836 27748
rect 10780 27020 10836 27076
rect 9772 26796 9828 26852
rect 11564 26796 11620 26852
rect 11900 27020 11956 27076
rect 11004 26124 11060 26180
rect 6972 25228 7028 25284
rect 9324 25282 9380 25284
rect 9324 25230 9326 25282
rect 9326 25230 9378 25282
rect 9378 25230 9380 25282
rect 9324 25228 9380 25230
rect 10108 24892 10164 24948
rect 9436 24780 9492 24836
rect 7980 24668 8036 24724
rect 10220 24780 10276 24836
rect 10108 24722 10164 24724
rect 10108 24670 10110 24722
rect 10110 24670 10162 24722
rect 10162 24670 10164 24722
rect 10108 24668 10164 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6748 24108 6804 24164
rect 4060 24050 4116 24052
rect 4060 23998 4062 24050
rect 4062 23998 4114 24050
rect 4114 23998 4116 24050
rect 4060 23996 4116 23998
rect 9996 23938 10052 23940
rect 9996 23886 9998 23938
rect 9998 23886 10050 23938
rect 10050 23886 10052 23938
rect 9996 23884 10052 23886
rect 12236 26962 12292 26964
rect 12236 26910 12238 26962
rect 12238 26910 12290 26962
rect 12290 26910 12292 26962
rect 12236 26908 12292 26910
rect 12796 26796 12852 26852
rect 12572 26124 12628 26180
rect 14476 29372 14532 29428
rect 17388 31666 17444 31668
rect 17388 31614 17390 31666
rect 17390 31614 17442 31666
rect 17442 31614 17444 31666
rect 17388 31612 17444 31614
rect 17164 31052 17220 31108
rect 16380 28476 16436 28532
rect 13916 27074 13972 27076
rect 13916 27022 13918 27074
rect 13918 27022 13970 27074
rect 13970 27022 13972 27074
rect 13916 27020 13972 27022
rect 14812 26962 14868 26964
rect 14812 26910 14814 26962
rect 14814 26910 14866 26962
rect 14866 26910 14868 26962
rect 14812 26908 14868 26910
rect 12908 26012 12964 26068
rect 14812 26290 14868 26292
rect 14812 26238 14814 26290
rect 14814 26238 14866 26290
rect 14866 26238 14868 26290
rect 14812 26236 14868 26238
rect 15148 26178 15204 26180
rect 15148 26126 15150 26178
rect 15150 26126 15202 26178
rect 15202 26126 15204 26178
rect 15148 26124 15204 26126
rect 16828 27746 16884 27748
rect 16828 27694 16830 27746
rect 16830 27694 16882 27746
rect 16882 27694 16884 27746
rect 16828 27692 16884 27694
rect 15596 26236 15652 26292
rect 14028 25676 14084 25732
rect 13356 25452 13412 25508
rect 13244 25340 13300 25396
rect 11004 24050 11060 24052
rect 11004 23998 11006 24050
rect 11006 23998 11058 24050
rect 11058 23998 11060 24050
rect 11004 23996 11060 23998
rect 11900 24162 11956 24164
rect 11900 24110 11902 24162
rect 11902 24110 11954 24162
rect 11954 24110 11956 24162
rect 11900 24108 11956 24110
rect 4060 23266 4116 23268
rect 4060 23214 4062 23266
rect 4062 23214 4114 23266
rect 4114 23214 4116 23266
rect 4060 23212 4116 23214
rect 5180 23042 5236 23044
rect 5180 22990 5182 23042
rect 5182 22990 5234 23042
rect 5234 22990 5236 23042
rect 5180 22988 5236 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4060 22482 4116 22484
rect 4060 22430 4062 22482
rect 4062 22430 4114 22482
rect 4114 22430 4116 22482
rect 4060 22428 4116 22430
rect 3612 22092 3668 22148
rect 4060 21868 4116 21924
rect 2044 19122 2100 19124
rect 2044 19070 2046 19122
rect 2046 19070 2098 19122
rect 2098 19070 2100 19122
rect 2044 19068 2100 19070
rect 1708 18844 1764 18900
rect 3052 21308 3108 21364
rect 6076 21868 6132 21924
rect 9212 23772 9268 23828
rect 6972 23324 7028 23380
rect 6860 22204 6916 22260
rect 4732 21586 4788 21588
rect 4732 21534 4734 21586
rect 4734 21534 4786 21586
rect 4786 21534 4788 21586
rect 4732 21532 4788 21534
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 6860 21532 6916 21588
rect 5404 21362 5460 21364
rect 5404 21310 5406 21362
rect 5406 21310 5458 21362
rect 5458 21310 5460 21362
rect 5404 21308 5460 21310
rect 5068 20188 5124 20244
rect 3276 20130 3332 20132
rect 3276 20078 3278 20130
rect 3278 20078 3330 20130
rect 3330 20078 3332 20130
rect 3276 20076 3332 20078
rect 5964 20076 6020 20132
rect 1596 16658 1652 16660
rect 1596 16606 1598 16658
rect 1598 16606 1650 16658
rect 1650 16606 1652 16658
rect 1596 16604 1652 16606
rect 1932 16098 1988 16100
rect 1932 16046 1934 16098
rect 1934 16046 1986 16098
rect 1986 16046 1988 16098
rect 1932 16044 1988 16046
rect 1820 15932 1876 15988
rect 2268 16828 2324 16884
rect 2380 16604 2436 16660
rect 3052 18396 3108 18452
rect 3052 18172 3108 18228
rect 3948 19180 4004 19236
rect 3948 17778 4004 17780
rect 3948 17726 3950 17778
rect 3950 17726 4002 17778
rect 4002 17726 4004 17778
rect 3948 17724 4004 17726
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 6076 19292 6132 19348
rect 5516 18396 5572 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5740 18226 5796 18228
rect 5740 18174 5742 18226
rect 5742 18174 5794 18226
rect 5794 18174 5796 18226
rect 5740 18172 5796 18174
rect 4284 17724 4340 17780
rect 4060 16828 4116 16884
rect 4732 16940 4788 16996
rect 5068 16882 5124 16884
rect 5068 16830 5070 16882
rect 5070 16830 5122 16882
rect 5122 16830 5124 16882
rect 5068 16828 5124 16830
rect 6300 17442 6356 17444
rect 6300 17390 6302 17442
rect 6302 17390 6354 17442
rect 6354 17390 6356 17442
rect 6300 17388 6356 17390
rect 2716 16492 2772 16548
rect 3500 16492 3556 16548
rect 2940 16156 2996 16212
rect 2716 15986 2772 15988
rect 2716 15934 2718 15986
rect 2718 15934 2770 15986
rect 2770 15934 2772 15986
rect 2716 15932 2772 15934
rect 2716 14140 2772 14196
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 3836 16210 3892 16212
rect 3836 16158 3838 16210
rect 3838 16158 3890 16210
rect 3890 16158 3892 16210
rect 3836 16156 3892 16158
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3612 14140 3668 14196
rect 5740 15090 5796 15092
rect 5740 15038 5742 15090
rect 5742 15038 5794 15090
rect 5794 15038 5796 15090
rect 5740 15036 5796 15038
rect 6188 16044 6244 16100
rect 6300 15148 6356 15204
rect 7980 22876 8036 22932
rect 9436 23266 9492 23268
rect 9436 23214 9438 23266
rect 9438 23214 9490 23266
rect 9490 23214 9492 23266
rect 9436 23212 9492 23214
rect 9884 22988 9940 23044
rect 8540 22428 8596 22484
rect 7980 20802 8036 20804
rect 7980 20750 7982 20802
rect 7982 20750 8034 20802
rect 8034 20750 8036 20802
rect 7980 20748 8036 20750
rect 7420 20690 7476 20692
rect 7420 20638 7422 20690
rect 7422 20638 7474 20690
rect 7474 20638 7476 20690
rect 7420 20636 7476 20638
rect 7196 20188 7252 20244
rect 6972 19346 7028 19348
rect 6972 19294 6974 19346
rect 6974 19294 7026 19346
rect 7026 19294 7028 19346
rect 6972 19292 7028 19294
rect 7980 20188 8036 20244
rect 8316 19906 8372 19908
rect 8316 19854 8318 19906
rect 8318 19854 8370 19906
rect 8370 19854 8372 19906
rect 8316 19852 8372 19854
rect 7980 19292 8036 19348
rect 7756 19234 7812 19236
rect 7756 19182 7758 19234
rect 7758 19182 7810 19234
rect 7810 19182 7812 19234
rect 7756 19180 7812 19182
rect 11340 21980 11396 22036
rect 10220 21756 10276 21812
rect 9100 20748 9156 20804
rect 8988 20636 9044 20692
rect 9996 21644 10052 21700
rect 9996 20748 10052 20804
rect 12572 23996 12628 24052
rect 12012 23100 12068 23156
rect 11788 21644 11844 21700
rect 11900 21756 11956 21812
rect 11004 20972 11060 21028
rect 12124 21644 12180 21700
rect 12124 20860 12180 20916
rect 9996 20524 10052 20580
rect 11676 20578 11732 20580
rect 11676 20526 11678 20578
rect 11678 20526 11730 20578
rect 11730 20526 11732 20578
rect 11676 20524 11732 20526
rect 10108 19852 10164 19908
rect 11228 19180 11284 19236
rect 7196 16940 7252 16996
rect 8428 16156 8484 16212
rect 7420 16044 7476 16100
rect 8876 16882 8932 16884
rect 8876 16830 8878 16882
rect 8878 16830 8930 16882
rect 8930 16830 8932 16882
rect 8876 16828 8932 16830
rect 9436 16882 9492 16884
rect 9436 16830 9438 16882
rect 9438 16830 9490 16882
rect 9490 16830 9492 16882
rect 9436 16828 9492 16830
rect 8540 16044 8596 16100
rect 13580 25394 13636 25396
rect 13580 25342 13582 25394
rect 13582 25342 13634 25394
rect 13634 25342 13636 25394
rect 13580 25340 13636 25342
rect 13468 24892 13524 24948
rect 14924 25618 14980 25620
rect 14924 25566 14926 25618
rect 14926 25566 14978 25618
rect 14978 25566 14980 25618
rect 14924 25564 14980 25566
rect 15820 26178 15876 26180
rect 15820 26126 15822 26178
rect 15822 26126 15874 26178
rect 15874 26126 15876 26178
rect 15820 26124 15876 26126
rect 13692 23996 13748 24052
rect 15484 23996 15540 24052
rect 13020 22988 13076 23044
rect 13020 21868 13076 21924
rect 12796 20860 12852 20916
rect 12460 19964 12516 20020
rect 13804 23154 13860 23156
rect 13804 23102 13806 23154
rect 13806 23102 13858 23154
rect 13858 23102 13860 23154
rect 13804 23100 13860 23102
rect 13580 22988 13636 23044
rect 13804 22876 13860 22932
rect 14924 22540 14980 22596
rect 15820 22988 15876 23044
rect 14364 22258 14420 22260
rect 14364 22206 14366 22258
rect 14366 22206 14418 22258
rect 14418 22206 14420 22258
rect 14364 22204 14420 22206
rect 13916 21980 13972 22036
rect 13356 21026 13412 21028
rect 13356 20974 13358 21026
rect 13358 20974 13410 21026
rect 13410 20974 13412 21026
rect 13356 20972 13412 20974
rect 14364 21868 14420 21924
rect 13244 19964 13300 20020
rect 12236 19180 12292 19236
rect 11452 19122 11508 19124
rect 11452 19070 11454 19122
rect 11454 19070 11506 19122
rect 11506 19070 11508 19122
rect 11452 19068 11508 19070
rect 10892 16940 10948 16996
rect 11116 17388 11172 17444
rect 9996 15260 10052 15316
rect 8428 15036 8484 15092
rect 4956 13468 5012 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5964 13522 6020 13524
rect 5964 13470 5966 13522
rect 5966 13470 6018 13522
rect 6018 13470 6020 13522
rect 5964 13468 6020 13470
rect 10668 16156 10724 16212
rect 10220 15426 10276 15428
rect 10220 15374 10222 15426
rect 10222 15374 10274 15426
rect 10274 15374 10276 15426
rect 10220 15372 10276 15374
rect 11340 16828 11396 16884
rect 12572 19068 12628 19124
rect 12348 16940 12404 16996
rect 11452 15820 11508 15876
rect 12124 15874 12180 15876
rect 12124 15822 12126 15874
rect 12126 15822 12178 15874
rect 12178 15822 12180 15874
rect 12124 15820 12180 15822
rect 11452 15426 11508 15428
rect 11452 15374 11454 15426
rect 11454 15374 11506 15426
rect 11506 15374 11508 15426
rect 11452 15372 11508 15374
rect 11564 15260 11620 15316
rect 10108 13020 10164 13076
rect 13468 19122 13524 19124
rect 13468 19070 13470 19122
rect 13470 19070 13522 19122
rect 13522 19070 13524 19122
rect 13468 19068 13524 19070
rect 13804 19122 13860 19124
rect 13804 19070 13806 19122
rect 13806 19070 13858 19122
rect 13858 19070 13860 19122
rect 13804 19068 13860 19070
rect 12684 16828 12740 16884
rect 14140 18284 14196 18340
rect 12908 16044 12964 16100
rect 13244 16882 13300 16884
rect 13244 16830 13246 16882
rect 13246 16830 13298 16882
rect 13298 16830 13300 16882
rect 13244 16828 13300 16830
rect 13132 16658 13188 16660
rect 13132 16606 13134 16658
rect 13134 16606 13186 16658
rect 13186 16606 13188 16658
rect 13132 16604 13188 16606
rect 13020 15820 13076 15876
rect 12460 15708 12516 15764
rect 13916 16940 13972 16996
rect 14140 16604 14196 16660
rect 12460 14588 12516 14644
rect 14028 14642 14084 14644
rect 14028 14590 14030 14642
rect 14030 14590 14082 14642
rect 14082 14590 14084 14642
rect 14028 14588 14084 14590
rect 11676 13580 11732 13636
rect 12460 13580 12516 13636
rect 14252 16044 14308 16100
rect 16268 25228 16324 25284
rect 16716 26124 16772 26180
rect 16492 25676 16548 25732
rect 17052 25564 17108 25620
rect 16828 25506 16884 25508
rect 16828 25454 16830 25506
rect 16830 25454 16882 25506
rect 16882 25454 16884 25506
rect 16828 25452 16884 25454
rect 16940 25228 16996 25284
rect 16940 24722 16996 24724
rect 16940 24670 16942 24722
rect 16942 24670 16994 24722
rect 16994 24670 16996 24722
rect 16940 24668 16996 24670
rect 17948 30098 18004 30100
rect 17948 30046 17950 30098
rect 17950 30046 18002 30098
rect 18002 30046 18004 30098
rect 17948 30044 18004 30046
rect 17500 29426 17556 29428
rect 17500 29374 17502 29426
rect 17502 29374 17554 29426
rect 17554 29374 17556 29426
rect 17500 29372 17556 29374
rect 20300 31836 20356 31892
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 22316 31890 22372 31892
rect 22316 31838 22318 31890
rect 22318 31838 22370 31890
rect 22370 31838 22372 31890
rect 22316 31836 22372 31838
rect 21532 31612 21588 31668
rect 20300 30380 20356 30436
rect 20188 30098 20244 30100
rect 20188 30046 20190 30098
rect 20190 30046 20242 30098
rect 20242 30046 20244 30098
rect 20188 30044 20244 30046
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 29372 19684 29428
rect 23548 31666 23604 31668
rect 23548 31614 23550 31666
rect 23550 31614 23602 31666
rect 23602 31614 23604 31666
rect 23548 31612 23604 31614
rect 44044 31666 44100 31668
rect 44044 31614 44046 31666
rect 44046 31614 44098 31666
rect 44098 31614 44100 31666
rect 44044 31612 44100 31614
rect 28028 31052 28084 31108
rect 27020 30828 27076 30884
rect 22540 30380 22596 30436
rect 21756 30268 21812 30324
rect 21644 29484 21700 29540
rect 19404 28642 19460 28644
rect 19404 28590 19406 28642
rect 19406 28590 19458 28642
rect 19458 28590 19460 28642
rect 19404 28588 19460 28590
rect 19180 28476 19236 28532
rect 17724 27746 17780 27748
rect 17724 27694 17726 27746
rect 17726 27694 17778 27746
rect 17778 27694 17780 27746
rect 17724 27692 17780 27694
rect 17724 27020 17780 27076
rect 19404 27186 19460 27188
rect 19404 27134 19406 27186
rect 19406 27134 19458 27186
rect 19458 27134 19460 27186
rect 19404 27132 19460 27134
rect 18844 26348 18900 26404
rect 19068 26908 19124 26964
rect 19180 26796 19236 26852
rect 21308 28476 21364 28532
rect 20524 28364 20580 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19852 27074 19908 27076
rect 19852 27022 19854 27074
rect 19854 27022 19906 27074
rect 19906 27022 19908 27074
rect 19852 27020 19908 27022
rect 19628 26962 19684 26964
rect 19628 26910 19630 26962
rect 19630 26910 19682 26962
rect 19682 26910 19684 26962
rect 19628 26908 19684 26910
rect 23100 30322 23156 30324
rect 23100 30270 23102 30322
rect 23102 30270 23154 30322
rect 23154 30270 23156 30322
rect 23100 30268 23156 30270
rect 24668 30268 24724 30324
rect 23324 30044 23380 30100
rect 24108 30098 24164 30100
rect 24108 30046 24110 30098
rect 24110 30046 24162 30098
rect 24162 30046 24164 30098
rect 24108 30044 24164 30046
rect 24220 29650 24276 29652
rect 24220 29598 24222 29650
rect 24222 29598 24274 29650
rect 24274 29598 24276 29650
rect 24220 29596 24276 29598
rect 22316 28754 22372 28756
rect 22316 28702 22318 28754
rect 22318 28702 22370 28754
rect 22370 28702 22372 28754
rect 22316 28700 22372 28702
rect 25900 30322 25956 30324
rect 25900 30270 25902 30322
rect 25902 30270 25954 30322
rect 25954 30270 25956 30322
rect 25900 30268 25956 30270
rect 24780 30044 24836 30100
rect 26908 30098 26964 30100
rect 26908 30046 26910 30098
rect 26910 30046 26962 30098
rect 26962 30046 26964 30098
rect 26908 30044 26964 30046
rect 25340 29650 25396 29652
rect 25340 29598 25342 29650
rect 25342 29598 25394 29650
rect 25394 29598 25396 29650
rect 25340 29596 25396 29598
rect 25228 29538 25284 29540
rect 25228 29486 25230 29538
rect 25230 29486 25282 29538
rect 25282 29486 25284 29538
rect 25228 29484 25284 29486
rect 25788 29260 25844 29316
rect 21644 28364 21700 28420
rect 20636 27074 20692 27076
rect 20636 27022 20638 27074
rect 20638 27022 20690 27074
rect 20690 27022 20692 27074
rect 20636 27020 20692 27022
rect 19516 26796 19572 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 26348 19684 26404
rect 19180 26124 19236 26180
rect 19628 26178 19684 26180
rect 19628 26126 19630 26178
rect 19630 26126 19682 26178
rect 19682 26126 19684 26178
rect 19628 26124 19684 26126
rect 17948 25228 18004 25284
rect 16380 24050 16436 24052
rect 16380 23998 16382 24050
rect 16382 23998 16434 24050
rect 16434 23998 16436 24050
rect 16380 23996 16436 23998
rect 17612 23996 17668 24052
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 25618 20356 25620
rect 20300 25566 20302 25618
rect 20302 25566 20354 25618
rect 20354 25566 20356 25618
rect 20300 25564 20356 25566
rect 20412 25228 20468 25284
rect 19628 24668 19684 24724
rect 18396 24444 18452 24500
rect 16940 23714 16996 23716
rect 16940 23662 16942 23714
rect 16942 23662 16994 23714
rect 16994 23662 16996 23714
rect 16940 23660 16996 23662
rect 16380 23436 16436 23492
rect 15932 22428 15988 22484
rect 18396 23660 18452 23716
rect 19404 24610 19460 24612
rect 19404 24558 19406 24610
rect 19406 24558 19458 24610
rect 19458 24558 19460 24610
rect 19404 24556 19460 24558
rect 20300 24722 20356 24724
rect 20300 24670 20302 24722
rect 20302 24670 20354 24722
rect 20354 24670 20356 24722
rect 20300 24668 20356 24670
rect 23436 27916 23492 27972
rect 23548 27132 23604 27188
rect 23996 28476 24052 28532
rect 23996 27970 24052 27972
rect 23996 27918 23998 27970
rect 23998 27918 24050 27970
rect 24050 27918 24052 27970
rect 23996 27916 24052 27918
rect 23884 27804 23940 27860
rect 25116 27858 25172 27860
rect 25116 27806 25118 27858
rect 25118 27806 25170 27858
rect 25170 27806 25172 27858
rect 25116 27804 25172 27806
rect 27804 29260 27860 29316
rect 27356 28924 27412 28980
rect 26236 27804 26292 27860
rect 22092 26796 22148 26852
rect 23212 26796 23268 26852
rect 21868 26290 21924 26292
rect 21868 26238 21870 26290
rect 21870 26238 21922 26290
rect 21922 26238 21924 26290
rect 21868 26236 21924 26238
rect 21756 25564 21812 25620
rect 23772 26178 23828 26180
rect 23772 26126 23774 26178
rect 23774 26126 23826 26178
rect 23826 26126 23828 26178
rect 23772 26124 23828 26126
rect 22876 25618 22932 25620
rect 22876 25566 22878 25618
rect 22878 25566 22930 25618
rect 22930 25566 22932 25618
rect 22876 25564 22932 25566
rect 23324 25340 23380 25396
rect 21532 24444 21588 24500
rect 23324 24050 23380 24052
rect 23324 23998 23326 24050
rect 23326 23998 23378 24050
rect 23378 23998 23380 24050
rect 23324 23996 23380 23998
rect 20860 23938 20916 23940
rect 20860 23886 20862 23938
rect 20862 23886 20914 23938
rect 20914 23886 20916 23938
rect 20860 23884 20916 23886
rect 19068 23436 19124 23492
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 16940 23378 16996 23380
rect 16940 23326 16942 23378
rect 16942 23326 16994 23378
rect 16994 23326 16996 23378
rect 16940 23324 16996 23326
rect 16828 22988 16884 23044
rect 16940 22540 16996 22596
rect 16604 22258 16660 22260
rect 16604 22206 16606 22258
rect 16606 22206 16658 22258
rect 16658 22206 16660 22258
rect 16604 22204 16660 22206
rect 17724 22428 17780 22484
rect 15372 21532 15428 21588
rect 15036 18956 15092 19012
rect 15372 16828 15428 16884
rect 15260 15820 15316 15876
rect 14700 15708 14756 15764
rect 14364 15148 14420 15204
rect 15036 15148 15092 15204
rect 16156 20018 16212 20020
rect 16156 19966 16158 20018
rect 16158 19966 16210 20018
rect 16210 19966 16212 20018
rect 16156 19964 16212 19966
rect 19068 23100 19124 23156
rect 20860 23154 20916 23156
rect 20860 23102 20862 23154
rect 20862 23102 20914 23154
rect 20914 23102 20916 23154
rect 20860 23100 20916 23102
rect 19740 22204 19796 22260
rect 20860 22146 20916 22148
rect 20860 22094 20862 22146
rect 20862 22094 20914 22146
rect 20914 22094 20916 22146
rect 20860 22092 20916 22094
rect 21420 22092 21476 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 18060 21756 18116 21812
rect 17500 20188 17556 20244
rect 15820 19068 15876 19124
rect 16716 19068 16772 19124
rect 16492 18338 16548 18340
rect 16492 18286 16494 18338
rect 16494 18286 16546 18338
rect 16546 18286 16548 18338
rect 16492 18284 16548 18286
rect 16828 18956 16884 19012
rect 17052 18396 17108 18452
rect 17612 18450 17668 18452
rect 17612 18398 17614 18450
rect 17614 18398 17666 18450
rect 17666 18398 17668 18450
rect 17612 18396 17668 18398
rect 15932 15202 15988 15204
rect 15932 15150 15934 15202
rect 15934 15150 15986 15202
rect 15986 15150 15988 15202
rect 15932 15148 15988 15150
rect 18844 21586 18900 21588
rect 18844 21534 18846 21586
rect 18846 21534 18898 21586
rect 18898 21534 18900 21586
rect 18844 21532 18900 21534
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19964 20188 20020 20244
rect 20188 20130 20244 20132
rect 20188 20078 20190 20130
rect 20190 20078 20242 20130
rect 20242 20078 20244 20130
rect 20188 20076 20244 20078
rect 20300 19404 20356 19460
rect 20300 19234 20356 19236
rect 20300 19182 20302 19234
rect 20302 19182 20354 19234
rect 20354 19182 20356 19234
rect 20300 19180 20356 19182
rect 20748 19010 20804 19012
rect 20748 18958 20750 19010
rect 20750 18958 20802 19010
rect 20802 18958 20804 19010
rect 20748 18956 20804 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 17052 16828 17108 16884
rect 16828 16716 16884 16772
rect 16380 15484 16436 15540
rect 16604 14700 16660 14756
rect 15260 13074 15316 13076
rect 15260 13022 15262 13074
rect 15262 13022 15314 13074
rect 15314 13022 15316 13074
rect 15260 13020 15316 13022
rect 16716 14364 16772 14420
rect 18060 17052 18116 17108
rect 17724 16268 17780 16324
rect 17836 16770 17892 16772
rect 17836 16718 17838 16770
rect 17838 16718 17890 16770
rect 17890 16718 17892 16770
rect 17836 16716 17892 16718
rect 17724 15484 17780 15540
rect 17836 15148 17892 15204
rect 18396 18396 18452 18452
rect 20524 17724 20580 17780
rect 18396 17388 18452 17444
rect 20188 17388 20244 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 17052 19908 17108
rect 18844 16380 18900 16436
rect 19516 16940 19572 16996
rect 18172 15820 18228 15876
rect 18844 16044 18900 16100
rect 18060 15202 18116 15204
rect 18060 15150 18062 15202
rect 18062 15150 18114 15202
rect 18114 15150 18116 15202
rect 18060 15148 18116 15150
rect 17948 14700 18004 14756
rect 19068 15820 19124 15876
rect 18508 14418 18564 14420
rect 18508 14366 18510 14418
rect 18510 14366 18562 14418
rect 18562 14366 18564 14418
rect 18508 14364 18564 14366
rect 19740 16098 19796 16100
rect 19740 16046 19742 16098
rect 19742 16046 19794 16098
rect 19794 16046 19796 16098
rect 19740 16044 19796 16046
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21980 21810 22036 21812
rect 21980 21758 21982 21810
rect 21982 21758 22034 21810
rect 22034 21758 22036 21810
rect 21980 21756 22036 21758
rect 22092 21532 22148 21588
rect 23100 22988 23156 23044
rect 22652 22876 22708 22932
rect 23212 22204 23268 22260
rect 21420 19404 21476 19460
rect 21084 18396 21140 18452
rect 22092 20076 22148 20132
rect 21644 19180 21700 19236
rect 22428 19234 22484 19236
rect 22428 19182 22430 19234
rect 22430 19182 22482 19234
rect 22482 19182 22484 19234
rect 22428 19180 22484 19182
rect 22540 18396 22596 18452
rect 21084 18226 21140 18228
rect 21084 18174 21086 18226
rect 21086 18174 21138 18226
rect 21138 18174 21140 18226
rect 21084 18172 21140 18174
rect 21420 17778 21476 17780
rect 21420 17726 21422 17778
rect 21422 17726 21474 17778
rect 21474 17726 21476 17778
rect 21420 17724 21476 17726
rect 20860 16828 20916 16884
rect 20972 16604 21028 16660
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21196 15932 21252 15988
rect 21308 16828 21364 16884
rect 21308 15484 21364 15540
rect 21420 16268 21476 16324
rect 24332 25564 24388 25620
rect 23884 25394 23940 25396
rect 23884 25342 23886 25394
rect 23886 25342 23938 25394
rect 23938 25342 23940 25394
rect 23884 25340 23940 25342
rect 28028 30098 28084 30100
rect 28028 30046 28030 30098
rect 28030 30046 28082 30098
rect 28082 30046 28084 30098
rect 28028 30044 28084 30046
rect 31500 31106 31556 31108
rect 31500 31054 31502 31106
rect 31502 31054 31554 31106
rect 31554 31054 31556 31106
rect 31500 31052 31556 31054
rect 32732 31052 32788 31108
rect 30492 30882 30548 30884
rect 30492 30830 30494 30882
rect 30494 30830 30546 30882
rect 30546 30830 30548 30882
rect 30492 30828 30548 30830
rect 29484 30098 29540 30100
rect 29484 30046 29486 30098
rect 29486 30046 29538 30098
rect 29538 30046 29540 30098
rect 29484 30044 29540 30046
rect 29708 29260 29764 29316
rect 28700 28924 28756 28980
rect 29596 29036 29652 29092
rect 26572 26962 26628 26964
rect 26572 26910 26574 26962
rect 26574 26910 26626 26962
rect 26626 26910 26628 26962
rect 26572 26908 26628 26910
rect 27580 26962 27636 26964
rect 27580 26910 27582 26962
rect 27582 26910 27634 26962
rect 27634 26910 27636 26962
rect 27580 26908 27636 26910
rect 27916 26962 27972 26964
rect 27916 26910 27918 26962
rect 27918 26910 27970 26962
rect 27970 26910 27972 26962
rect 27916 26908 27972 26910
rect 28588 27804 28644 27860
rect 29036 27858 29092 27860
rect 29036 27806 29038 27858
rect 29038 27806 29090 27858
rect 29090 27806 29092 27858
rect 29036 27804 29092 27806
rect 29932 29202 29988 29204
rect 29932 29150 29934 29202
rect 29934 29150 29986 29202
rect 29986 29150 29988 29202
rect 29932 29148 29988 29150
rect 31052 29036 31108 29092
rect 31164 28700 31220 28756
rect 26796 26178 26852 26180
rect 26796 26126 26798 26178
rect 26798 26126 26850 26178
rect 26850 26126 26852 26178
rect 26796 26124 26852 26126
rect 25676 25618 25732 25620
rect 25676 25566 25678 25618
rect 25678 25566 25730 25618
rect 25730 25566 25732 25618
rect 25676 25564 25732 25566
rect 24780 25340 24836 25396
rect 26908 25394 26964 25396
rect 26908 25342 26910 25394
rect 26910 25342 26962 25394
rect 26962 25342 26964 25394
rect 26908 25340 26964 25342
rect 27020 25116 27076 25172
rect 26460 24722 26516 24724
rect 26460 24670 26462 24722
rect 26462 24670 26514 24722
rect 26514 24670 26516 24722
rect 26460 24668 26516 24670
rect 23884 24610 23940 24612
rect 23884 24558 23886 24610
rect 23886 24558 23938 24610
rect 23938 24558 23940 24610
rect 23884 24556 23940 24558
rect 24444 24556 24500 24612
rect 24332 24444 24388 24500
rect 26236 24444 26292 24500
rect 25228 23996 25284 24052
rect 24556 23938 24612 23940
rect 24556 23886 24558 23938
rect 24558 23886 24610 23938
rect 24610 23886 24612 23938
rect 24556 23884 24612 23886
rect 25788 23884 25844 23940
rect 24556 23154 24612 23156
rect 24556 23102 24558 23154
rect 24558 23102 24610 23154
rect 24610 23102 24612 23154
rect 24556 23100 24612 23102
rect 25452 23100 25508 23156
rect 24332 23042 24388 23044
rect 24332 22990 24334 23042
rect 24334 22990 24386 23042
rect 24386 22990 24388 23042
rect 24332 22988 24388 22990
rect 23996 22930 24052 22932
rect 23996 22878 23998 22930
rect 23998 22878 24050 22930
rect 24050 22878 24052 22930
rect 23996 22876 24052 22878
rect 25340 21586 25396 21588
rect 25340 21534 25342 21586
rect 25342 21534 25394 21586
rect 25394 21534 25396 21586
rect 25340 21532 25396 21534
rect 23660 20748 23716 20804
rect 25340 20802 25396 20804
rect 25340 20750 25342 20802
rect 25342 20750 25394 20802
rect 25394 20750 25396 20802
rect 25340 20748 25396 20750
rect 23548 18956 23604 19012
rect 23884 18956 23940 19012
rect 23548 18172 23604 18228
rect 21756 16882 21812 16884
rect 21756 16830 21758 16882
rect 21758 16830 21810 16882
rect 21810 16830 21812 16882
rect 21756 16828 21812 16830
rect 22092 16380 22148 16436
rect 22316 15932 22372 15988
rect 21980 15148 22036 15204
rect 21644 14476 21700 14532
rect 21980 14476 22036 14532
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 22764 15484 22820 15540
rect 23436 15484 23492 15540
rect 23324 14028 23380 14084
rect 22988 13634 23044 13636
rect 22988 13582 22990 13634
rect 22990 13582 23042 13634
rect 23042 13582 23044 13634
rect 22988 13580 23044 13582
rect 23324 13356 23380 13412
rect 21756 11452 21812 11508
rect 24332 19852 24388 19908
rect 27132 24668 27188 24724
rect 26460 23884 26516 23940
rect 26236 23772 26292 23828
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 28812 25340 28868 25396
rect 31388 26908 31444 26964
rect 31388 26012 31444 26068
rect 29932 25004 29988 25060
rect 28588 24668 28644 24724
rect 29036 24668 29092 24724
rect 26460 21586 26516 21588
rect 26460 21534 26462 21586
rect 26462 21534 26514 21586
rect 26514 21534 26516 21586
rect 26460 21532 26516 21534
rect 27916 22482 27972 22484
rect 27916 22430 27918 22482
rect 27918 22430 27970 22482
rect 27970 22430 27972 22482
rect 27916 22428 27972 22430
rect 28252 23714 28308 23716
rect 28252 23662 28254 23714
rect 28254 23662 28306 23714
rect 28306 23662 28308 23714
rect 28252 23660 28308 23662
rect 28924 22988 28980 23044
rect 28476 22482 28532 22484
rect 28476 22430 28478 22482
rect 28478 22430 28530 22482
rect 28530 22430 28532 22482
rect 28476 22428 28532 22430
rect 27580 20860 27636 20916
rect 27020 20748 27076 20804
rect 24556 18956 24612 19012
rect 24556 18732 24612 18788
rect 26012 18956 26068 19012
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 25116 16658 25172 16660
rect 25116 16606 25118 16658
rect 25118 16606 25170 16658
rect 25170 16606 25172 16658
rect 25116 16604 25172 16606
rect 26012 18338 26068 18340
rect 26012 18286 26014 18338
rect 26014 18286 26066 18338
rect 26066 18286 26068 18338
rect 26012 18284 26068 18286
rect 26012 17890 26068 17892
rect 26012 17838 26014 17890
rect 26014 17838 26066 17890
rect 26066 17838 26068 17890
rect 26012 17836 26068 17838
rect 29372 22876 29428 22932
rect 31500 27580 31556 27636
rect 31052 24722 31108 24724
rect 31052 24670 31054 24722
rect 31054 24670 31106 24722
rect 31106 24670 31108 24722
rect 31052 24668 31108 24670
rect 31612 24668 31668 24724
rect 30156 24610 30212 24612
rect 30156 24558 30158 24610
rect 30158 24558 30210 24610
rect 30210 24558 30212 24610
rect 30156 24556 30212 24558
rect 30044 23884 30100 23940
rect 29932 23212 29988 23268
rect 29708 22540 29764 22596
rect 29820 22876 29876 22932
rect 29372 22428 29428 22484
rect 29484 21362 29540 21364
rect 29484 21310 29486 21362
rect 29486 21310 29538 21362
rect 29538 21310 29540 21362
rect 29484 21308 29540 21310
rect 31500 23266 31556 23268
rect 31500 23214 31502 23266
rect 31502 23214 31554 23266
rect 31554 23214 31556 23266
rect 31500 23212 31556 23214
rect 32620 30044 32676 30100
rect 34636 31106 34692 31108
rect 34636 31054 34638 31106
rect 34638 31054 34690 31106
rect 34690 31054 34692 31106
rect 34636 31052 34692 31054
rect 42476 31052 42532 31108
rect 43820 31106 43876 31108
rect 43820 31054 43822 31106
rect 43822 31054 43874 31106
rect 43874 31054 43876 31106
rect 43820 31052 43876 31054
rect 43596 30994 43652 30996
rect 43596 30942 43598 30994
rect 43598 30942 43650 30994
rect 43650 30942 43652 30994
rect 43596 30940 43652 30942
rect 44156 30994 44212 30996
rect 44156 30942 44158 30994
rect 44158 30942 44210 30994
rect 44210 30942 44212 30994
rect 44156 30940 44212 30942
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 33516 28812 33572 28868
rect 32956 27634 33012 27636
rect 32956 27582 32958 27634
rect 32958 27582 33010 27634
rect 33010 27582 33012 27634
rect 32956 27580 33012 27582
rect 34860 30098 34916 30100
rect 34860 30046 34862 30098
rect 34862 30046 34914 30098
rect 34914 30046 34916 30098
rect 34860 30044 34916 30046
rect 34188 29484 34244 29540
rect 34076 29314 34132 29316
rect 34076 29262 34078 29314
rect 34078 29262 34130 29314
rect 34130 29262 34132 29314
rect 34076 29260 34132 29262
rect 33852 28700 33908 28756
rect 33068 26908 33124 26964
rect 33404 26290 33460 26292
rect 33404 26238 33406 26290
rect 33406 26238 33458 26290
rect 33458 26238 33460 26290
rect 33404 26236 33460 26238
rect 32172 26124 32228 26180
rect 32172 25282 32228 25284
rect 32172 25230 32174 25282
rect 32174 25230 32226 25282
rect 32226 25230 32228 25282
rect 32172 25228 32228 25230
rect 32956 25116 33012 25172
rect 33628 25228 33684 25284
rect 32284 24722 32340 24724
rect 32284 24670 32286 24722
rect 32286 24670 32338 24722
rect 32338 24670 32340 24722
rect 32284 24668 32340 24670
rect 33516 25004 33572 25060
rect 32060 24556 32116 24612
rect 31948 23660 32004 23716
rect 30828 23042 30884 23044
rect 30828 22990 30830 23042
rect 30830 22990 30882 23042
rect 30882 22990 30884 23042
rect 30828 22988 30884 22990
rect 31164 23042 31220 23044
rect 31164 22990 31166 23042
rect 31166 22990 31218 23042
rect 31218 22990 31220 23042
rect 31164 22988 31220 22990
rect 31612 22988 31668 23044
rect 30492 22370 30548 22372
rect 30492 22318 30494 22370
rect 30494 22318 30546 22370
rect 30546 22318 30548 22370
rect 30492 22316 30548 22318
rect 30156 20914 30212 20916
rect 30156 20862 30158 20914
rect 30158 20862 30210 20914
rect 30210 20862 30212 20914
rect 30156 20860 30212 20862
rect 32844 23938 32900 23940
rect 32844 23886 32846 23938
rect 32846 23886 32898 23938
rect 32898 23886 32900 23938
rect 32844 23884 32900 23886
rect 35308 29148 35364 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34076 26908 34132 26964
rect 34860 26908 34916 26964
rect 33964 25394 34020 25396
rect 33964 25342 33966 25394
rect 33966 25342 34018 25394
rect 34018 25342 34020 25394
rect 33964 25340 34020 25342
rect 33852 25228 33908 25284
rect 34524 26796 34580 26852
rect 34076 23884 34132 23940
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 32508 23324 32564 23380
rect 32508 23042 32564 23044
rect 32508 22990 32510 23042
rect 32510 22990 32562 23042
rect 32562 22990 32564 23042
rect 32508 22988 32564 22990
rect 32956 23436 33012 23492
rect 33516 23378 33572 23380
rect 33516 23326 33518 23378
rect 33518 23326 33570 23378
rect 33570 23326 33572 23378
rect 33516 23324 33572 23326
rect 32732 22204 32788 22260
rect 33180 22540 33236 22596
rect 32508 21532 32564 21588
rect 30716 21474 30772 21476
rect 30716 21422 30718 21474
rect 30718 21422 30770 21474
rect 30770 21422 30772 21474
rect 30716 21420 30772 21422
rect 30604 20636 30660 20692
rect 31164 21308 31220 21364
rect 33516 22594 33572 22596
rect 33516 22542 33518 22594
rect 33518 22542 33570 22594
rect 33570 22542 33572 22594
rect 33516 22540 33572 22542
rect 34748 22482 34804 22484
rect 34748 22430 34750 22482
rect 34750 22430 34802 22482
rect 34802 22430 34804 22482
rect 34748 22428 34804 22430
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36540 30044 36596 30100
rect 37884 29538 37940 29540
rect 37884 29486 37886 29538
rect 37886 29486 37938 29538
rect 37938 29486 37940 29538
rect 37884 29484 37940 29486
rect 36876 28812 36932 28868
rect 37548 28700 37604 28756
rect 36316 26962 36372 26964
rect 36316 26910 36318 26962
rect 36318 26910 36370 26962
rect 36370 26910 36372 26962
rect 36316 26908 36372 26910
rect 35644 26236 35700 26292
rect 35644 25618 35700 25620
rect 35644 25566 35646 25618
rect 35646 25566 35698 25618
rect 35698 25566 35700 25618
rect 35644 25564 35700 25566
rect 35532 23996 35588 24052
rect 36988 25618 37044 25620
rect 36988 25566 36990 25618
rect 36990 25566 37042 25618
rect 37042 25566 37044 25618
rect 36988 25564 37044 25566
rect 37548 27692 37604 27748
rect 39004 30098 39060 30100
rect 39004 30046 39006 30098
rect 39006 30046 39058 30098
rect 39058 30046 39060 30098
rect 39004 30044 39060 30046
rect 41804 28754 41860 28756
rect 41804 28702 41806 28754
rect 41806 28702 41858 28754
rect 41858 28702 41860 28754
rect 41804 28700 41860 28702
rect 40796 28476 40852 28532
rect 37996 26796 38052 26852
rect 38220 27132 38276 27188
rect 37548 26402 37604 26404
rect 37548 26350 37550 26402
rect 37550 26350 37602 26402
rect 37602 26350 37604 26402
rect 37548 26348 37604 26350
rect 37436 26124 37492 26180
rect 37100 25282 37156 25284
rect 37100 25230 37102 25282
rect 37102 25230 37154 25282
rect 37154 25230 37156 25282
rect 37100 25228 37156 25230
rect 37436 24556 37492 24612
rect 37212 23996 37268 24052
rect 35644 23884 35700 23940
rect 36428 23884 36484 23940
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35756 22258 35812 22260
rect 35756 22206 35758 22258
rect 35758 22206 35810 22258
rect 35810 22206 35812 22258
rect 35756 22204 35812 22206
rect 33404 21586 33460 21588
rect 33404 21534 33406 21586
rect 33406 21534 33458 21586
rect 33458 21534 33460 21586
rect 33404 21532 33460 21534
rect 33852 21586 33908 21588
rect 33852 21534 33854 21586
rect 33854 21534 33906 21586
rect 33906 21534 33908 21586
rect 33852 21532 33908 21534
rect 33628 20748 33684 20804
rect 26460 18844 26516 18900
rect 26460 18450 26516 18452
rect 26460 18398 26462 18450
rect 26462 18398 26514 18450
rect 26514 18398 26516 18450
rect 26460 18396 26516 18398
rect 29596 19794 29652 19796
rect 29596 19742 29598 19794
rect 29598 19742 29650 19794
rect 29650 19742 29652 19794
rect 29596 19740 29652 19742
rect 27692 19010 27748 19012
rect 27692 18958 27694 19010
rect 27694 18958 27746 19010
rect 27746 18958 27748 19010
rect 27692 18956 27748 18958
rect 27356 17948 27412 18004
rect 26348 16940 26404 16996
rect 25900 16156 25956 16212
rect 25340 15538 25396 15540
rect 25340 15486 25342 15538
rect 25342 15486 25394 15538
rect 25394 15486 25396 15538
rect 25340 15484 25396 15486
rect 24220 15372 24276 15428
rect 25788 15426 25844 15428
rect 25788 15374 25790 15426
rect 25790 15374 25842 15426
rect 25842 15374 25844 15426
rect 25788 15372 25844 15374
rect 26124 15426 26180 15428
rect 26124 15374 26126 15426
rect 26126 15374 26178 15426
rect 26178 15374 26180 15426
rect 26124 15372 26180 15374
rect 26348 15874 26404 15876
rect 26348 15822 26350 15874
rect 26350 15822 26402 15874
rect 26402 15822 26404 15874
rect 26348 15820 26404 15822
rect 26348 15148 26404 15204
rect 24108 13580 24164 13636
rect 24780 13580 24836 13636
rect 26124 14028 26180 14084
rect 25676 12012 25732 12068
rect 27804 16210 27860 16212
rect 27804 16158 27806 16210
rect 27806 16158 27858 16210
rect 27858 16158 27860 16210
rect 27804 16156 27860 16158
rect 26684 15932 26740 15988
rect 27468 15986 27524 15988
rect 27468 15934 27470 15986
rect 27470 15934 27522 15986
rect 27522 15934 27524 15986
rect 27468 15932 27524 15934
rect 28364 17500 28420 17556
rect 28588 18956 28644 19012
rect 28364 16940 28420 16996
rect 28252 16882 28308 16884
rect 28252 16830 28254 16882
rect 28254 16830 28306 16882
rect 28306 16830 28308 16882
rect 28252 16828 28308 16830
rect 28140 15986 28196 15988
rect 28140 15934 28142 15986
rect 28142 15934 28194 15986
rect 28194 15934 28196 15986
rect 28140 15932 28196 15934
rect 26684 15372 26740 15428
rect 27132 15484 27188 15540
rect 27356 15148 27412 15204
rect 26572 13356 26628 13412
rect 26908 12796 26964 12852
rect 27244 13580 27300 13636
rect 26684 11506 26740 11508
rect 26684 11454 26686 11506
rect 26686 11454 26738 11506
rect 26738 11454 26740 11506
rect 26684 11452 26740 11454
rect 30828 19906 30884 19908
rect 30828 19854 30830 19906
rect 30830 19854 30882 19906
rect 30882 19854 30884 19906
rect 30828 19852 30884 19854
rect 30044 18956 30100 19012
rect 29036 18732 29092 18788
rect 29148 17948 29204 18004
rect 29036 16716 29092 16772
rect 29148 15596 29204 15652
rect 33516 20018 33572 20020
rect 33516 19966 33518 20018
rect 33518 19966 33570 20018
rect 33570 19966 33572 20018
rect 33516 19964 33572 19966
rect 32172 19852 32228 19908
rect 32732 19234 32788 19236
rect 32732 19182 32734 19234
rect 32734 19182 32786 19234
rect 32786 19182 32788 19234
rect 32732 19180 32788 19182
rect 33964 20690 34020 20692
rect 33964 20638 33966 20690
rect 33966 20638 34018 20690
rect 34018 20638 34020 20690
rect 33964 20636 34020 20638
rect 34300 21532 34356 21588
rect 36540 23714 36596 23716
rect 36540 23662 36542 23714
rect 36542 23662 36594 23714
rect 36594 23662 36596 23714
rect 36540 23660 36596 23662
rect 36092 22988 36148 23044
rect 38780 25564 38836 25620
rect 38444 23996 38500 24052
rect 37548 23884 37604 23940
rect 38108 23938 38164 23940
rect 38108 23886 38110 23938
rect 38110 23886 38162 23938
rect 38162 23886 38164 23938
rect 38108 23884 38164 23886
rect 35980 22092 36036 22148
rect 36988 22092 37044 22148
rect 34860 21756 34916 21812
rect 35756 21532 35812 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34748 20860 34804 20916
rect 36428 20914 36484 20916
rect 36428 20862 36430 20914
rect 36430 20862 36482 20914
rect 36482 20862 36484 20914
rect 36428 20860 36484 20862
rect 37212 21644 37268 21700
rect 37212 20860 37268 20916
rect 34188 19964 34244 20020
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34188 19180 34244 19236
rect 35980 19516 36036 19572
rect 33964 19068 34020 19124
rect 32844 19010 32900 19012
rect 32844 18958 32846 19010
rect 32846 18958 32898 19010
rect 32898 18958 32900 19010
rect 32844 18956 32900 18958
rect 35644 18956 35700 19012
rect 32060 18450 32116 18452
rect 32060 18398 32062 18450
rect 32062 18398 32114 18450
rect 32114 18398 32116 18450
rect 32060 18396 32116 18398
rect 32508 18450 32564 18452
rect 32508 18398 32510 18450
rect 32510 18398 32562 18450
rect 32562 18398 32564 18450
rect 32508 18396 32564 18398
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 31948 17836 32004 17892
rect 29596 17500 29652 17556
rect 32172 17052 32228 17108
rect 29596 16268 29652 16324
rect 30044 16828 30100 16884
rect 29708 14588 29764 14644
rect 27804 11452 27860 11508
rect 28028 12684 28084 12740
rect 30940 16268 30996 16324
rect 30268 15820 30324 15876
rect 30268 15372 30324 15428
rect 30156 15148 30212 15204
rect 29372 12684 29428 12740
rect 30828 14476 30884 14532
rect 31388 15932 31444 15988
rect 31052 15426 31108 15428
rect 31052 15374 31054 15426
rect 31054 15374 31106 15426
rect 31106 15374 31108 15426
rect 31052 15372 31108 15374
rect 32620 17500 32676 17556
rect 32844 17442 32900 17444
rect 32844 17390 32846 17442
rect 32846 17390 32898 17442
rect 32898 17390 32900 17442
rect 32844 17388 32900 17390
rect 32508 16716 32564 16772
rect 31836 15484 31892 15540
rect 31948 15596 32004 15652
rect 31724 15426 31780 15428
rect 31724 15374 31726 15426
rect 31726 15374 31778 15426
rect 31778 15374 31780 15426
rect 31724 15372 31780 15374
rect 33180 16716 33236 16772
rect 31164 12850 31220 12852
rect 31164 12798 31166 12850
rect 31166 12798 31218 12850
rect 31218 12798 31220 12850
rect 31164 12796 31220 12798
rect 29036 12066 29092 12068
rect 29036 12014 29038 12066
rect 29038 12014 29090 12066
rect 29090 12014 29092 12066
rect 29036 12012 29092 12014
rect 33068 15426 33124 15428
rect 33068 15374 33070 15426
rect 33070 15374 33122 15426
rect 33122 15374 33124 15426
rect 33068 15372 33124 15374
rect 33292 15314 33348 15316
rect 33292 15262 33294 15314
rect 33294 15262 33346 15314
rect 33346 15262 33348 15314
rect 33292 15260 33348 15262
rect 35532 17388 35588 17444
rect 34972 16716 35028 16772
rect 33740 15314 33796 15316
rect 33740 15262 33742 15314
rect 33742 15262 33794 15314
rect 33794 15262 33796 15314
rect 33740 15260 33796 15262
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 33964 15202 34020 15204
rect 33964 15150 33966 15202
rect 33966 15150 34018 15202
rect 34018 15150 34020 15202
rect 33964 15148 34020 15150
rect 34748 15202 34804 15204
rect 34748 15150 34750 15202
rect 34750 15150 34802 15202
rect 34802 15150 34804 15202
rect 34748 15148 34804 15150
rect 34300 14642 34356 14644
rect 34300 14590 34302 14642
rect 34302 14590 34354 14642
rect 34354 14590 34356 14642
rect 34300 14588 34356 14590
rect 33516 14252 33572 14308
rect 34300 14252 34356 14308
rect 32732 13468 32788 13524
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35308 14418 35364 14420
rect 35308 14366 35310 14418
rect 35310 14366 35362 14418
rect 35362 14366 35364 14418
rect 35308 14364 35364 14366
rect 35644 14140 35700 14196
rect 35420 13468 35476 13524
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34860 12684 34916 12740
rect 32508 12012 32564 12068
rect 34076 12066 34132 12068
rect 34076 12014 34078 12066
rect 34078 12014 34130 12066
rect 34130 12014 34132 12066
rect 34076 12012 34132 12014
rect 33516 11506 33572 11508
rect 33516 11454 33518 11506
rect 33518 11454 33570 11506
rect 33570 11454 33572 11506
rect 33516 11452 33572 11454
rect 36092 18956 36148 19012
rect 35980 17724 36036 17780
rect 38892 25004 38948 25060
rect 39004 24668 39060 24724
rect 39676 24722 39732 24724
rect 39676 24670 39678 24722
rect 39678 24670 39730 24722
rect 39730 24670 39732 24722
rect 39676 24668 39732 24670
rect 39004 23996 39060 24052
rect 40460 27970 40516 27972
rect 40460 27918 40462 27970
rect 40462 27918 40514 27970
rect 40514 27918 40516 27970
rect 40460 27916 40516 27918
rect 40572 27580 40628 27636
rect 42812 28530 42868 28532
rect 42812 28478 42814 28530
rect 42814 28478 42866 28530
rect 42866 28478 42868 28530
rect 42812 28476 42868 28478
rect 42924 27970 42980 27972
rect 42924 27918 42926 27970
rect 42926 27918 42978 27970
rect 42978 27918 42980 27970
rect 42924 27916 42980 27918
rect 41916 27746 41972 27748
rect 41916 27694 41918 27746
rect 41918 27694 41970 27746
rect 41970 27694 41972 27746
rect 41916 27692 41972 27694
rect 42812 27580 42868 27636
rect 41804 27186 41860 27188
rect 41804 27134 41806 27186
rect 41806 27134 41858 27186
rect 41858 27134 41860 27186
rect 41804 27132 41860 27134
rect 40124 26460 40180 26516
rect 40684 26908 40740 26964
rect 42924 26402 42980 26404
rect 42924 26350 42926 26402
rect 42926 26350 42978 26402
rect 42978 26350 42980 26402
rect 42924 26348 42980 26350
rect 41916 26178 41972 26180
rect 41916 26126 41918 26178
rect 41918 26126 41970 26178
rect 41970 26126 41972 26178
rect 41916 26124 41972 26126
rect 43932 26962 43988 26964
rect 43932 26910 43934 26962
rect 43934 26910 43986 26962
rect 43986 26910 43988 26962
rect 43932 26908 43988 26910
rect 43820 26514 43876 26516
rect 43820 26462 43822 26514
rect 43822 26462 43874 26514
rect 43874 26462 43876 26514
rect 43820 26460 43876 26462
rect 42476 25618 42532 25620
rect 42476 25566 42478 25618
rect 42478 25566 42530 25618
rect 42530 25566 42532 25618
rect 42476 25564 42532 25566
rect 41244 25394 41300 25396
rect 41244 25342 41246 25394
rect 41246 25342 41298 25394
rect 41298 25342 41300 25394
rect 41244 25340 41300 25342
rect 41916 24610 41972 24612
rect 41916 24558 41918 24610
rect 41918 24558 41970 24610
rect 41970 24558 41972 24610
rect 41916 24556 41972 24558
rect 42252 23996 42308 24052
rect 41244 23772 41300 23828
rect 42028 23826 42084 23828
rect 42028 23774 42030 23826
rect 42030 23774 42082 23826
rect 42082 23774 42084 23826
rect 42028 23772 42084 23774
rect 39788 23436 39844 23492
rect 38444 21698 38500 21700
rect 38444 21646 38446 21698
rect 38446 21646 38498 21698
rect 38498 21646 38500 21698
rect 38444 21644 38500 21646
rect 39452 21698 39508 21700
rect 39452 21646 39454 21698
rect 39454 21646 39506 21698
rect 39506 21646 39508 21698
rect 39452 21644 39508 21646
rect 37548 21420 37604 21476
rect 37884 21362 37940 21364
rect 37884 21310 37886 21362
rect 37886 21310 37938 21362
rect 37938 21310 37940 21362
rect 37884 21308 37940 21310
rect 38444 20860 38500 20916
rect 36204 18396 36260 18452
rect 36540 19234 36596 19236
rect 36540 19182 36542 19234
rect 36542 19182 36594 19234
rect 36594 19182 36596 19234
rect 36540 19180 36596 19182
rect 36652 17388 36708 17444
rect 38780 20748 38836 20804
rect 40012 22204 40068 22260
rect 40460 21644 40516 21700
rect 40572 20636 40628 20692
rect 40908 22092 40964 22148
rect 41468 21532 41524 21588
rect 38220 19906 38276 19908
rect 38220 19854 38222 19906
rect 38222 19854 38274 19906
rect 38274 19854 38276 19906
rect 38220 19852 38276 19854
rect 37884 19346 37940 19348
rect 37884 19294 37886 19346
rect 37886 19294 37938 19346
rect 37938 19294 37940 19346
rect 37884 19292 37940 19294
rect 39228 19740 39284 19796
rect 38892 19292 38948 19348
rect 37772 19180 37828 19236
rect 39116 19234 39172 19236
rect 39116 19182 39118 19234
rect 39118 19182 39170 19234
rect 39170 19182 39172 19234
rect 39116 19180 39172 19182
rect 38780 19010 38836 19012
rect 38780 18958 38782 19010
rect 38782 18958 38834 19010
rect 38834 18958 38836 19010
rect 38780 18956 38836 18958
rect 39788 18508 39844 18564
rect 39340 18450 39396 18452
rect 39340 18398 39342 18450
rect 39342 18398 39394 18450
rect 39394 18398 39396 18450
rect 39340 18396 39396 18398
rect 38780 18284 38836 18340
rect 37100 16940 37156 16996
rect 37212 17052 37268 17108
rect 36988 16882 37044 16884
rect 36988 16830 36990 16882
rect 36990 16830 37042 16882
rect 37042 16830 37044 16882
rect 36988 16828 37044 16830
rect 36316 15148 36372 15204
rect 36876 14812 36932 14868
rect 36540 14252 36596 14308
rect 37548 16716 37604 16772
rect 37436 16156 37492 16212
rect 37660 16604 37716 16660
rect 38108 15372 38164 15428
rect 39564 18284 39620 18340
rect 40236 18284 40292 18340
rect 40348 16828 40404 16884
rect 38892 15426 38948 15428
rect 38892 15374 38894 15426
rect 38894 15374 38946 15426
rect 38946 15374 38948 15426
rect 38892 15372 38948 15374
rect 38780 15148 38836 15204
rect 39116 15148 39172 15204
rect 38220 14812 38276 14868
rect 37660 14418 37716 14420
rect 37660 14366 37662 14418
rect 37662 14366 37714 14418
rect 37714 14366 37716 14418
rect 37660 14364 37716 14366
rect 37996 14140 38052 14196
rect 40012 15036 40068 15092
rect 38668 13916 38724 13972
rect 39004 14252 39060 14308
rect 40572 15932 40628 15988
rect 42812 23660 42868 23716
rect 41916 23042 41972 23044
rect 41916 22990 41918 23042
rect 41918 22990 41970 23042
rect 41970 22990 41972 23042
rect 41916 22988 41972 22990
rect 42924 22540 42980 22596
rect 41804 21756 41860 21812
rect 42476 21532 42532 21588
rect 41916 21474 41972 21476
rect 41916 21422 41918 21474
rect 41918 21422 41970 21474
rect 41970 21422 41972 21474
rect 41916 21420 41972 21422
rect 42252 21420 42308 21476
rect 41580 20076 41636 20132
rect 41916 19516 41972 19572
rect 41916 19068 41972 19124
rect 41692 18508 41748 18564
rect 42700 20914 42756 20916
rect 42700 20862 42702 20914
rect 42702 20862 42754 20914
rect 42754 20862 42756 20914
rect 42700 20860 42756 20862
rect 42924 21698 42980 21700
rect 42924 21646 42926 21698
rect 42926 21646 42978 21698
rect 42978 21646 42980 21698
rect 42924 21644 42980 21646
rect 43708 25394 43764 25396
rect 43708 25342 43710 25394
rect 43710 25342 43762 25394
rect 43762 25342 43764 25394
rect 43708 25340 43764 25342
rect 43596 23996 43652 24052
rect 43484 22316 43540 22372
rect 43932 22204 43988 22260
rect 43708 22146 43764 22148
rect 43708 22094 43710 22146
rect 43710 22094 43762 22146
rect 43762 22094 43764 22146
rect 43708 22092 43764 22094
rect 43596 21532 43652 21588
rect 43932 21474 43988 21476
rect 43932 21422 43934 21474
rect 43934 21422 43986 21474
rect 43986 21422 43988 21474
rect 43932 21420 43988 21422
rect 43148 21308 43204 21364
rect 43708 20690 43764 20692
rect 43708 20638 43710 20690
rect 43710 20638 43762 20690
rect 43762 20638 43764 20690
rect 43708 20636 43764 20638
rect 42924 20130 42980 20132
rect 42924 20078 42926 20130
rect 42926 20078 42978 20130
rect 42978 20078 42980 20130
rect 42924 20076 42980 20078
rect 41804 17778 41860 17780
rect 41804 17726 41806 17778
rect 41806 17726 41858 17778
rect 41858 17726 41860 17778
rect 41804 17724 41860 17726
rect 42812 17554 42868 17556
rect 42812 17502 42814 17554
rect 42814 17502 42866 17554
rect 42866 17502 42868 17554
rect 42812 17500 42868 17502
rect 43596 18284 43652 18340
rect 42924 17388 42980 17444
rect 42924 16994 42980 16996
rect 42924 16942 42926 16994
rect 42926 16942 42978 16994
rect 42978 16942 42980 16994
rect 42924 16940 42980 16942
rect 41916 16770 41972 16772
rect 41916 16718 41918 16770
rect 41918 16718 41970 16770
rect 41970 16718 41972 16770
rect 41916 16716 41972 16718
rect 43932 16604 43988 16660
rect 41804 16210 41860 16212
rect 41804 16158 41806 16210
rect 41806 16158 41858 16210
rect 41858 16158 41860 16210
rect 41804 16156 41860 16158
rect 41468 15372 41524 15428
rect 40460 15148 40516 15204
rect 42812 15986 42868 15988
rect 42812 15934 42814 15986
rect 42814 15934 42866 15986
rect 42866 15934 42868 15986
rect 42812 15932 42868 15934
rect 42924 15426 42980 15428
rect 42924 15374 42926 15426
rect 42926 15374 42978 15426
rect 42978 15374 42980 15426
rect 42924 15372 42980 15374
rect 42924 15148 42980 15204
rect 41804 15036 41860 15092
rect 44044 14364 44100 14420
rect 42028 13916 42084 13972
rect 40012 13020 40068 13076
rect 40796 13074 40852 13076
rect 40796 13022 40798 13074
rect 40798 13022 40850 13074
rect 40850 13022 40852 13074
rect 40796 13020 40852 13022
rect 36876 12684 36932 12740
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 43596 8930 43652 8932
rect 43596 8878 43598 8930
rect 43598 8878 43650 8930
rect 43650 8878 43652 8930
rect 43596 8876 43652 8878
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19516 4226 19572 4228
rect 19516 4174 19518 4226
rect 19518 4174 19570 4226
rect 19570 4174 19572 4226
rect 19516 4172 19572 4174
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 20188 4060 20244 4116
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21532 3276 21588 3332
rect 22652 3330 22708 3332
rect 22652 3278 22654 3330
rect 22654 3278 22706 3330
rect 22706 3278 22708 3330
rect 22652 3276 22708 3278
rect 23660 3276 23716 3332
rect 24892 4284 24948 4340
rect 24556 3330 24612 3332
rect 24556 3278 24558 3330
rect 24558 3278 24610 3330
rect 24610 3278 24612 3330
rect 24556 3276 24612 3278
rect 25564 4338 25620 4340
rect 25564 4286 25566 4338
rect 25566 4286 25618 4338
rect 25618 4286 25620 4338
rect 25564 4284 25620 4286
rect 25564 3612 25620 3668
rect 26236 4226 26292 4228
rect 26236 4174 26238 4226
rect 26238 4174 26290 4226
rect 26290 4174 26292 4226
rect 26236 4172 26292 4174
rect 27356 4172 27412 4228
rect 26572 3666 26628 3668
rect 26572 3614 26574 3666
rect 26574 3614 26626 3666
rect 26626 3614 26628 3666
rect 26572 3612 26628 3614
rect 27580 3612 27636 3668
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 41804 5852 41860 5908
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35756 5180 35812 5236
rect 28812 3666 28868 3668
rect 28812 3614 28814 3666
rect 28814 3614 28866 3666
rect 28866 3614 28868 3666
rect 28812 3612 28868 3614
rect 31612 3612 31668 3668
rect 32172 4226 32228 4228
rect 32172 4174 32174 4226
rect 32174 4174 32226 4226
rect 32226 4174 32228 4226
rect 32172 4172 32228 4174
rect 32956 4172 33012 4228
rect 32620 3666 32676 3668
rect 32620 3614 32622 3666
rect 32622 3614 32674 3666
rect 32674 3614 32676 3666
rect 32620 3612 32676 3614
rect 37884 5180 37940 5236
rect 36428 5068 36484 5124
rect 38108 5122 38164 5124
rect 38108 5070 38110 5122
rect 38110 5070 38162 5122
rect 38162 5070 38164 5122
rect 38108 5068 38164 5070
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34972 3500 35028 3556
rect 36092 3500 36148 3556
rect 39228 5010 39284 5012
rect 39228 4958 39230 5010
rect 39230 4958 39282 5010
rect 39282 4958 39284 5010
rect 39228 4956 39284 4958
rect 40908 4956 40964 5012
rect 37996 4396 38052 4452
rect 37660 4226 37716 4228
rect 37660 4174 37662 4226
rect 37662 4174 37714 4226
rect 37714 4174 37716 4226
rect 37660 4172 37716 4174
rect 38556 4172 38612 4228
rect 38220 3500 38276 3556
rect 39004 3612 39060 3668
rect 39564 3388 39620 3444
rect 40236 3666 40292 3668
rect 40236 3614 40238 3666
rect 40238 3614 40290 3666
rect 40290 3614 40292 3666
rect 40236 3612 40292 3614
rect 39788 3554 39844 3556
rect 39788 3502 39790 3554
rect 39790 3502 39842 3554
rect 39842 3502 39844 3554
rect 39788 3500 39844 3502
rect 41468 4508 41524 4564
rect 41580 4450 41636 4452
rect 41580 4398 41582 4450
rect 41582 4398 41634 4450
rect 41634 4398 41636 4450
rect 41580 4396 41636 4398
rect 42588 6748 42644 6804
rect 42252 4844 42308 4900
rect 42140 4172 42196 4228
rect 42924 5906 42980 5908
rect 42924 5854 42926 5906
rect 42926 5854 42978 5906
rect 42978 5854 42980 5906
rect 42924 5852 42980 5854
rect 43036 4732 43092 4788
rect 44156 8764 44212 8820
rect 44044 8146 44100 8148
rect 44044 8094 44046 8146
rect 44046 8094 44098 8146
rect 44098 8094 44100 8146
rect 44044 8092 44100 8094
rect 44044 7474 44100 7476
rect 44044 7422 44046 7474
rect 44046 7422 44098 7474
rect 44098 7422 44100 7474
rect 44044 7420 44100 7422
rect 44044 6076 44100 6132
rect 44044 5404 44100 5460
rect 44156 4844 44212 4900
rect 43148 4620 43204 4676
rect 43820 4620 43876 4676
rect 43036 4508 43092 4564
rect 42700 4284 42756 4340
rect 42364 4060 42420 4116
rect 41804 3442 41860 3444
rect 41804 3390 41806 3442
rect 41806 3390 41858 3442
rect 41858 3390 41860 3442
rect 41804 3388 41860 3390
rect 44044 4338 44100 4340
rect 44044 4286 44046 4338
rect 44046 4286 44098 4338
rect 44098 4286 44100 4338
rect 44044 4284 44100 4286
rect 43820 4172 43876 4228
rect 44156 3442 44212 3444
rect 44156 3390 44158 3442
rect 44158 3390 44210 3442
rect 44210 3390 44212 3442
rect 44156 3388 44212 3390
rect 44380 4284 44436 4340
rect 43148 2716 43204 2772
rect 44380 2044 44436 2100
<< metal3 >>
rect 45200 45780 46000 45808
rect 41906 45724 41916 45780
rect 41972 45724 46000 45780
rect 45200 45696 46000 45724
rect 45200 45108 46000 45136
rect 44258 45052 44268 45108
rect 44324 45052 46000 45108
rect 45200 45024 46000 45052
rect 45200 44436 46000 44464
rect 43922 44380 43932 44436
rect 43988 44380 46000 44436
rect 45200 44352 46000 44380
rect 45200 43764 46000 43792
rect 43698 43708 43708 43764
rect 43764 43708 46000 43764
rect 45200 43680 46000 43708
rect 45200 43092 46000 43120
rect 44370 43036 44380 43092
rect 44436 43036 46000 43092
rect 45200 43008 46000 43036
rect 45200 42420 46000 42448
rect 43474 42364 43484 42420
rect 43540 42364 46000 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 45200 42336 46000 42364
rect 14578 41916 14588 41972
rect 14644 41916 15260 41972
rect 15316 41916 15326 41972
rect 16370 41916 16380 41972
rect 16436 41916 17388 41972
rect 17444 41916 17454 41972
rect 26226 41916 26236 41972
rect 26292 41916 26908 41972
rect 26964 41916 26974 41972
rect 27906 41916 27916 41972
rect 27972 41916 28588 41972
rect 28644 41916 28654 41972
rect 38994 41916 39004 41972
rect 39060 41916 40348 41972
rect 40404 41916 40414 41972
rect 43138 41804 43148 41860
rect 43204 41804 44156 41860
rect 44212 41804 44492 41860
rect 44548 41804 44558 41860
rect 45200 41748 46000 41776
rect 44034 41692 44044 41748
rect 44100 41692 46000 41748
rect 45200 41664 46000 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 18162 41356 18172 41412
rect 18228 41356 19292 41412
rect 19348 41356 19358 41412
rect 24882 41244 24892 41300
rect 24948 41244 26012 41300
rect 26068 41244 26078 41300
rect 15138 41132 15148 41188
rect 15204 41132 16940 41188
rect 16996 41132 17006 41188
rect 18834 41132 18844 41188
rect 18900 41132 20244 41188
rect 20188 41076 20244 41132
rect 45200 41076 46000 41104
rect 20178 41020 20188 41076
rect 20244 41020 20254 41076
rect 44482 41020 44492 41076
rect 44548 41020 46000 41076
rect 45200 40992 46000 41020
rect 38210 40908 38220 40964
rect 38276 40908 39788 40964
rect 39844 40908 39854 40964
rect 41682 40908 41692 40964
rect 41748 40908 43708 40964
rect 40114 40796 40124 40852
rect 40180 40796 41804 40852
rect 41860 40796 41870 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 43652 40628 43708 40908
rect 39554 40572 39564 40628
rect 39620 40572 43316 40628
rect 43652 40572 43820 40628
rect 43876 40572 43886 40628
rect 43260 40516 43316 40572
rect 14466 40460 14476 40516
rect 14532 40460 15484 40516
rect 15540 40460 15550 40516
rect 36306 40460 36316 40516
rect 36372 40460 38780 40516
rect 38836 40460 38846 40516
rect 41906 40460 41916 40516
rect 41972 40460 42924 40516
rect 42980 40460 42990 40516
rect 43260 40460 43708 40516
rect 43652 40404 43708 40460
rect 45200 40404 46000 40432
rect 41682 40348 41692 40404
rect 41748 40348 43484 40404
rect 43540 40348 43550 40404
rect 43652 40348 46000 40404
rect 45200 40320 46000 40348
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 45200 39732 46000 39760
rect 40338 39676 40348 39732
rect 40404 39676 46000 39732
rect 45200 39648 46000 39676
rect 37538 39564 37548 39620
rect 37604 39564 39116 39620
rect 39172 39564 39182 39620
rect 39890 39564 39900 39620
rect 39956 39564 40908 39620
rect 40964 39564 40974 39620
rect 42802 39452 42812 39508
rect 42868 39452 43820 39508
rect 43876 39452 43886 39508
rect 42242 39340 42252 39396
rect 42308 39340 43372 39396
rect 43428 39340 43438 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 45200 39060 46000 39088
rect 42354 39004 42364 39060
rect 42420 39004 46000 39060
rect 45200 38976 46000 39004
rect 26226 38556 26236 38612
rect 26292 38556 28364 38612
rect 28420 38556 28430 38612
rect 42802 38556 42812 38612
rect 42868 38556 43708 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 43652 38388 43708 38556
rect 45200 38388 46000 38416
rect 43652 38332 46000 38388
rect 45200 38304 46000 38332
rect 43138 38108 43148 38164
rect 43204 38108 44044 38164
rect 44100 38108 44380 38164
rect 44436 38108 44446 38164
rect 43474 37772 43484 37828
rect 43540 37772 43708 37828
rect 43652 37716 43708 37772
rect 45200 37716 46000 37744
rect 43652 37660 46000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 45200 37632 46000 37660
rect 45200 37044 46000 37072
rect 44146 36988 44156 37044
rect 44212 36988 46000 37044
rect 45200 36960 46000 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 45200 36372 46000 36400
rect 43698 36316 43708 36372
rect 43764 36316 46000 36372
rect 45200 36288 46000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 21634 35868 21644 35924
rect 21700 35868 22428 35924
rect 22484 35868 22494 35924
rect 26450 35868 26460 35924
rect 26516 35868 27132 35924
rect 27188 35868 27198 35924
rect 43652 35756 44156 35812
rect 44212 35756 44222 35812
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 43652 35028 43708 35756
rect 45200 35700 46000 35728
rect 44258 35644 44268 35700
rect 44324 35644 46000 35700
rect 45200 35616 46000 35644
rect 45200 35028 46000 35056
rect 43652 34972 46000 35028
rect 45200 34944 46000 34972
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 20290 31836 20300 31892
rect 20356 31836 22316 31892
rect 22372 31836 22382 31892
rect 45200 31668 46000 31696
rect 11554 31612 11564 31668
rect 11620 31612 12460 31668
rect 12516 31612 12526 31668
rect 16594 31612 16604 31668
rect 16660 31612 17388 31668
rect 17444 31612 17454 31668
rect 21522 31612 21532 31668
rect 21588 31612 23548 31668
rect 23604 31612 23614 31668
rect 44034 31612 44044 31668
rect 44100 31612 46000 31668
rect 45200 31584 46000 31612
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 14130 31052 14140 31108
rect 14196 31052 17164 31108
rect 17220 31052 17230 31108
rect 28018 31052 28028 31108
rect 28084 31052 31500 31108
rect 31556 31052 31566 31108
rect 32722 31052 32732 31108
rect 32788 31052 34636 31108
rect 34692 31052 34702 31108
rect 42466 31052 42476 31108
rect 42532 31052 43820 31108
rect 43876 31052 43886 31108
rect 45200 30996 46000 31024
rect 43586 30940 43596 30996
rect 43652 30940 44156 30996
rect 44212 30940 46000 30996
rect 45200 30912 46000 30940
rect 27010 30828 27020 30884
rect 27076 30828 30492 30884
rect 30548 30828 30558 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 20290 30380 20300 30436
rect 20356 30380 22540 30436
rect 22596 30380 22606 30436
rect 11218 30268 11228 30324
rect 11284 30268 12124 30324
rect 12180 30268 12190 30324
rect 21746 30268 21756 30324
rect 21812 30268 23100 30324
rect 23156 30268 23166 30324
rect 24658 30268 24668 30324
rect 24724 30268 25900 30324
rect 25956 30268 25966 30324
rect 5282 30044 5292 30100
rect 5348 30044 7644 30100
rect 7700 30044 7710 30100
rect 17938 30044 17948 30100
rect 18004 30044 20188 30100
rect 20244 30044 20254 30100
rect 23314 30044 23324 30100
rect 23380 30044 24108 30100
rect 24164 30044 24174 30100
rect 24770 30044 24780 30100
rect 24836 30044 26908 30100
rect 26964 30044 26974 30100
rect 28018 30044 28028 30100
rect 28084 30044 29484 30100
rect 29540 30044 29550 30100
rect 32610 30044 32620 30100
rect 32676 30044 34860 30100
rect 34916 30044 34926 30100
rect 36530 30044 36540 30100
rect 36596 30044 39004 30100
rect 39060 30044 39070 30100
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 24210 29596 24220 29652
rect 24276 29596 25340 29652
rect 25396 29596 25406 29652
rect 21634 29484 21644 29540
rect 21700 29484 25228 29540
rect 25284 29484 25294 29540
rect 34178 29484 34188 29540
rect 34244 29484 37884 29540
rect 37940 29484 37950 29540
rect 9986 29372 9996 29428
rect 10052 29372 11452 29428
rect 11508 29372 11518 29428
rect 14466 29372 14476 29428
rect 14532 29372 17500 29428
rect 17556 29372 19628 29428
rect 19684 29372 19694 29428
rect 6178 29260 6188 29316
rect 6244 29260 7532 29316
rect 7588 29260 7598 29316
rect 25778 29260 25788 29316
rect 25844 29260 27804 29316
rect 27860 29260 27870 29316
rect 29698 29260 29708 29316
rect 29764 29260 34076 29316
rect 34132 29260 34142 29316
rect 29922 29148 29932 29204
rect 29988 29148 35308 29204
rect 35364 29148 35374 29204
rect 29586 29036 29596 29092
rect 29652 29036 31052 29092
rect 31108 29036 31118 29092
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 3612 28980
rect 3668 28924 3678 28980
rect 27346 28924 27356 28980
rect 27412 28924 28700 28980
rect 28756 28924 28766 28980
rect 0 28896 800 28924
rect 33506 28812 33516 28868
rect 33572 28812 36876 28868
rect 36932 28812 36942 28868
rect 3042 28700 3052 28756
rect 3108 28700 4956 28756
rect 5012 28700 5022 28756
rect 20132 28700 22316 28756
rect 22372 28700 22382 28756
rect 31154 28700 31164 28756
rect 31220 28700 33852 28756
rect 33908 28700 33918 28756
rect 37538 28700 37548 28756
rect 37604 28700 41804 28756
rect 41860 28700 41870 28756
rect 20132 28644 20188 28700
rect 1810 28588 1820 28644
rect 1876 28588 4004 28644
rect 4834 28588 4844 28644
rect 4900 28588 5740 28644
rect 5796 28588 6748 28644
rect 6804 28588 7420 28644
rect 7476 28588 7486 28644
rect 19394 28588 19404 28644
rect 19460 28588 20188 28644
rect 3948 28532 4004 28588
rect 3938 28476 3948 28532
rect 4004 28476 4014 28532
rect 16370 28476 16380 28532
rect 16436 28476 19180 28532
rect 19236 28476 19246 28532
rect 21298 28476 21308 28532
rect 21364 28476 23996 28532
rect 24052 28476 24062 28532
rect 40786 28476 40796 28532
rect 40852 28476 42812 28532
rect 42868 28476 42878 28532
rect 20514 28364 20524 28420
rect 20580 28364 21644 28420
rect 21700 28364 21710 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 5506 27916 5516 27972
rect 5572 27916 6636 27972
rect 6692 27916 6702 27972
rect 23426 27916 23436 27972
rect 23492 27916 23996 27972
rect 24052 27916 24062 27972
rect 40450 27916 40460 27972
rect 40516 27916 42924 27972
rect 42980 27916 42990 27972
rect 3826 27804 3836 27860
rect 3892 27804 5292 27860
rect 5348 27804 5358 27860
rect 5730 27804 5740 27860
rect 5796 27804 7868 27860
rect 7924 27804 9324 27860
rect 9380 27804 9390 27860
rect 23874 27804 23884 27860
rect 23940 27804 25116 27860
rect 25172 27804 26236 27860
rect 26292 27804 28588 27860
rect 28644 27804 29036 27860
rect 29092 27804 29102 27860
rect 3042 27692 3052 27748
rect 3108 27692 4284 27748
rect 4340 27692 4350 27748
rect 7634 27692 7644 27748
rect 7700 27692 8540 27748
rect 8596 27692 8606 27748
rect 9874 27692 9884 27748
rect 9940 27692 10780 27748
rect 10836 27692 10846 27748
rect 16818 27692 16828 27748
rect 16884 27692 17724 27748
rect 17780 27692 17790 27748
rect 37538 27692 37548 27748
rect 37604 27692 41916 27748
rect 41972 27692 41982 27748
rect 0 27636 800 27664
rect 0 27580 1708 27636
rect 1764 27580 1774 27636
rect 31490 27580 31500 27636
rect 31556 27580 32956 27636
rect 33012 27580 33022 27636
rect 40562 27580 40572 27636
rect 40628 27580 42812 27636
rect 42868 27580 42878 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 8372 27356 9548 27412
rect 9604 27356 9614 27412
rect 8372 27076 8428 27356
rect 19394 27132 19404 27188
rect 19460 27132 23548 27188
rect 23604 27132 23614 27188
rect 38210 27132 38220 27188
rect 38276 27132 41804 27188
rect 41860 27132 41870 27188
rect 3938 27020 3948 27076
rect 4004 27020 5516 27076
rect 5572 27020 5582 27076
rect 6290 27020 6300 27076
rect 6356 27020 8428 27076
rect 10770 27020 10780 27076
rect 10836 27020 11900 27076
rect 11956 27020 13916 27076
rect 13972 27020 13982 27076
rect 17714 27020 17724 27076
rect 17780 27020 19852 27076
rect 19908 27020 20636 27076
rect 20692 27020 20702 27076
rect 12226 26908 12236 26964
rect 12292 26908 14812 26964
rect 14868 26908 14878 26964
rect 19058 26908 19068 26964
rect 19124 26908 19628 26964
rect 19684 26908 19694 26964
rect 26562 26908 26572 26964
rect 26628 26908 27580 26964
rect 27636 26908 27646 26964
rect 27906 26908 27916 26964
rect 27972 26908 29260 26964
rect 29316 26908 31388 26964
rect 31444 26908 31454 26964
rect 33058 26908 33068 26964
rect 33124 26908 34076 26964
rect 34132 26908 34142 26964
rect 34850 26908 34860 26964
rect 34916 26908 36316 26964
rect 36372 26908 36382 26964
rect 40674 26908 40684 26964
rect 40740 26908 43932 26964
rect 43988 26908 43998 26964
rect 9762 26796 9772 26852
rect 9828 26796 11564 26852
rect 11620 26796 12796 26852
rect 12852 26796 12862 26852
rect 19170 26796 19180 26852
rect 19236 26796 19516 26852
rect 19572 26796 19582 26852
rect 22082 26796 22092 26852
rect 22148 26796 23212 26852
rect 23268 26796 23278 26852
rect 34514 26796 34524 26852
rect 34580 26796 37996 26852
rect 38052 26796 38062 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 40114 26460 40124 26516
rect 40180 26460 43820 26516
rect 43876 26460 43886 26516
rect 18834 26348 18844 26404
rect 18900 26348 19628 26404
rect 19684 26348 19694 26404
rect 37538 26348 37548 26404
rect 37604 26348 42924 26404
rect 42980 26348 42990 26404
rect 14802 26236 14812 26292
rect 14868 26236 15596 26292
rect 15652 26236 21868 26292
rect 21924 26236 23828 26292
rect 33394 26236 33404 26292
rect 33460 26236 35644 26292
rect 35700 26236 35710 26292
rect 23772 26180 23828 26236
rect 2818 26124 2828 26180
rect 2884 26124 3724 26180
rect 3780 26124 3790 26180
rect 8372 26124 8876 26180
rect 8932 26124 11004 26180
rect 11060 26124 11070 26180
rect 12562 26124 12572 26180
rect 12628 26124 15148 26180
rect 15204 26124 15214 26180
rect 15810 26124 15820 26180
rect 15876 26124 16716 26180
rect 16772 26124 16782 26180
rect 19170 26124 19180 26180
rect 19236 26124 19628 26180
rect 19684 26124 19694 26180
rect 23762 26124 23772 26180
rect 23828 26124 26796 26180
rect 26852 26124 32172 26180
rect 32228 26124 32238 26180
rect 7410 26012 7420 26068
rect 7476 26012 8316 26068
rect 8372 26012 8428 26124
rect 33404 26068 33460 26236
rect 37426 26124 37436 26180
rect 37492 26124 41916 26180
rect 41972 26124 41982 26180
rect 8642 26012 8652 26068
rect 8708 26012 12908 26068
rect 12964 26012 12974 26068
rect 31378 26012 31388 26068
rect 31444 26012 33460 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14018 25676 14028 25732
rect 14084 25676 16492 25732
rect 16548 25676 16558 25732
rect 3714 25564 3724 25620
rect 3780 25564 4508 25620
rect 4564 25564 7420 25620
rect 7476 25564 7486 25620
rect 14914 25564 14924 25620
rect 14980 25564 16884 25620
rect 17042 25564 17052 25620
rect 17108 25564 20300 25620
rect 20356 25564 20366 25620
rect 21746 25564 21756 25620
rect 21812 25564 22876 25620
rect 22932 25564 22942 25620
rect 24322 25564 24332 25620
rect 24388 25564 25676 25620
rect 25732 25564 25742 25620
rect 35634 25564 35644 25620
rect 35700 25564 36988 25620
rect 37044 25564 37054 25620
rect 38770 25564 38780 25620
rect 38836 25564 42476 25620
rect 42532 25564 42542 25620
rect 16828 25508 16884 25564
rect 13346 25452 13356 25508
rect 13412 25452 15148 25508
rect 16818 25452 16828 25508
rect 16884 25452 16894 25508
rect 13234 25340 13244 25396
rect 13300 25340 13580 25396
rect 13636 25340 13646 25396
rect 15092 25284 15148 25452
rect 23314 25340 23324 25396
rect 23380 25340 23884 25396
rect 23940 25340 23950 25396
rect 24770 25340 24780 25396
rect 24836 25340 26908 25396
rect 26964 25340 26974 25396
rect 28802 25340 28812 25396
rect 28868 25340 33964 25396
rect 34020 25340 34030 25396
rect 41234 25340 41244 25396
rect 41300 25340 43708 25396
rect 43764 25340 43774 25396
rect 6962 25228 6972 25284
rect 7028 25228 9324 25284
rect 9380 25228 9390 25284
rect 15092 25228 16268 25284
rect 16324 25228 16940 25284
rect 16996 25228 17006 25284
rect 17938 25228 17948 25284
rect 18004 25228 20412 25284
rect 20468 25228 20478 25284
rect 32162 25228 32172 25284
rect 32228 25228 33628 25284
rect 33684 25228 33694 25284
rect 33842 25228 33852 25284
rect 33908 25228 37100 25284
rect 37156 25228 37166 25284
rect 27010 25116 27020 25172
rect 27076 25116 32956 25172
rect 33012 25116 33022 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 20300 25004 29932 25060
rect 29988 25004 29998 25060
rect 33506 25004 33516 25060
rect 33572 25004 38892 25060
rect 38948 25004 38958 25060
rect 10098 24892 10108 24948
rect 10164 24892 13468 24948
rect 13524 24892 13534 24948
rect 9426 24780 9436 24836
rect 9492 24780 10220 24836
rect 10276 24780 10286 24836
rect 20300 24724 20356 25004
rect 7970 24668 7980 24724
rect 8036 24668 10108 24724
rect 10164 24668 10174 24724
rect 16930 24668 16940 24724
rect 16996 24668 19628 24724
rect 19684 24668 19694 24724
rect 20290 24668 20300 24724
rect 20356 24668 20366 24724
rect 26450 24668 26460 24724
rect 26516 24668 27132 24724
rect 27188 24668 28588 24724
rect 28644 24668 29036 24724
rect 29092 24668 29102 24724
rect 31042 24668 31052 24724
rect 31108 24668 31612 24724
rect 31668 24668 32284 24724
rect 32340 24668 32350 24724
rect 38994 24668 39004 24724
rect 39060 24668 39676 24724
rect 39732 24668 39742 24724
rect 19394 24556 19404 24612
rect 19460 24556 23884 24612
rect 23940 24556 24444 24612
rect 24500 24556 24510 24612
rect 30146 24556 30156 24612
rect 30212 24556 32060 24612
rect 32116 24556 32126 24612
rect 37426 24556 37436 24612
rect 37492 24556 41916 24612
rect 41972 24556 41982 24612
rect 18386 24444 18396 24500
rect 18452 24444 21532 24500
rect 21588 24444 24332 24500
rect 24388 24444 26236 24500
rect 26292 24444 26302 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 6738 24108 6748 24164
rect 6804 24108 11900 24164
rect 11956 24108 11966 24164
rect 4050 23996 4060 24052
rect 4116 23996 8428 24052
rect 10994 23996 11004 24052
rect 11060 23996 12572 24052
rect 12628 23996 13692 24052
rect 13748 23996 15484 24052
rect 15540 23996 16380 24052
rect 16436 23996 17612 24052
rect 17668 23996 17678 24052
rect 23314 23996 23324 24052
rect 23380 23996 25228 24052
rect 25284 23996 25294 24052
rect 35522 23996 35532 24052
rect 35588 23996 37212 24052
rect 37268 23996 38444 24052
rect 38500 23996 39004 24052
rect 39060 23996 42252 24052
rect 42308 23996 43596 24052
rect 43652 23996 43662 24052
rect 8372 23940 8428 23996
rect 8372 23884 9996 23940
rect 10052 23884 10062 23940
rect 20850 23884 20860 23940
rect 20916 23884 24556 23940
rect 24612 23884 25788 23940
rect 25844 23884 26460 23940
rect 26516 23884 26526 23940
rect 30034 23884 30044 23940
rect 30100 23884 32844 23940
rect 32900 23884 34076 23940
rect 34132 23884 35644 23940
rect 35700 23884 36428 23940
rect 36484 23884 37548 23940
rect 37604 23884 38108 23940
rect 38164 23884 38174 23940
rect 3042 23772 3052 23828
rect 3108 23772 9212 23828
rect 9268 23772 9278 23828
rect 26226 23772 26236 23828
rect 26292 23772 31948 23828
rect 32004 23772 32014 23828
rect 41234 23772 41244 23828
rect 41300 23772 42028 23828
rect 42084 23772 42094 23828
rect 16930 23660 16940 23716
rect 16996 23660 18396 23716
rect 18452 23660 18462 23716
rect 28242 23660 28252 23716
rect 28308 23660 31948 23716
rect 32004 23660 32014 23716
rect 36530 23660 36540 23716
rect 36596 23660 42812 23716
rect 42868 23660 42878 23716
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 16370 23436 16380 23492
rect 16436 23436 19068 23492
rect 19124 23436 19134 23492
rect 32946 23436 32956 23492
rect 33012 23436 39788 23492
rect 39844 23436 39854 23492
rect 6962 23324 6972 23380
rect 7028 23324 16940 23380
rect 16996 23324 17006 23380
rect 32498 23324 32508 23380
rect 32564 23324 33516 23380
rect 33572 23324 33582 23380
rect 4050 23212 4060 23268
rect 4116 23212 9436 23268
rect 9492 23212 9502 23268
rect 29922 23212 29932 23268
rect 29988 23212 31500 23268
rect 31556 23212 31566 23268
rect 12002 23100 12012 23156
rect 12068 23100 13804 23156
rect 13860 23100 13870 23156
rect 19058 23100 19068 23156
rect 19124 23100 20860 23156
rect 20916 23100 20926 23156
rect 24546 23100 24556 23156
rect 24612 23100 25452 23156
rect 25508 23100 25518 23156
rect 5170 22988 5180 23044
rect 5236 22988 9884 23044
rect 9940 22988 9950 23044
rect 13010 22988 13020 23044
rect 13076 22988 13580 23044
rect 13636 22988 15820 23044
rect 15876 22988 16828 23044
rect 16884 22988 16894 23044
rect 23090 22988 23100 23044
rect 23156 22988 24332 23044
rect 24388 22988 24398 23044
rect 28914 22988 28924 23044
rect 28980 22988 30828 23044
rect 30884 22988 30894 23044
rect 31154 22988 31164 23044
rect 31220 22988 31612 23044
rect 31668 22988 32508 23044
rect 32564 22988 32574 23044
rect 36082 22988 36092 23044
rect 36148 22988 41916 23044
rect 41972 22988 41982 23044
rect 31164 22932 31220 22988
rect 7970 22876 7980 22932
rect 8036 22876 13804 22932
rect 13860 22876 13870 22932
rect 22642 22876 22652 22932
rect 22708 22876 23996 22932
rect 24052 22876 24062 22932
rect 29362 22876 29372 22932
rect 29428 22876 29820 22932
rect 29876 22876 31220 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14914 22540 14924 22596
rect 14980 22540 16940 22596
rect 16996 22540 17006 22596
rect 29698 22540 29708 22596
rect 29764 22540 33180 22596
rect 33236 22540 33246 22596
rect 33506 22540 33516 22596
rect 33572 22540 42924 22596
rect 42980 22540 42990 22596
rect 4050 22428 4060 22484
rect 4116 22428 8540 22484
rect 8596 22428 8606 22484
rect 15922 22428 15932 22484
rect 15988 22428 17724 22484
rect 17780 22428 17790 22484
rect 27906 22428 27916 22484
rect 27972 22428 28476 22484
rect 28532 22428 29372 22484
rect 29428 22428 29438 22484
rect 31892 22428 34748 22484
rect 34804 22428 34814 22484
rect 31892 22372 31948 22428
rect 30482 22316 30492 22372
rect 30548 22316 31948 22372
rect 43474 22316 43484 22372
rect 43540 22316 44548 22372
rect 44492 22260 44548 22316
rect 45200 22260 46000 22288
rect 3042 22204 3052 22260
rect 3108 22204 6860 22260
rect 6916 22204 6926 22260
rect 14354 22204 14364 22260
rect 14420 22204 16604 22260
rect 16660 22204 16670 22260
rect 19730 22204 19740 22260
rect 19796 22204 23212 22260
rect 23268 22204 23278 22260
rect 32722 22204 32732 22260
rect 32788 22204 35756 22260
rect 35812 22204 35822 22260
rect 40002 22204 40012 22260
rect 40068 22204 43932 22260
rect 43988 22204 43998 22260
rect 44492 22204 46000 22260
rect 45200 22176 46000 22204
rect 3602 22092 3612 22148
rect 3668 22092 20860 22148
rect 20916 22092 21420 22148
rect 21476 22092 21486 22148
rect 35970 22092 35980 22148
rect 36036 22092 36988 22148
rect 37044 22092 37054 22148
rect 40898 22092 40908 22148
rect 40964 22092 43708 22148
rect 43764 22092 43774 22148
rect 11330 21980 11340 22036
rect 11396 21980 13916 22036
rect 13972 21980 13982 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 4050 21868 4060 21924
rect 4116 21868 6076 21924
rect 6132 21868 6142 21924
rect 13010 21868 13020 21924
rect 13076 21868 14364 21924
rect 14420 21868 14430 21924
rect 10210 21756 10220 21812
rect 10276 21756 11900 21812
rect 11956 21756 11966 21812
rect 18050 21756 18060 21812
rect 18116 21756 21980 21812
rect 22036 21756 22046 21812
rect 34850 21756 34860 21812
rect 34916 21756 41804 21812
rect 41860 21756 41870 21812
rect 9986 21644 9996 21700
rect 10052 21644 11788 21700
rect 11844 21644 12124 21700
rect 12180 21644 12190 21700
rect 37202 21644 37212 21700
rect 37268 21644 38444 21700
rect 38500 21644 39452 21700
rect 39508 21644 39518 21700
rect 40450 21644 40460 21700
rect 40516 21644 42924 21700
rect 42980 21644 42990 21700
rect 4722 21532 4732 21588
rect 4788 21532 6860 21588
rect 6916 21532 6926 21588
rect 15362 21532 15372 21588
rect 15428 21532 18844 21588
rect 18900 21532 18910 21588
rect 22082 21532 22092 21588
rect 22148 21532 25340 21588
rect 25396 21532 25406 21588
rect 26450 21532 26460 21588
rect 26516 21532 26908 21588
rect 32498 21532 32508 21588
rect 32564 21532 33404 21588
rect 33460 21532 33852 21588
rect 33908 21532 34300 21588
rect 34356 21532 35756 21588
rect 35812 21532 41468 21588
rect 41524 21532 42476 21588
rect 42532 21532 43596 21588
rect 43652 21532 43662 21588
rect 26852 21476 26908 21532
rect 26852 21420 30716 21476
rect 30772 21420 30782 21476
rect 37538 21420 37548 21476
rect 37604 21420 41916 21476
rect 41972 21420 41982 21476
rect 42242 21420 42252 21476
rect 42308 21420 43932 21476
rect 43988 21420 43998 21476
rect 3042 21308 3052 21364
rect 3108 21308 5404 21364
rect 5460 21308 5470 21364
rect 29474 21308 29484 21364
rect 29540 21308 31164 21364
rect 31220 21308 31230 21364
rect 37874 21308 37884 21364
rect 37940 21308 43148 21364
rect 43204 21308 43214 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 10994 20972 11004 21028
rect 11060 20972 13356 21028
rect 13412 20972 13422 21028
rect 12114 20860 12124 20916
rect 12180 20860 12796 20916
rect 12852 20860 12862 20916
rect 27570 20860 27580 20916
rect 27636 20860 30156 20916
rect 30212 20860 30222 20916
rect 31948 20860 34748 20916
rect 34804 20860 36428 20916
rect 36484 20860 37212 20916
rect 37268 20860 37278 20916
rect 38434 20860 38444 20916
rect 38500 20860 42700 20916
rect 42756 20860 42766 20916
rect 31948 20804 32004 20860
rect 7970 20748 7980 20804
rect 8036 20748 9100 20804
rect 9156 20748 9166 20804
rect 9986 20748 9996 20804
rect 10052 20748 10062 20804
rect 23650 20748 23660 20804
rect 23716 20748 25340 20804
rect 25396 20748 25406 20804
rect 27010 20748 27020 20804
rect 27076 20748 31948 20804
rect 32004 20748 32014 20804
rect 33618 20748 33628 20804
rect 33684 20748 38780 20804
rect 38836 20748 38846 20804
rect 9996 20692 10052 20748
rect 7410 20636 7420 20692
rect 7476 20636 8988 20692
rect 9044 20636 10052 20692
rect 30594 20636 30604 20692
rect 30660 20636 33964 20692
rect 34020 20636 34030 20692
rect 40562 20636 40572 20692
rect 40628 20636 43708 20692
rect 43764 20636 43774 20692
rect 9986 20524 9996 20580
rect 10052 20524 11676 20580
rect 11732 20524 11742 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 5058 20188 5068 20244
rect 5124 20188 7196 20244
rect 7252 20188 7980 20244
rect 8036 20188 8046 20244
rect 17490 20188 17500 20244
rect 17556 20188 19964 20244
rect 20020 20188 20030 20244
rect 3266 20076 3276 20132
rect 3332 20076 5964 20132
rect 6020 20076 6030 20132
rect 20178 20076 20188 20132
rect 20244 20076 22092 20132
rect 22148 20076 22158 20132
rect 41570 20076 41580 20132
rect 41636 20076 42924 20132
rect 42980 20076 42990 20132
rect 12450 19964 12460 20020
rect 12516 19964 13244 20020
rect 13300 19964 16156 20020
rect 16212 19964 16222 20020
rect 33506 19964 33516 20020
rect 33572 19964 34188 20020
rect 34244 19964 34254 20020
rect 8306 19852 8316 19908
rect 8372 19852 10108 19908
rect 10164 19852 10174 19908
rect 24322 19852 24332 19908
rect 24388 19852 30828 19908
rect 30884 19852 30894 19908
rect 32162 19852 32172 19908
rect 32228 19852 38220 19908
rect 38276 19852 38286 19908
rect 29586 19740 29596 19796
rect 29652 19740 39228 19796
rect 39284 19740 39294 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 35970 19516 35980 19572
rect 36036 19516 41916 19572
rect 41972 19516 41982 19572
rect 20290 19404 20300 19460
rect 20356 19404 21420 19460
rect 21476 19404 21486 19460
rect 6066 19292 6076 19348
rect 6132 19292 6972 19348
rect 7028 19292 7980 19348
rect 8036 19292 8046 19348
rect 37874 19292 37884 19348
rect 37940 19292 38892 19348
rect 38948 19292 38958 19348
rect 3938 19180 3948 19236
rect 4004 19180 7756 19236
rect 7812 19180 7822 19236
rect 11218 19180 11228 19236
rect 11284 19180 12236 19236
rect 12292 19180 12302 19236
rect 20290 19180 20300 19236
rect 20356 19180 21644 19236
rect 21700 19180 22428 19236
rect 22484 19180 22494 19236
rect 32722 19180 32732 19236
rect 32788 19180 34188 19236
rect 34244 19180 36540 19236
rect 36596 19180 37772 19236
rect 37828 19180 39116 19236
rect 39172 19180 39182 19236
rect 2034 19068 2044 19124
rect 2100 19068 11452 19124
rect 11508 19068 11518 19124
rect 12562 19068 12572 19124
rect 12628 19068 13468 19124
rect 13524 19068 13534 19124
rect 13794 19068 13804 19124
rect 13860 19068 15820 19124
rect 15876 19068 16716 19124
rect 16772 19068 16782 19124
rect 33954 19068 33964 19124
rect 34020 19068 41916 19124
rect 41972 19068 41982 19124
rect 15026 18956 15036 19012
rect 15092 18956 16828 19012
rect 16884 18956 20748 19012
rect 20804 18956 23548 19012
rect 23604 18956 23614 19012
rect 23874 18956 23884 19012
rect 23940 18956 24556 19012
rect 24612 18956 26012 19012
rect 26068 18956 27692 19012
rect 27748 18956 28588 19012
rect 28644 18956 30044 19012
rect 30100 18956 30110 19012
rect 32834 18956 32844 19012
rect 32900 18956 35644 19012
rect 35700 18956 35710 19012
rect 36082 18956 36092 19012
rect 36148 18956 38780 19012
rect 38836 18956 38846 19012
rect 0 18900 800 18928
rect 23548 18900 23604 18956
rect 0 18844 1708 18900
rect 1764 18844 1774 18900
rect 23548 18844 26460 18900
rect 26516 18844 26526 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 24546 18732 24556 18788
rect 24612 18732 29036 18788
rect 29092 18732 29102 18788
rect 39778 18508 39788 18564
rect 39844 18508 41692 18564
rect 41748 18508 41758 18564
rect 3042 18396 3052 18452
rect 3108 18396 5516 18452
rect 5572 18396 5582 18452
rect 17042 18396 17052 18452
rect 17108 18396 17612 18452
rect 17668 18396 18396 18452
rect 18452 18396 18462 18452
rect 21074 18396 21084 18452
rect 21140 18396 22540 18452
rect 22596 18396 22606 18452
rect 26450 18396 26460 18452
rect 26516 18396 32060 18452
rect 32116 18396 32508 18452
rect 32564 18396 32574 18452
rect 36194 18396 36204 18452
rect 36260 18396 39340 18452
rect 39396 18396 39406 18452
rect 14130 18284 14140 18340
rect 14196 18284 16492 18340
rect 16548 18284 16558 18340
rect 25330 18284 25340 18340
rect 25396 18284 26012 18340
rect 26068 18284 26078 18340
rect 38770 18284 38780 18340
rect 38836 18284 39564 18340
rect 39620 18284 40236 18340
rect 40292 18284 43596 18340
rect 43652 18284 43662 18340
rect 3042 18172 3052 18228
rect 3108 18172 5740 18228
rect 5796 18172 5806 18228
rect 21074 18172 21084 18228
rect 21140 18172 23548 18228
rect 23604 18172 23614 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 27346 17948 27356 18004
rect 27412 17948 29148 18004
rect 29204 17948 29214 18004
rect 26002 17836 26012 17892
rect 26068 17836 31948 17892
rect 32004 17836 32014 17892
rect 3938 17724 3948 17780
rect 4004 17724 4284 17780
rect 4340 17724 4350 17780
rect 20514 17724 20524 17780
rect 20580 17724 21420 17780
rect 21476 17724 21486 17780
rect 35970 17724 35980 17780
rect 36036 17724 41804 17780
rect 41860 17724 41870 17780
rect 28354 17500 28364 17556
rect 28420 17500 29596 17556
rect 29652 17500 29662 17556
rect 32610 17500 32620 17556
rect 32676 17500 42812 17556
rect 42868 17500 42878 17556
rect 6290 17388 6300 17444
rect 6356 17388 11116 17444
rect 11172 17388 11182 17444
rect 18386 17388 18396 17444
rect 18452 17388 20188 17444
rect 20244 17388 20254 17444
rect 32834 17388 32844 17444
rect 32900 17388 35532 17444
rect 35588 17388 35598 17444
rect 36642 17388 36652 17444
rect 36708 17388 42924 17444
rect 42980 17388 42990 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 18050 17052 18060 17108
rect 18116 17052 19852 17108
rect 19908 17052 19918 17108
rect 32162 17052 32172 17108
rect 32228 17052 37212 17108
rect 37268 17052 37278 17108
rect 4722 16940 4732 16996
rect 4788 16940 7196 16996
rect 7252 16940 7262 16996
rect 10882 16940 10892 16996
rect 10948 16940 12348 16996
rect 12404 16940 12414 16996
rect 13906 16940 13916 16996
rect 13972 16940 19516 16996
rect 19572 16940 19582 16996
rect 26338 16940 26348 16996
rect 26404 16940 28364 16996
rect 28420 16940 28430 16996
rect 37090 16940 37100 16996
rect 37156 16940 42924 16996
rect 42980 16940 42990 16996
rect 2258 16828 2268 16884
rect 2324 16828 4060 16884
rect 4116 16828 5068 16884
rect 5124 16828 8876 16884
rect 8932 16828 9436 16884
rect 9492 16828 9502 16884
rect 11330 16828 11340 16884
rect 11396 16828 12684 16884
rect 12740 16828 13244 16884
rect 13300 16828 15372 16884
rect 15428 16828 17052 16884
rect 17108 16828 17118 16884
rect 20850 16828 20860 16884
rect 20916 16828 21308 16884
rect 21364 16828 21756 16884
rect 21812 16828 21822 16884
rect 28242 16828 28252 16884
rect 28308 16828 30044 16884
rect 30100 16828 30110 16884
rect 35308 16828 36988 16884
rect 37044 16828 40348 16884
rect 40404 16828 40414 16884
rect 35308 16772 35364 16828
rect 16818 16716 16828 16772
rect 16884 16716 17836 16772
rect 17892 16716 17902 16772
rect 29026 16716 29036 16772
rect 29092 16716 32508 16772
rect 32564 16716 32574 16772
rect 33170 16716 33180 16772
rect 33236 16716 34972 16772
rect 35028 16716 35364 16772
rect 37538 16716 37548 16772
rect 37604 16716 41916 16772
rect 41972 16716 41982 16772
rect 1586 16604 1596 16660
rect 1652 16604 2380 16660
rect 2436 16604 2446 16660
rect 13122 16604 13132 16660
rect 13188 16604 14140 16660
rect 14196 16604 14206 16660
rect 20962 16604 20972 16660
rect 21028 16604 25116 16660
rect 25172 16604 25182 16660
rect 37650 16604 37660 16660
rect 37716 16604 43932 16660
rect 43988 16604 43998 16660
rect 2706 16492 2716 16548
rect 2772 16492 3500 16548
rect 3556 16492 3566 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 18834 16380 18844 16436
rect 18900 16380 22092 16436
rect 22148 16380 22158 16436
rect 17714 16268 17724 16324
rect 17780 16268 21420 16324
rect 21476 16268 21486 16324
rect 29586 16268 29596 16324
rect 29652 16268 30940 16324
rect 30996 16268 31006 16324
rect 2930 16156 2940 16212
rect 2996 16156 3836 16212
rect 3892 16156 3902 16212
rect 8418 16156 8428 16212
rect 8484 16156 10668 16212
rect 10724 16156 10734 16212
rect 25890 16156 25900 16212
rect 25956 16156 27804 16212
rect 27860 16156 27870 16212
rect 37426 16156 37436 16212
rect 37492 16156 41804 16212
rect 41860 16156 41870 16212
rect 1922 16044 1932 16100
rect 1988 16044 6188 16100
rect 6244 16044 6254 16100
rect 7410 16044 7420 16100
rect 7476 16044 8540 16100
rect 8596 16044 8606 16100
rect 12898 16044 12908 16100
rect 12964 16044 14252 16100
rect 14308 16044 14318 16100
rect 18834 16044 18844 16100
rect 18900 16044 19740 16100
rect 19796 16044 19806 16100
rect 1810 15932 1820 15988
rect 1876 15932 2716 15988
rect 2772 15932 2782 15988
rect 21186 15932 21196 15988
rect 21252 15932 22316 15988
rect 22372 15932 22382 15988
rect 26674 15932 26684 15988
rect 26740 15932 27468 15988
rect 27524 15932 28140 15988
rect 28196 15932 31388 15988
rect 31444 15932 31454 15988
rect 40562 15932 40572 15988
rect 40628 15932 42812 15988
rect 42868 15932 42878 15988
rect 11442 15820 11452 15876
rect 11508 15820 12124 15876
rect 12180 15820 12190 15876
rect 13010 15820 13020 15876
rect 13076 15820 15260 15876
rect 15316 15820 15326 15876
rect 18162 15820 18172 15876
rect 18228 15820 19068 15876
rect 19124 15820 19134 15876
rect 26338 15820 26348 15876
rect 26404 15820 30268 15876
rect 30324 15820 30334 15876
rect 12450 15708 12460 15764
rect 12516 15708 14700 15764
rect 14756 15708 14766 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 29138 15596 29148 15652
rect 29204 15596 31948 15652
rect 32004 15596 32014 15652
rect 16370 15484 16380 15540
rect 16436 15484 17724 15540
rect 17780 15484 17790 15540
rect 21298 15484 21308 15540
rect 21364 15484 22764 15540
rect 22820 15484 23436 15540
rect 23492 15484 25340 15540
rect 25396 15484 27132 15540
rect 27188 15484 27198 15540
rect 31826 15484 31836 15540
rect 31892 15484 33124 15540
rect 33068 15428 33124 15484
rect 8372 15372 10220 15428
rect 10276 15372 11452 15428
rect 11508 15372 11518 15428
rect 24210 15372 24220 15428
rect 24276 15372 25788 15428
rect 25844 15372 25854 15428
rect 26114 15372 26124 15428
rect 26180 15372 26684 15428
rect 26740 15372 26750 15428
rect 30258 15372 30268 15428
rect 30324 15372 31052 15428
rect 31108 15372 31118 15428
rect 31714 15372 31724 15428
rect 31780 15372 31948 15428
rect 33058 15372 33068 15428
rect 33124 15372 33134 15428
rect 38098 15372 38108 15428
rect 38164 15372 38892 15428
rect 38948 15372 38958 15428
rect 41458 15372 41468 15428
rect 41524 15372 42924 15428
rect 42980 15372 42990 15428
rect 8372 15204 8428 15372
rect 31892 15316 31948 15372
rect 9986 15260 9996 15316
rect 10052 15260 11564 15316
rect 11620 15260 11630 15316
rect 31892 15260 33292 15316
rect 33348 15260 33740 15316
rect 33796 15260 33806 15316
rect 6290 15148 6300 15204
rect 6356 15148 8428 15204
rect 14354 15148 14364 15204
rect 14420 15148 15036 15204
rect 15092 15148 15932 15204
rect 15988 15148 17836 15204
rect 17892 15148 18060 15204
rect 18116 15148 21980 15204
rect 22036 15148 22046 15204
rect 26338 15148 26348 15204
rect 26404 15148 27356 15204
rect 27412 15148 27422 15204
rect 30146 15148 30156 15204
rect 30212 15148 33964 15204
rect 34020 15148 34030 15204
rect 34738 15148 34748 15204
rect 34804 15148 36316 15204
rect 36372 15148 38780 15204
rect 38836 15148 39116 15204
rect 39172 15148 39182 15204
rect 40450 15148 40460 15204
rect 40516 15148 42924 15204
rect 42980 15148 42990 15204
rect 5730 15036 5740 15092
rect 5796 15036 8428 15092
rect 8484 15036 8494 15092
rect 40002 15036 40012 15092
rect 40068 15036 41804 15092
rect 41860 15036 41870 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 36866 14812 36876 14868
rect 36932 14812 38220 14868
rect 38276 14812 38286 14868
rect 16594 14700 16604 14756
rect 16660 14700 17948 14756
rect 18004 14700 18014 14756
rect 12450 14588 12460 14644
rect 12516 14588 14028 14644
rect 14084 14588 14094 14644
rect 29698 14588 29708 14644
rect 29764 14588 34300 14644
rect 34356 14588 34366 14644
rect 21634 14476 21644 14532
rect 21700 14476 21980 14532
rect 22036 14476 22046 14532
rect 30818 14476 30828 14532
rect 30884 14476 31948 14532
rect 31892 14420 31948 14476
rect 16706 14364 16716 14420
rect 16772 14364 18508 14420
rect 18564 14364 18574 14420
rect 31892 14364 35308 14420
rect 35364 14364 35374 14420
rect 37650 14364 37660 14420
rect 37716 14364 44044 14420
rect 44100 14364 44110 14420
rect 33506 14252 33516 14308
rect 33572 14252 34300 14308
rect 34356 14252 34366 14308
rect 36530 14252 36540 14308
rect 36596 14252 39004 14308
rect 39060 14252 39070 14308
rect 2706 14140 2716 14196
rect 2772 14140 3612 14196
rect 3668 14140 3678 14196
rect 35634 14140 35644 14196
rect 35700 14140 37996 14196
rect 38052 14140 38062 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 23314 14028 23324 14084
rect 23380 14028 26124 14084
rect 26180 14028 26190 14084
rect 38658 13916 38668 13972
rect 38724 13916 42028 13972
rect 42084 13916 42094 13972
rect 11666 13580 11676 13636
rect 11732 13580 12460 13636
rect 12516 13580 12526 13636
rect 22978 13580 22988 13636
rect 23044 13580 24108 13636
rect 24164 13580 24174 13636
rect 24770 13580 24780 13636
rect 24836 13580 27244 13636
rect 27300 13580 27310 13636
rect 4946 13468 4956 13524
rect 5012 13468 5964 13524
rect 6020 13468 6030 13524
rect 32722 13468 32732 13524
rect 32788 13468 35420 13524
rect 35476 13468 35486 13524
rect 23314 13356 23324 13412
rect 23380 13356 26572 13412
rect 26628 13356 26638 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 10098 13020 10108 13076
rect 10164 13020 15260 13076
rect 15316 13020 15326 13076
rect 40002 13020 40012 13076
rect 40068 13020 40796 13076
rect 40852 13020 40862 13076
rect 26898 12796 26908 12852
rect 26964 12796 31164 12852
rect 31220 12796 31230 12852
rect 28018 12684 28028 12740
rect 28084 12684 29372 12740
rect 29428 12684 29438 12740
rect 34850 12684 34860 12740
rect 34916 12684 36876 12740
rect 36932 12684 36942 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 25666 12012 25676 12068
rect 25732 12012 29036 12068
rect 29092 12012 29102 12068
rect 32498 12012 32508 12068
rect 32564 12012 34076 12068
rect 34132 12012 34142 12068
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 21746 11452 21756 11508
rect 21812 11452 26684 11508
rect 26740 11452 26750 11508
rect 27794 11452 27804 11508
rect 27860 11452 33516 11508
rect 33572 11452 33582 11508
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 43586 8876 43596 8932
rect 43652 8820 43708 8932
rect 45200 8820 46000 8848
rect 43652 8764 44156 8820
rect 44212 8764 46000 8820
rect 45200 8736 46000 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 45200 8148 46000 8176
rect 44034 8092 44044 8148
rect 44100 8092 46000 8148
rect 45200 8064 46000 8092
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 45200 7476 46000 7504
rect 44034 7420 44044 7476
rect 44100 7420 46000 7476
rect 45200 7392 46000 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 45200 6804 46000 6832
rect 42578 6748 42588 6804
rect 42644 6748 46000 6804
rect 45200 6720 46000 6748
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 45200 6132 46000 6160
rect 44034 6076 44044 6132
rect 44100 6076 46000 6132
rect 45200 6048 46000 6076
rect 41794 5852 41804 5908
rect 41860 5852 42924 5908
rect 42980 5852 42990 5908
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 45200 5460 46000 5488
rect 44034 5404 44044 5460
rect 44100 5404 46000 5460
rect 45200 5376 46000 5404
rect 35746 5180 35756 5236
rect 35812 5180 37884 5236
rect 37940 5180 37950 5236
rect 36418 5068 36428 5124
rect 36484 5068 38108 5124
rect 38164 5068 38174 5124
rect 39218 4956 39228 5012
rect 39284 4956 40908 5012
rect 40964 4956 40974 5012
rect 42242 4844 42252 4900
rect 42308 4844 44156 4900
rect 44212 4844 44222 4900
rect 45200 4788 46000 4816
rect 43026 4732 43036 4788
rect 43092 4732 46000 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 45200 4704 46000 4732
rect 43138 4620 43148 4676
rect 43204 4620 43820 4676
rect 43876 4620 43886 4676
rect 41458 4508 41468 4564
rect 41524 4508 43036 4564
rect 43092 4508 43102 4564
rect 37986 4396 37996 4452
rect 38052 4396 41580 4452
rect 41636 4396 41646 4452
rect 24882 4284 24892 4340
rect 24948 4284 25564 4340
rect 25620 4284 25630 4340
rect 42690 4284 42700 4340
rect 42756 4284 44044 4340
rect 44100 4284 44380 4340
rect 44436 4284 44446 4340
rect 19506 4172 19516 4228
rect 19572 4172 20188 4228
rect 26226 4172 26236 4228
rect 26292 4172 27356 4228
rect 27412 4172 27422 4228
rect 32162 4172 32172 4228
rect 32228 4172 32956 4228
rect 33012 4172 33022 4228
rect 37650 4172 37660 4228
rect 37716 4172 38556 4228
rect 38612 4172 38622 4228
rect 42130 4172 42140 4228
rect 42196 4172 43820 4228
rect 43876 4172 43886 4228
rect 20132 4060 20188 4172
rect 45200 4116 46000 4144
rect 20244 4060 20254 4116
rect 42354 4060 42364 4116
rect 42420 4060 46000 4116
rect 45200 4032 46000 4060
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 25554 3612 25564 3668
rect 25620 3612 26572 3668
rect 26628 3612 26638 3668
rect 27570 3612 27580 3668
rect 27636 3612 28812 3668
rect 28868 3612 28878 3668
rect 31602 3612 31612 3668
rect 31668 3612 32620 3668
rect 32676 3612 32686 3668
rect 38994 3612 39004 3668
rect 39060 3612 40236 3668
rect 40292 3612 40302 3668
rect 34962 3500 34972 3556
rect 35028 3500 36092 3556
rect 36148 3500 36158 3556
rect 38210 3500 38220 3556
rect 38276 3500 39788 3556
rect 39844 3500 39854 3556
rect 45200 3444 46000 3472
rect 39554 3388 39564 3444
rect 39620 3388 41804 3444
rect 41860 3388 41870 3444
rect 44146 3388 44156 3444
rect 44212 3388 46000 3444
rect 45200 3360 46000 3388
rect 21522 3276 21532 3332
rect 21588 3276 22652 3332
rect 22708 3276 22718 3332
rect 23650 3276 23660 3332
rect 23716 3276 24556 3332
rect 24612 3276 24622 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 45200 2772 46000 2800
rect 43138 2716 43148 2772
rect 43204 2716 46000 2772
rect 45200 2688 46000 2716
rect 45200 2100 46000 2128
rect 44370 2044 44380 2100
rect 44436 2044 46000 2100
rect 45200 2016 46000 2044
rect 45200 0 46000 112
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 31948 23772 32004 23828
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 31948 20748 32004 20804
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 31948 23828 32004 23838
rect 31948 20804 32004 23772
rect 31948 20738 32004 20748
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _123_
timestamp 1698431365
transform -1 0 18816 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _125_
timestamp 1698431365
transform -1 0 15680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _126_
timestamp 1698431365
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _127_
timestamp 1698431365
transform -1 0 9184 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _128_
timestamp 1698431365
transform 1 0 6496 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _129_
timestamp 1698431365
transform 1 0 4592 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _130_
timestamp 1698431365
transform -1 0 3920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _131_
timestamp 1698431365
transform 1 0 2576 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _132_
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _133_
timestamp 1698431365
transform 1 0 10864 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _134_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _135_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _136_
timestamp 1698431365
transform -1 0 12432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _137_
timestamp 1698431365
transform 1 0 9744 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _138_
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _139_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _140_
timestamp 1698431365
transform -1 0 6944 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _141_
timestamp 1698431365
transform 1 0 13664 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _142_
timestamp 1698431365
transform 1 0 14336 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _143_
timestamp 1698431365
transform 1 0 10528 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _144_
timestamp 1698431365
transform -1 0 10080 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _145_
timestamp 1698431365
transform 1 0 21392 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _146_
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _147_
timestamp 1698431365
transform -1 0 20160 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _148_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _149_
timestamp 1698431365
transform 1 0 20272 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _150_
timestamp 1698431365
transform -1 0 21840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _151_
timestamp 1698431365
transform -1 0 20720 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _152_
timestamp 1698431365
transform 1 0 17584 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _153_
timestamp 1698431365
transform -1 0 17024 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _154_
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _155_
timestamp 1698431365
transform -1 0 23520 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _156_
timestamp 1698431365
transform 1 0 34608 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _157_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _158_
timestamp 1698431365
transform 1 0 31360 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _159_
timestamp 1698431365
transform -1 0 29680 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _160_
timestamp 1698431365
transform -1 0 28224 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _161_
timestamp 1698431365
transform 1 0 35504 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _162_
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _163_
timestamp 1698431365
transform 1 0 31248 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _164_
timestamp 1698431365
transform 1 0 29120 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _165_
timestamp 1698431365
transform 1 0 27776 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _166_
timestamp 1698431365
transform -1 0 28112 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _167_
timestamp 1698431365
transform -1 0 26656 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _168_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _169_
timestamp 1698431365
transform -1 0 25760 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _170_
timestamp 1698431365
transform -1 0 22288 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _171_
timestamp 1698431365
transform -1 0 22624 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _172_
timestamp 1698431365
transform -1 0 21840 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _173_
timestamp 1698431365
transform -1 0 19600 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _174_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _175_
timestamp 1698431365
transform -1 0 24080 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _176_
timestamp 1698431365
transform -1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _177_
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _178_
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _179_
timestamp 1698431365
transform 1 0 29120 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _180_
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _181_
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _182_
timestamp 1698431365
transform -1 0 33600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _183_
timestamp 1698431365
transform -1 0 32704 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _184_
timestamp 1698431365
transform -1 0 32032 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _185_
timestamp 1698431365
transform -1 0 31360 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _186_
timestamp 1698431365
transform -1 0 28672 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _187_
timestamp 1698431365
transform 1 0 43568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _188_
timestamp 1698431365
transform 1 0 43456 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _189_
timestamp 1698431365
transform 1 0 34496 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _190_
timestamp 1698431365
transform 1 0 43568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _191_
timestamp 1698431365
transform 1 0 39312 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _192_
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _193_
timestamp 1698431365
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _194_
timestamp 1698431365
transform -1 0 42560 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _195_
timestamp 1698431365
transform 1 0 43456 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _196_
timestamp 1698431365
transform 1 0 43568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _197_
timestamp 1698431365
transform 1 0 39536 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _198_
timestamp 1698431365
transform 1 0 38864 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _199_
timestamp 1698431365
transform -1 0 37520 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _200_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _201_
timestamp 1698431365
transform 1 0 43456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _202_
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _203_
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _204_
timestamp 1698431365
transform -1 0 39872 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _205_
timestamp 1698431365
transform -1 0 39088 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _206_
timestamp 1698431365
transform -1 0 39312 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _207_
timestamp 1698431365
transform 1 0 43568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _208_
timestamp 1698431365
transform -1 0 39424 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _209_
timestamp 1698431365
transform -1 0 36624 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _210_
timestamp 1698431365
transform -1 0 34944 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _211_
timestamp 1698431365
transform 1 0 27216 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _212_
timestamp 1698431365
transform -1 0 33600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _213_
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _214_
timestamp 1698431365
transform -1 0 27104 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _215_
timestamp 1698431365
transform -1 0 26992 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _216_
timestamp 1698431365
transform -1 0 26320 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _217_
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _218_
timestamp 1698431365
transform 1 0 31584 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _219_
timestamp 1698431365
transform -1 0 31584 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _220_
timestamp 1698431365
transform -1 0 28336 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _221_
timestamp 1698431365
transform -1 0 27664 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _222_
timestamp 1698431365
transform -1 0 16576 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _223_
timestamp 1698431365
transform -1 0 18032 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _224_
timestamp 1698431365
transform -1 0 18256 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _225_
timestamp 1698431365
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _226_
timestamp 1698431365
transform -1 0 21840 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _227_
timestamp 1698431365
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _228_
timestamp 1698431365
transform 1 0 21840 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _229_
timestamp 1698431365
transform -1 0 15232 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _230_
timestamp 1698431365
transform -1 0 14560 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _231_
timestamp 1698431365
transform -1 0 17024 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _232_
timestamp 1698431365
transform -1 0 16128 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _233_
timestamp 1698431365
transform 1 0 11424 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _234_
timestamp 1698431365
transform -1 0 11648 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _235_
timestamp 1698431365
transform -1 0 7168 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _236_
timestamp 1698431365
transform -1 0 10416 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _237_
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _238_
timestamp 1698431365
transform -1 0 6496 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _239_
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _240_
timestamp 1698431365
transform 1 0 1792 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _241_
timestamp 1698431365
transform 1 0 3136 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _242_
timestamp 1698431365
transform 1 0 5824 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _243_
timestamp 1698431365
transform -1 0 6160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _244_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _245_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _246_
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _247_
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _248_
timestamp 1698431365
transform 1 0 3920 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _249_
timestamp 1698431365
transform -1 0 6048 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _250_
timestamp 1698431365
transform -1 0 5824 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _251_
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _252_
timestamp 1698431365
transform 1 0 13216 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _253_
timestamp 1698431365
transform -1 0 17136 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _254_
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _255_
timestamp 1698431365
transform -1 0 13216 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _256_
timestamp 1698431365
transform 1 0 7952 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _257_
timestamp 1698431365
transform -1 0 10752 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _258_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _259_
timestamp 1698431365
transform -1 0 9184 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _260_
timestamp 1698431365
transform 1 0 11536 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _261_
timestamp 1698431365
transform 1 0 9296 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _262_
timestamp 1698431365
transform 1 0 7840 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _263_
timestamp 1698431365
transform -1 0 9296 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _264_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _265_
timestamp 1698431365
transform 1 0 16128 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _266_
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _267_
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _268_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _269_
timestamp 1698431365
transform -1 0 20048 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _270_
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _271_
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _272_
timestamp 1698431365
transform 1 0 21056 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _273_
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _274_
timestamp 1698431365
transform -1 0 36736 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _275_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _276_
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _277_
timestamp 1698431365
transform 1 0 23968 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _278_
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _279_
timestamp 1698431365
transform 1 0 30464 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _280_
timestamp 1698431365
transform 1 0 28896 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _281_
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _282_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _283_
timestamp 1698431365
transform 1 0 23632 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _284_
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _285_
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _286_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _287_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _288_
timestamp 1698431365
transform 1 0 17136 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _289_
timestamp 1698431365
transform 1 0 13216 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _290_
timestamp 1698431365
transform -1 0 26096 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _291_
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _292_
timestamp 1698431365
transform 1 0 18256 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _293_
timestamp 1698431365
transform -1 0 20384 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _294_
timestamp 1698431365
transform -1 0 32816 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _295_
timestamp 1698431365
transform 1 0 25872 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _296_
timestamp 1698431365
transform -1 0 36736 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _297_
timestamp 1698431365
transform 1 0 29792 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _298_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _299_
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _300_
timestamp 1698431365
transform 1 0 25760 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _301_
timestamp 1698431365
transform 1 0 24528 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _302_
timestamp 1698431365
transform 1 0 39088 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _303_
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _304_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _305_
timestamp 1698431365
transform 1 0 36736 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _306_
timestamp 1698431365
transform 1 0 34160 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _307_
timestamp 1698431365
transform 1 0 32816 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _308_
timestamp 1698431365
transform 1 0 38080 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _309_
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _310_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _311_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _312_
timestamp 1698431365
transform 1 0 36736 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _313_
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _314_
timestamp 1698431365
transform -1 0 40656 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _315_
timestamp 1698431365
transform 1 0 36736 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _316_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _317_
timestamp 1698431365
transform 1 0 33264 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _318_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _319_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _320_
timestamp 1698431365
transform -1 0 40656 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _321_
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _322_
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _323_
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _324_
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _325_
timestamp 1698431365
transform -1 0 32816 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _326_
timestamp 1698431365
transform -1 0 26320 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _327_
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _328_
timestamp 1698431365
transform 1 0 21056 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _329_
timestamp 1698431365
transform -1 0 33152 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _330_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _331_
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _332_
timestamp 1698431365
transform -1 0 28896 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _333_
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _334_
timestamp 1698431365
transform -1 0 20496 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _335_
timestamp 1698431365
transform 1 0 13216 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _336_
timestamp 1698431365
transform 1 0 17360 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _337_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _338_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _339_
timestamp 1698431365
transform -1 0 21840 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _340_
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _341_
timestamp 1698431365
transform -1 0 15456 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _342_
timestamp 1698431365
transform -1 0 17136 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _343_
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _344_
timestamp 1698431365
transform -1 0 9296 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _345_
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _346_
timestamp 1698431365
transform -1 0 11424 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _347_
timestamp 1698431365
transform 1 0 7168 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _348_
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _349_
timestamp 1698431365
transform -1 0 5376 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _350_
timestamp 1698431365
transform -1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _351_
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _352_
timestamp 1698431365
transform 1 0 3808 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _353_
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _379_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_
timestamp 1698431365
transform -1 0 39984 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1698431365
transform 1 0 38976 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _382_
timestamp 1698431365
transform 1 0 42000 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1698431365
transform 1 0 24304 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _384_
timestamp 1698431365
transform 1 0 19264 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1698431365
transform 1 0 39088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1698431365
transform 1 0 42224 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1698431365
transform -1 0 37744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1698431365
transform 1 0 42112 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _391_
timestamp 1698431365
transform 1 0 19600 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1698431365
transform -1 0 43008 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _393_
timestamp 1698431365
transform 1 0 14672 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1698431365
transform 1 0 31696 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _395_
timestamp 1698431365
transform 1 0 33152 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1698431365
transform 1 0 20272 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1698431365
transform 1 0 38416 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1698431365
transform 1 0 24864 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1698431365
transform 1 0 41328 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _400_
timestamp 1698431365
transform 1 0 15344 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1698431365
transform 1 0 18368 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _402_
timestamp 1698431365
transform 1 0 38640 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _403_
timestamp 1698431365
transform -1 0 38416 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _406_
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _408_
timestamp 1698431365
transform -1 0 43344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1698431365
transform -1 0 44016 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _412_
timestamp 1698431365
transform 1 0 39648 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1698431365
transform 1 0 41664 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__I
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1698431365
transform 1 0 15456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1698431365
transform 1 0 16352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1698431365
transform 1 0 8288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__I
timestamp 1698431365
transform 1 0 7392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1698431365
transform 1 0 5712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__I
timestamp 1698431365
transform -1 0 2576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1698431365
transform -1 0 12656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I
timestamp 1698431365
transform -1 0 21056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__I
timestamp 1698431365
transform 1 0 24304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1698431365
transform -1 0 29456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1698431365
transform -1 0 32816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1698431365
transform 1 0 34272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1698431365
transform 1 0 33824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1698431365
transform 1 0 31024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1698431365
transform -1 0 28000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I
timestamp 1698431365
transform -1 0 42560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1698431365
transform 1 0 41440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1698431365
transform 1 0 37296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I
timestamp 1698431365
transform -1 0 26992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1698431365
transform 1 0 15792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__CLK
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__CLK
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__CLK
timestamp 1698431365
transform -1 0 30128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__CLK
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__CLK
timestamp 1698431365
transform -1 0 30576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__CLK
timestamp 1698431365
transform -1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__CLK
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__CLK
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__CLK
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__CLK
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__CLK
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__CLK
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_prog_clk_I
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_prog_clk_I
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_prog_clk_I
timestamp 1698431365
transform -1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_prog_clk_I
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_prog_clk_I
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_prog_clk_I
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_prog_clk_I
timestamp 1698431365
transform 1 0 26768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_prog_clk_I
timestamp 1698431365
transform 1 0 32144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 42784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 14336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 37744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 20272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 32256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 31024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 19600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 26320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 43680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 35952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 16912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 15232 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 23632 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 40768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 19936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 42336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 43232 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 37296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 24976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 44128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 19152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 41216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 43904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 43680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 43232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 40768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 32592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1698431365
transform -1 0 22848 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1698431365
transform -1 0 32256 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1698431365
transform -1 0 32592 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1698431365
transform 1 0 33264 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_154 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_216
timestamp 1698431365
transform 1 0 25536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_230 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_250
timestamp 1698431365
transform 1 0 29344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_258
timestamp 1698431365
transform 1 0 30240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_262
timestamp 1698431365
transform 1 0 30688 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_284
timestamp 1698431365
transform 1 0 33152 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_288
timestamp 1698431365
transform 1 0 33600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_299
timestamp 1698431365
transform 1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_326
timestamp 1698431365
transform 1 0 37856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_352
timestamp 1698431365
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_358
timestamp 1698431365
transform 1 0 41440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_370
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_159
timestamp 1698431365
transform 1 0 19152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_175
timestamp 1698431365
transform 1 0 20944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_191
timestamp 1698431365
transform 1 0 22736 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_199
timestamp 1698431365
transform 1 0 23632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_227
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_235
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_267
timestamp 1698431365
transform 1 0 31248 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_271
timestamp 1698431365
transform 1 0 31696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_273
timestamp 1698431365
transform 1 0 31920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_289
timestamp 1698431365
transform 1 0 33712 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_297
timestamp 1698431365
transform 1 0 34608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_321
timestamp 1698431365
transform 1 0 37296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_337
timestamp 1698431365
transform 1 0 39088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_341
timestamp 1698431365
transform 1 0 39536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_209
timestamp 1698431365
transform 1 0 24752 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_216
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_232
timestamp 1698431365
transform 1 0 27328 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_240
timestamp 1698431365
transform 1 0 28224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_263
timestamp 1698431365
transform 1 0 30800 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_277
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_281
timestamp 1698431365
transform 1 0 32816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_283
timestamp 1698431365
transform 1 0 33040 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_290
timestamp 1698431365
transform 1 0 33824 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_306
timestamp 1698431365
transform 1 0 35616 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_309
timestamp 1698431365
transform 1 0 35952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_343
timestamp 1698431365
transform 1 0 39760 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_347
timestamp 1698431365
transform 1 0 40208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_349
timestamp 1698431365
transform 1 0 40432 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_352
timestamp 1698431365
transform 1 0 40768 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_356
timestamp 1698431365
transform 1 0 41216 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_360
timestamp 1698431365
transform 1 0 41664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_366
timestamp 1698431365
transform 1 0 42336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_193
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_201
timestamp 1698431365
transform 1 0 23856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_211
timestamp 1698431365
transform 1 0 24976 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_349
timestamp 1698431365
transform 1 0 40432 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_365
timestamp 1698431365
transform 1 0 42224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_369
timestamp 1698431365
transform 1 0 42672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_360
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_364
timestamp 1698431365
transform 1 0 42112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_225
timestamp 1698431365
transform 1 0 26544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_233
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_349
timestamp 1698431365
transform 1 0 40432 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_365
timestamp 1698431365
transform 1 0 42224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_369
timestamp 1698431365
transform 1 0 42672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_162
timestamp 1698431365
transform 1 0 19488 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_169
timestamp 1698431365
transform 1 0 20272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_176
timestamp 1698431365
transform 1 0 21056 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_368
timestamp 1698431365
transform 1 0 42560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_189
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_207
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_223
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_279
timestamp 1698431365
transform 1 0 32592 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_283
timestamp 1698431365
transform 1 0 33040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_285
timestamp 1698431365
transform 1 0 33264 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_302
timestamp 1698431365
transform 1 0 35168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_112
timestamp 1698431365
transform 1 0 13888 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_129
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_137
timestamp 1698431365
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_182
timestamp 1698431365
transform 1 0 21728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_202
timestamp 1698431365
transform 1 0 23968 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_237
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_245
timestamp 1698431365
transform 1 0 28784 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_262
timestamp 1698431365
transform 1 0 30688 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_307
timestamp 1698431365
transform 1 0 35728 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_339
timestamp 1698431365
transform 1 0 39312 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698431365
transform 1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_161
timestamp 1698431365
transform 1 0 19376 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_169
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_223
timestamp 1698431365
transform 1 0 26320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_272
timestamp 1698431365
transform 1 0 31808 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_288
timestamp 1698431365
transform 1 0 33600 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_292
timestamp 1698431365
transform 1 0 34048 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_309
timestamp 1698431365
transform 1 0 35952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_342
timestamp 1698431365
transform 1 0 39648 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_350
timestamp 1698431365
transform 1 0 40544 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_367
timestamp 1698431365
transform 1 0 42448 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_42
timestamp 1698431365
transform 1 0 6048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_50
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_88
timestamp 1698431365
transform 1 0 11200 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_105
timestamp 1698431365
transform 1 0 13104 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_113
timestamp 1698431365
transform 1 0 14000 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_130
timestamp 1698431365
transform 1 0 15904 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_162
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_236
timestamp 1698431365
transform 1 0 27776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_254
timestamp 1698431365
transform 1 0 29792 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_262
timestamp 1698431365
transform 1 0 30688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_310
timestamp 1698431365
transform 1 0 36064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_318
timestamp 1698431365
transform 1 0 36960 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_335
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_6
timestamp 1698431365
transform 1 0 2016 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_23
timestamp 1698431365
transform 1 0 3920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_39
timestamp 1698431365
transform 1 0 5712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_56
timestamp 1698431365
transform 1 0 7616 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_88
timestamp 1698431365
transform 1 0 11200 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_124
timestamp 1698431365
transform 1 0 15232 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_141
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_149
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_166
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_191
timestamp 1698431365
transform 1 0 22736 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_229
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_249
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_284
timestamp 1698431365
transform 1 0 33152 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_292
timestamp 1698431365
transform 1 0 34048 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_351
timestamp 1698431365
transform 1 0 40656 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_359
timestamp 1698431365
transform 1 0 41552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_376
timestamp 1698431365
transform 1 0 43456 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_40
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_48
timestamp 1698431365
transform 1 0 6720 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_74
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_81
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_85
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_132
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_144
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_151
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_159
timestamp 1698431365
transform 1 0 19152 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_229
timestamp 1698431365
transform 1 0 26992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_340
timestamp 1698431365
transform 1 0 39424 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_348
timestamp 1698431365
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_360
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_377
timestamp 1698431365
transform 1 0 43568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_381
timestamp 1698431365
transform 1 0 44016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_383
timestamp 1698431365
transform 1 0 44240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_39
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_46
timestamp 1698431365
transform 1 0 6496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_54
timestamp 1698431365
transform 1 0 7392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_128
timestamp 1698431365
transform 1 0 15680 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_136
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_189
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_224
timestamp 1698431365
transform 1 0 26432 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_226
timestamp 1698431365
transform 1 0 26656 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_351
timestamp 1698431365
transform 1 0 40656 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_359
timestamp 1698431365
transform 1 0 41552 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_376
timestamp 1698431365
transform 1 0 43456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_183
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_383
timestamp 1698431365
transform 1 0 44240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_183
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_221
timestamp 1698431365
transform 1 0 26096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_223
timestamp 1698431365
transform 1 0 26320 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_351
timestamp 1698431365
transform 1 0 40656 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_359
timestamp 1698431365
transform 1 0 41552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_382
timestamp 1698431365
transform 1 0 44128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_44
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_61
timestamp 1698431365
transform 1 0 8176 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_90
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_98
timestamp 1698431365
transform 1 0 12320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_133
timestamp 1698431365
transform 1 0 16240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_193
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_377
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_381
timestamp 1698431365
transform 1 0 44016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_383
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_39
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_86
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_88
timestamp 1698431365
transform 1 0 11200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_190
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_198
timestamp 1698431365
transform 1 0 23520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_233
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_237
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_371
timestamp 1698431365
transform 1 0 42896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_379
timestamp 1698431365
transform 1 0 43792 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_10
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_14
timestamp 1698431365
transform 1 0 2912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_56
timestamp 1698431365
transform 1 0 7616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_253
timestamp 1698431365
transform 1 0 29680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_257
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_261
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_284
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_319
timestamp 1698431365
transform 1 0 37072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_323
timestamp 1698431365
transform 1 0 37520 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_327
timestamp 1698431365
transform 1 0 37968 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_344
timestamp 1698431365
transform 1 0 39872 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_348
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_360
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_377
timestamp 1698431365
transform 1 0 43568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_381
timestamp 1698431365
transform 1 0 44016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_383
timestamp 1698431365
transform 1 0 44240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_43
timestamp 1698431365
transform 1 0 6160 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_51
timestamp 1698431365
transform 1 0 7056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_221
timestamp 1698431365
transform 1 0 26096 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_237
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_272
timestamp 1698431365
transform 1 0 31808 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_280
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_323
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_359
timestamp 1698431365
transform 1 0 41552 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_363
timestamp 1698431365
transform 1 0 42000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_365
timestamp 1698431365
transform 1 0 42224 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_74
timestamp 1698431365
transform 1 0 9632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_97
timestamp 1698431365
transform 1 0 12208 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_101
timestamp 1698431365
transform 1 0 12656 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_105
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_201
timestamp 1698431365
transform 1 0 23856 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_252
timestamp 1698431365
transform 1 0 29568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_256
timestamp 1698431365
transform 1 0 30016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_260
timestamp 1698431365
transform 1 0 30464 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_288
timestamp 1698431365
transform 1 0 33600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_292
timestamp 1698431365
transform 1 0 34048 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_345
timestamp 1698431365
transform 1 0 39984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_383
timestamp 1698431365
transform 1 0 44240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_127
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_170
timestamp 1698431365
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_235
timestamp 1698431365
transform 1 0 27664 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_288
timestamp 1698431365
transform 1 0 33600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_292
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_296
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_313
timestamp 1698431365
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_351
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_355
timestamp 1698431365
transform 1 0 41104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_357
timestamp 1698431365
transform 1 0 41328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_382
timestamp 1698431365
transform 1 0 44128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_36
timestamp 1698431365
transform 1 0 5376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_61
timestamp 1698431365
transform 1 0 8176 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_160
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_383
timestamp 1698431365
transform 1 0 44240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_84
timestamp 1698431365
transform 1 0 10752 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_115
timestamp 1698431365
transform 1 0 14224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_132
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_136
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_198
timestamp 1698431365
transform 1 0 23520 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_202
timestamp 1698431365
transform 1 0 23968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_204
timestamp 1698431365
transform 1 0 24192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_323
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_327
timestamp 1698431365
transform 1 0 37968 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_368
timestamp 1698431365
transform 1 0 42560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_380
timestamp 1698431365
transform 1 0 43904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_40
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_44
timestamp 1698431365
transform 1 0 6272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_61
timestamp 1698431365
transform 1 0 8176 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_156
timestamp 1698431365
transform 1 0 18816 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_258
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_264
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_273
timestamp 1698431365
transform 1 0 31920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_284
timestamp 1698431365
transform 1 0 33152 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_377
timestamp 1698431365
transform 1 0 43568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_381
timestamp 1698431365
transform 1 0 44016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_383
timestamp 1698431365
transform 1 0 44240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_30
timestamp 1698431365
transform 1 0 4704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_128
timestamp 1698431365
transform 1 0 15680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_207
timestamp 1698431365
transform 1 0 24528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698431365
transform 1 0 25424 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_232
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_272
timestamp 1698431365
transform 1 0 31808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_274
timestamp 1698431365
transform 1 0 32032 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_277
timestamp 1698431365
transform 1 0 32368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_357
timestamp 1698431365
transform 1 0 41328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_365
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_6
timestamp 1698431365
transform 1 0 2016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_57
timestamp 1698431365
transform 1 0 7728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_61
timestamp 1698431365
transform 1 0 8176 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_198
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_224
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_324
timestamp 1698431365
transform 1 0 37632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_332
timestamp 1698431365
transform 1 0 38528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_383
timestamp 1698431365
transform 1 0 44240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_6
timestamp 1698431365
transform 1 0 2016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_109
timestamp 1698431365
transform 1 0 13552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_122
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_168
timestamp 1698431365
transform 1 0 20160 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698431365
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_254
timestamp 1698431365
transform 1 0 29792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_258
timestamp 1698431365
transform 1 0 30240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_294
timestamp 1698431365
transform 1 0 34272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_310
timestamp 1698431365
transform 1 0 36064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_351
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_359
timestamp 1698431365
transform 1 0 41552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_42
timestamp 1698431365
transform 1 0 6048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_44
timestamp 1698431365
transform 1 0 6272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_61
timestamp 1698431365
transform 1 0 8176 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_88
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_90
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_129
timestamp 1698431365
transform 1 0 15792 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_167
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698431365
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_173
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_360
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_377
timestamp 1698431365
transform 1 0 43568 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_381
timestamp 1698431365
transform 1 0 44016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_383
timestamp 1698431365
transform 1 0 44240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_18
timestamp 1698431365
transform 1 0 3360 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_26
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_52
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_56
timestamp 1698431365
transform 1 0 7616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_92
timestamp 1698431365
transform 1 0 11648 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_100
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_124
timestamp 1698431365
transform 1 0 15232 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_132
timestamp 1698431365
transform 1 0 16128 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_167
timestamp 1698431365
transform 1 0 20048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_351
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_359
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_376
timestamp 1698431365
transform 1 0 43456 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_36
timestamp 1698431365
transform 1 0 5376 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_52
timestamp 1698431365
transform 1 0 7168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_98
timestamp 1698431365
transform 1 0 12320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_115
timestamp 1698431365
transform 1 0 14224 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_123
timestamp 1698431365
transform 1 0 15120 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_256
timestamp 1698431365
transform 1 0 30016 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_264
timestamp 1698431365
transform 1 0 30912 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_274
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_307
timestamp 1698431365
transform 1 0 35728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_315
timestamp 1698431365
transform 1 0 36624 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_332
timestamp 1698431365
transform 1 0 38528 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_348
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_62
timestamp 1698431365
transform 1 0 8288 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_70
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_90
timestamp 1698431365
transform 1 0 11424 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_98
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_102
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_149
timestamp 1698431365
transform 1 0 18032 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_157
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_217
timestamp 1698431365
transform 1 0 25648 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_240
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_253
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_261
timestamp 1698431365
transform 1 0 30576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_263
timestamp 1698431365
transform 1 0 30800 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_288
timestamp 1698431365
transform 1 0 33600 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_342
timestamp 1698431365
transform 1 0 39648 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_374
timestamp 1698431365
transform 1 0 43232 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_88
timestamp 1698431365
transform 1 0 11200 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_96
timestamp 1698431365
transform 1 0 12096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_100
timestamp 1698431365
transform 1 0 12544 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_117
timestamp 1698431365
transform 1 0 14448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_133
timestamp 1698431365
transform 1 0 16240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_158
timestamp 1698431365
transform 1 0 19040 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_162
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_205
timestamp 1698431365
transform 1 0 24304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_232
timestamp 1698431365
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_250
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_258
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_275
timestamp 1698431365
transform 1 0 32144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_311
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_343
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_364
timestamp 1698431365
transform 1 0 42112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_371
timestamp 1698431365
transform 1 0 42896 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_375
timestamp 1698431365
transform 1 0 43344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_139
timestamp 1698431365
transform 1 0 16912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_157
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_202
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_234
timestamp 1698431365
transform 1 0 27552 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_242
timestamp 1698431365
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_349
timestamp 1698431365
transform 1 0 40432 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_365
timestamp 1698431365
transform 1 0 42224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_369
timestamp 1698431365
transform 1 0 42672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_166
timestamp 1698431365
transform 1 0 19936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_168
timestamp 1698431365
transform 1 0 20160 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_175
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_183
timestamp 1698431365
transform 1 0 21840 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_199
timestamp 1698431365
transform 1 0 23632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_226
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_258
timestamp 1698431365
transform 1 0 30240 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_274
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_278
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_368
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_376
timestamp 1698431365
transform 1 0 43456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_349
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_365
timestamp 1698431365
transform 1 0 42224 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_373
timestamp 1698431365
transform 1 0 43120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_375
timestamp 1698431365
transform 1 0 43344 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_376
timestamp 1698431365
transform 1 0 43456 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_365
timestamp 1698431365
transform 1 0 42224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_369
timestamp 1698431365
transform 1 0 42672 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_371
timestamp 1698431365
transform 1 0 42896 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_360
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_139
timestamp 1698431365
transform 1 0 16912 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_155
timestamp 1698431365
transform 1 0 18704 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_163
timestamp 1698431365
transform 1 0 19600 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_166
timestamp 1698431365
transform 1 0 19936 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_335
timestamp 1698431365
transform 1 0 38864 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_348
timestamp 1698431365
transform 1 0 40320 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_352
timestamp 1698431365
transform 1 0 40768 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_372
timestamp 1698431365
transform 1 0 43008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_104
timestamp 1698431365
transform 1 0 12992 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_112
timestamp 1698431365
transform 1 0 13888 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_116
timestamp 1698431365
transform 1 0 14336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_118
timestamp 1698431365
transform 1 0 14560 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_131
timestamp 1698431365
transform 1 0 16016 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_158
timestamp 1698431365
transform 1 0 19040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_172
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_204
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_288
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_320
timestamp 1698431365
transform 1 0 37184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_328
timestamp 1698431365
transform 1 0 38080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_332
timestamp 1698431365
transform 1 0 38528 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_345
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_380
timestamp 1698431365
transform 1 0 43904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_115
timestamp 1698431365
transform 1 0 14224 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_118
timestamp 1698431365
transform 1 0 14560 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_134
timestamp 1698431365
transform 1 0 16352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_136
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_143
timestamp 1698431365
transform 1 0 17360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_151
timestamp 1698431365
transform 1 0 18256 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_165
timestamp 1698431365
transform 1 0 19824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_187
timestamp 1698431365
transform 1 0 22288 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_195
timestamp 1698431365
transform 1 0 23184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_205
timestamp 1698431365
transform 1 0 24304 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_215
timestamp 1698431365
transform 1 0 25424 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_223
timestamp 1698431365
transform 1 0 26320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_227
timestamp 1698431365
transform 1 0 26768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_239
timestamp 1698431365
transform 1 0 28112 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_243
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_263
timestamp 1698431365
transform 1 0 30800 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_275
timestamp 1698431365
transform 1 0 32144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_279
timestamp 1698431365
transform 1 0 32592 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_321
timestamp 1698431365
transform 1 0 37296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_331
timestamp 1698431365
transform 1 0 38416 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_353
timestamp 1698431365
transform 1 0 40880 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_357
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_359
timestamp 1698431365
transform 1 0 41552 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_70
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_108
timestamp 1698431365
transform 1 0 13440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_122
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_148
timestamp 1698431365
transform 1 0 17920 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_156
timestamp 1698431365
transform 1 0 18816 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_183
timestamp 1698431365
transform 1 0 21840 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_197
timestamp 1698431365
transform 1 0 23408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_201
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_220
timestamp 1698431365
transform 1 0 25984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_222
timestamp 1698431365
transform 1 0 26208 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_233
timestamp 1698431365
transform 1 0 27440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_235
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_246
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_262
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_264
timestamp 1698431365
transform 1 0 30912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_271
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_293
timestamp 1698431365
transform 1 0 34160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_301
timestamp 1698431365
transform 1 0 35056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_303
timestamp 1698431365
transform 1 0 35280 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_318
timestamp 1698431365
transform 1 0 36960 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_325
timestamp 1698431365
transform 1 0 37744 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_329
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_370
timestamp 1698431365
transform 1 0 42784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_376
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 23968 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform 1 0 18144 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform 1 0 3584 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 13440 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 24752 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 13104 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 35728 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 24528 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 35504 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 43568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform 1 0 10416 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 39872 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform -1 0 44352 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform 1 0 14336 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 43456 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 43456 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 36400 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform 1 0 34384 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 15904 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform 1 0 17584 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform -1 0 38864 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 8624 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 43568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 16912 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform 1 0 14000 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 28336 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 27552 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 35728 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform -1 0 43456 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform -1 0 27328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform -1 0 40432 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform -1 0 32592 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 43456 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform 1 0 5824 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold50
timestamp 1698431365
transform -1 0 43568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform -1 0 43568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform -1 0 32144 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform -1 0 44128 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform -1 0 29792 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 23968 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform -1 0 39648 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 34608 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform -1 0 14224 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform -1 0 35952 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform -1 0 42448 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform -1 0 35952 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 43456 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform -1 0 27888 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform 1 0 6384 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 38528 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform -1 0 23968 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold69
timestamp 1698431365
transform -1 0 29344 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold70
timestamp 1698431365
transform -1 0 35168 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold71
timestamp 1698431365
transform 1 0 17136 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold72
timestamp 1698431365
transform 1 0 13888 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold73
timestamp 1698431365
transform 1 0 9632 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold74
timestamp 1698431365
transform 1 0 2128 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold75
timestamp 1698431365
transform 1 0 6384 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold76
timestamp 1698431365
transform -1 0 8848 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold77
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold78
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold79
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold80
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold81
timestamp 1698431365
transform -1 0 36064 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold82
timestamp 1698431365
transform -1 0 13104 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold83
timestamp 1698431365
transform -1 0 43568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold84
timestamp 1698431365
transform -1 0 32480 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold85
timestamp 1698431365
transform -1 0 43568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold86
timestamp 1698431365
transform -1 0 31808 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold87
timestamp 1698431365
transform -1 0 32704 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold88
timestamp 1698431365
transform -1 0 31808 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold89
timestamp 1698431365
transform 1 0 6384 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold90
timestamp 1698431365
transform -1 0 21056 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold91
timestamp 1698431365
transform -1 0 43568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold92
timestamp 1698431365
transform 1 0 21728 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold93
timestamp 1698431365
transform -1 0 30688 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold94
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold95
timestamp 1698431365
transform 1 0 6384 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold96
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold97
timestamp 1698431365
transform -1 0 32368 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold98
timestamp 1698431365
transform -1 0 39648 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold99
timestamp 1698431365
transform -1 0 43456 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold100
timestamp 1698431365
transform -1 0 20832 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold101
timestamp 1698431365
transform -1 0 34608 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold102
timestamp 1698431365
transform -1 0 8288 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold103
timestamp 1698431365
transform -1 0 43568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold104
timestamp 1698431365
transform -1 0 43568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold105
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold106
timestamp 1698431365
transform -1 0 21392 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold107
timestamp 1698431365
transform -1 0 14448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold108
timestamp 1698431365
transform -1 0 24864 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold109
timestamp 1698431365
transform -1 0 31808 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 44352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 13664 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 43680 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 25760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 38416 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 20272 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 33040 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 20272 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 27664 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 44352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 22288 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 28896 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 35952 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 35840 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 17584 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 14336 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 23632 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 41440 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 20608 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 44352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 44352 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 37072 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 26320 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 44352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 19600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 42112 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 43680 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 44352 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 44352 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output39
timestamp 1698431365
transform -1 0 34160 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output40
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41
timestamp 1698431365
transform -1 0 20384 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42
timestamp 1698431365
transform -1 0 25536 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 39760 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform -1 0 39424 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform 1 0 26320 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform -1 0 42784 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output49
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output50
timestamp 1698431365
transform 1 0 42784 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output51
timestamp 1698431365
transform -1 0 37408 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output52
timestamp 1698431365
transform 1 0 42784 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform 1 0 41664 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform 1 0 18704 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output55
timestamp 1698431365
transform -1 0 16576 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output56
timestamp 1698431365
transform 1 0 42784 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output57
timestamp 1698431365
transform 1 0 25984 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform 1 0 20720 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output60
timestamp 1698431365
transform 1 0 33712 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output62
timestamp 1698431365
transform 1 0 42784 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output63
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output64
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform 1 0 22288 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform 1 0 26992 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform -1 0 35952 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output69
timestamp 1698431365
transform 1 0 43232 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output70
timestamp 1698431365
transform 1 0 41664 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output71
timestamp 1698431365
transform 1 0 42784 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output72
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output73
timestamp 1698431365
transform 1 0 42784 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_50 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__74 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25424 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__75
timestamp 1698431365
transform -1 0 22960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__76
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__77
timestamp 1698431365
transform 1 0 43456 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__78
timestamp 1698431365
transform -1 0 26768 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__79
timestamp 1698431365
transform -1 0 17360 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__80
timestamp 1698431365
transform -1 0 32144 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__81
timestamp 1698431365
transform 1 0 42560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__82
timestamp 1698431365
transform 1 0 42560 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__83
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__84
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__85
timestamp 1698431365
transform 1 0 39312 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__86
timestamp 1698431365
transform -1 0 40208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__87
timestamp 1698431365
transform 1 0 43904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__88
timestamp 1698431365
transform -1 0 36960 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__89
timestamp 1698431365
transform -1 0 41664 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__90
timestamp 1698431365
transform -1 0 31472 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__91
timestamp 1698431365
transform -1 0 37856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__92
timestamp 1698431365
transform 1 0 42112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__93
timestamp 1698431365
transform 1 0 43904 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__94
timestamp 1698431365
transform 1 0 41216 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__95
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__96
timestamp 1698431365
transform 1 0 42336 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__97
timestamp 1698431365
transform -1 0 35056 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__2__98
timestamp 1698431365
transform 1 0 43904 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_115
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_123
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_124
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_128
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_129
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_130
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_135
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_141
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_143
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_146
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_147
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_148
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_151
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_152
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_153
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_154
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_156
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_157
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_158
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_159
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_161
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_162
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_163
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_164
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_165
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_166
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_167
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_168
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_169
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_170
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_171
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_172
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_173
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_174
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_175
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_176
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_178
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_179
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_180
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_181
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_183
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_184
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_185
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_188
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_189
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_190
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_193
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_194
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_195
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_209
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_210
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_213
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_214
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_215
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_218
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_219
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_220
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_222
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_223
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_224
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_225
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_227
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_228
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_229
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_230
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_231
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_232
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_233
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_234
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_235
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_236
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_237
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_238
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_239
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_240
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_241
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_242
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_243
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_244
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_245
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_246
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_247
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_248
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_249
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_250
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_251
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_252
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_253
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_254
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_255
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_256
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_257
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_258
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_259
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_260
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_261
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_262
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_263
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_264
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_265
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_266
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_267
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_268
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_269
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_270
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_271
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_272
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_273
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_274
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_275
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_276
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_277
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_278
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_279
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_280
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_281
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_282
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_283
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_284
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_285
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_287
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_288
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_289
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_290
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_292
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_293
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_294
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_295
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_298
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_299
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_300
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_301
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_302
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_303
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_304
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_305
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_306
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_307
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_308
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_309
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_310
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_311
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_312
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_313
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_314
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_315
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_316
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_317
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_318
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_319
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_320
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_321
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_322
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_323
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_324
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_325
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_326
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_327
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_328
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_329
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_330
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_331
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_332
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_333
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_334
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_335
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_336
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_337
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_338
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_339
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_340
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_343
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_344
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_345
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_346
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_347
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_348
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_349
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_350
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_351
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_352
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_353
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_354
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_355
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_356
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_357
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_358
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_359
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_360
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_361
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 2 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 3 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 45200 22176 46000 22288 0 FreeSans 448 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal3 s 45200 2016 46000 2128 0 FreeSans 448 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 14112 45200 14224 46000 0 FreeSans 448 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 45200 2688 46000 2800 0 FreeSans 448 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 20160 45200 20272 46000 0 FreeSans 448 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 chanx_left_in[2]
port 18 nsew signal input
flabel metal3 s 45200 8736 46000 8848 0 FreeSans 448 0 0 0 chanx_left_in[3]
port 19 nsew signal input
flabel metal2 s 21504 45200 21616 46000 0 FreeSans 448 90 0 0 chanx_left_in[4]
port 20 nsew signal input
flabel metal2 s 27552 45200 27664 46000 0 FreeSans 448 90 0 0 chanx_left_in[5]
port 21 nsew signal input
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 chanx_left_in[6]
port 22 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 chanx_left_in[7]
port 23 nsew signal input
flabel metal2 s 35616 45200 35728 46000 0 FreeSans 448 90 0 0 chanx_left_in[8]
port 24 nsew signal input
flabel metal2 s 17472 45200 17584 46000 0 FreeSans 448 90 0 0 chanx_left_in[9]
port 25 nsew signal input
flabel metal3 s 45200 34944 46000 35056 0 FreeSans 448 0 0 0 chanx_left_out[0]
port 26 nsew signal tristate
flabel metal2 s 32928 45200 33040 46000 0 FreeSans 448 90 0 0 chanx_left_out[10]
port 27 nsew signal tristate
flabel metal2 s 24192 45200 24304 46000 0 FreeSans 448 90 0 0 chanx_left_out[11]
port 28 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 chanx_left_out[12]
port 29 nsew signal tristate
flabel metal2 s 19488 45200 19600 46000 0 FreeSans 448 90 0 0 chanx_left_out[13]
port 30 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 chanx_left_out[14]
port 31 nsew signal tristate
flabel metal3 s 45200 8064 46000 8176 0 FreeSans 448 0 0 0 chanx_left_out[15]
port 32 nsew signal tristate
flabel metal2 s 41664 45200 41776 46000 0 FreeSans 448 90 0 0 chanx_left_out[16]
port 33 nsew signal tristate
flabel metal2 s 39648 45200 39760 46000 0 FreeSans 448 90 0 0 chanx_left_out[17]
port 34 nsew signal tristate
flabel metal2 s 38304 45200 38416 46000 0 FreeSans 448 90 0 0 chanx_left_out[18]
port 35 nsew signal tristate
flabel metal2 s 26208 45200 26320 46000 0 FreeSans 448 90 0 0 chanx_left_out[19]
port 36 nsew signal tristate
flabel metal2 s 16128 45200 16240 46000 0 FreeSans 448 90 0 0 chanx_left_out[1]
port 37 nsew signal tristate
flabel metal3 s 45200 45696 46000 45808 0 FreeSans 448 0 0 0 chanx_left_out[2]
port 38 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chanx_left_out[3]
port 39 nsew signal tristate
flabel metal2 s 34272 45200 34384 46000 0 FreeSans 448 90 0 0 chanx_left_out[4]
port 40 nsew signal tristate
flabel metal3 s 45200 41664 46000 41776 0 FreeSans 448 0 0 0 chanx_left_out[5]
port 41 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 chanx_left_out[6]
port 42 nsew signal tristate
flabel metal3 s 45200 31584 46000 31696 0 FreeSans 448 0 0 0 chanx_left_out[7]
port 43 nsew signal tristate
flabel metal3 s 45200 6720 46000 6832 0 FreeSans 448 0 0 0 chanx_left_out[8]
port 44 nsew signal tristate
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 chanx_left_out[9]
port 45 nsew signal tristate
flabel metal2 s 14784 45200 14896 46000 0 FreeSans 448 90 0 0 chanx_right_in[0]
port 46 nsew signal input
flabel metal2 s 23520 45200 23632 46000 0 FreeSans 448 90 0 0 chanx_right_in[10]
port 47 nsew signal input
flabel metal2 s 40320 45200 40432 46000 0 FreeSans 448 90 0 0 chanx_right_in[11]
port 48 nsew signal input
flabel metal2 s 18816 45200 18928 46000 0 FreeSans 448 90 0 0 chanx_right_in[12]
port 49 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 chanx_right_in[13]
port 50 nsew signal input
flabel metal3 s 45200 3360 46000 3472 0 FreeSans 448 0 0 0 chanx_right_in[14]
port 51 nsew signal input
flabel metal3 s 45200 40992 46000 41104 0 FreeSans 448 0 0 0 chanx_right_in[15]
port 52 nsew signal input
flabel metal2 s 36960 45200 37072 46000 0 FreeSans 448 90 0 0 chanx_right_in[16]
port 53 nsew signal input
flabel metal2 s 37632 45200 37744 46000 0 FreeSans 448 90 0 0 chanx_right_in[17]
port 54 nsew signal input
flabel metal2 s 25536 45200 25648 46000 0 FreeSans 448 90 0 0 chanx_right_in[18]
port 55 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 chanx_right_in[19]
port 56 nsew signal input
flabel metal3 s 45200 44352 46000 44464 0 FreeSans 448 0 0 0 chanx_right_in[1]
port 57 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 chanx_right_in[2]
port 58 nsew signal input
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 chanx_right_in[3]
port 59 nsew signal input
flabel metal3 s 45200 42336 46000 42448 0 FreeSans 448 0 0 0 chanx_right_in[4]
port 60 nsew signal input
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 chanx_right_in[5]
port 61 nsew signal input
flabel metal3 s 45200 30912 46000 31024 0 FreeSans 448 0 0 0 chanx_right_in[6]
port 62 nsew signal input
flabel metal3 s 45200 43008 46000 43120 0 FreeSans 448 0 0 0 chanx_right_in[7]
port 63 nsew signal input
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 chanx_right_in[8]
port 64 nsew signal input
flabel metal2 s 32256 45200 32368 46000 0 FreeSans 448 90 0 0 chanx_right_in[9]
port 65 nsew signal input
flabel metal3 s 45200 36960 46000 37072 0 FreeSans 448 0 0 0 chanx_right_out[0]
port 66 nsew signal tristate
flabel metal2 s 18144 45200 18256 46000 0 FreeSans 448 90 0 0 chanx_right_out[10]
port 67 nsew signal tristate
flabel metal2 s 15456 45200 15568 46000 0 FreeSans 448 90 0 0 chanx_right_out[11]
port 68 nsew signal tristate
flabel metal2 s 30912 45200 31024 46000 0 FreeSans 448 90 0 0 chanx_right_out[12]
port 69 nsew signal tristate
flabel metal3 s 45200 5376 46000 5488 0 FreeSans 448 0 0 0 chanx_right_out[13]
port 70 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 chanx_right_out[14]
port 71 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 chanx_right_out[15]
port 72 nsew signal tristate
flabel metal2 s 40992 45200 41104 46000 0 FreeSans 448 90 0 0 chanx_right_out[16]
port 73 nsew signal tristate
flabel metal2 s 20832 45200 20944 46000 0 FreeSans 448 90 0 0 chanx_right_out[17]
port 74 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 chanx_right_out[18]
port 75 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 chanx_right_out[19]
port 76 nsew signal tristate
flabel metal3 s 45200 7392 46000 7504 0 FreeSans 448 0 0 0 chanx_right_out[1]
port 77 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 chanx_right_out[2]
port 78 nsew signal tristate
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 chanx_right_out[3]
port 79 nsew signal tristate
flabel metal3 s 45200 4032 46000 4144 0 FreeSans 448 0 0 0 chanx_right_out[4]
port 80 nsew signal tristate
flabel metal2 s 22176 45200 22288 46000 0 FreeSans 448 90 0 0 chanx_right_out[5]
port 81 nsew signal tristate
flabel metal2 s 26880 45200 26992 46000 0 FreeSans 448 90 0 0 chanx_right_out[6]
port 82 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 chanx_right_out[7]
port 83 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 chanx_right_out[8]
port 84 nsew signal tristate
flabel metal2 s 38976 45200 39088 46000 0 FreeSans 448 90 0 0 chanx_right_out[9]
port 85 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 chany_bottom_in[0]
port 86 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 chany_bottom_in[10]
port 87 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 chany_bottom_in[11]
port 88 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chany_bottom_in[12]
port 89 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chany_bottom_in[13]
port 90 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chany_bottom_in[14]
port 91 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chany_bottom_in[15]
port 92 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chany_bottom_in[16]
port 93 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chany_bottom_in[17]
port 94 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chany_bottom_in[18]
port 95 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 chany_bottom_in[19]
port 96 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chany_bottom_in[1]
port 97 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chany_bottom_in[2]
port 98 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chany_bottom_in[3]
port 99 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 chany_bottom_in[4]
port 100 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chany_bottom_in[5]
port 101 nsew signal input
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 chany_bottom_in[6]
port 102 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 chany_bottom_in[7]
port 103 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chany_bottom_in[8]
port 104 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 chany_bottom_in[9]
port 105 nsew signal input
flabel metal2 s 36288 45200 36400 46000 0 FreeSans 448 90 0 0 chany_bottom_out[0]
port 106 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 chany_bottom_out[10]
port 107 nsew signal tristate
flabel metal3 s 45200 36288 46000 36400 0 FreeSans 448 0 0 0 chany_bottom_out[11]
port 108 nsew signal tristate
flabel metal3 s 45200 37632 46000 37744 0 FreeSans 448 0 0 0 chany_bottom_out[12]
port 109 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 chany_bottom_out[13]
port 110 nsew signal tristate
flabel metal2 s 24864 45200 24976 46000 0 FreeSans 448 90 0 0 chany_bottom_out[14]
port 111 nsew signal tristate
flabel metal3 s 45200 45024 46000 45136 0 FreeSans 448 0 0 0 chany_bottom_out[15]
port 112 nsew signal tristate
flabel metal2 s 42336 45200 42448 46000 0 FreeSans 448 90 0 0 chany_bottom_out[16]
port 113 nsew signal tristate
flabel metal3 s 45200 43680 46000 43792 0 FreeSans 448 0 0 0 chany_bottom_out[17]
port 114 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 chany_bottom_out[18]
port 115 nsew signal tristate
flabel metal3 s 45200 6048 46000 6160 0 FreeSans 448 0 0 0 chany_bottom_out[19]
port 116 nsew signal tristate
flabel metal3 s 45200 35616 46000 35728 0 FreeSans 448 0 0 0 chany_bottom_out[1]
port 117 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal3 s 45200 40320 46000 40432 0 FreeSans 448 0 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal3 s 45200 39648 46000 39760 0 FreeSans 448 0 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal3 s 45200 38976 46000 39088 0 FreeSans 448 0 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal3 s 45200 38304 46000 38416 0 FreeSans 448 0 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal3 s 45200 4704 46000 4816 0 FreeSans 448 0 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 31584 45200 31696 46000 0 FreeSans 448 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 16800 45200 16912 46000 0 FreeSans 448 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 126 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 127 nsew signal input
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 128 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 129 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 131 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 pReset
port 132 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 prog_clk
port 133 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 134 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 135 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 138 nsew signal input
flabel metal3 s 45200 0 46000 112 0 FreeSans 448 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 139 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal2 14056 25312 14056 25312 0 _000_
rlabel metal2 12600 25536 12600 25536 0 _001_
rlabel metal2 13496 24472 13496 24472 0 _002_
rlabel metal2 8680 26600 8680 26600 0 _003_
rlabel metal2 7000 27496 7000 27496 0 _004_
rlabel metal2 3080 28392 3080 28392 0 _005_
rlabel metal2 2856 25200 2856 25200 0 _006_
rlabel metal2 3080 27048 3080 27048 0 _007_
rlabel metal2 16184 24752 16184 24752 0 _008_
rlabel metal2 13944 21280 13944 21280 0 _009_
rlabel metal2 12488 20888 12488 20888 0 _010_
rlabel metal2 11928 21336 11928 21336 0 _011_
rlabel metal2 10920 21056 10920 21056 0 _012_
rlabel metal2 7672 22288 7672 22288 0 _013_
rlabel metal2 8680 21112 8680 21112 0 _014_
rlabel metal2 6216 22792 6216 22792 0 _015_
rlabel metal2 14168 27552 14168 27552 0 _016_
rlabel metal3 13552 26936 13552 26936 0 _017_
rlabel metal2 10808 28224 10808 28224 0 _018_
rlabel metal2 6328 26208 6328 26208 0 _019_
rlabel metal3 19208 25256 19208 25256 0 _020_
rlabel metal2 19096 26152 19096 26152 0 _021_
rlabel metal3 24808 29624 24808 29624 0 _022_
rlabel metal2 20664 29064 20664 29064 0 _023_
rlabel metal2 20440 29848 20440 29848 0 _024_
rlabel metal3 18704 25592 18704 25592 0 _025_
rlabel metal2 18648 27328 18648 27328 0 _026_
rlabel metal2 16744 29008 16744 29008 0 _027_
rlabel metal2 23464 27552 23464 27552 0 _028_
rlabel metal2 22792 25536 22792 25536 0 _029_
rlabel metal3 35504 25256 35504 25256 0 _030_
rlabel metal2 31864 28896 31864 28896 0 _031_
rlabel metal2 29400 29792 29400 29792 0 _032_
rlabel metal2 27160 29232 27160 29232 0 _033_
rlabel metal2 35784 29232 35784 29232 0 _034_
rlabel metal2 33432 26656 33432 26656 0 _035_
rlabel metal2 31808 24808 31808 24808 0 _036_
rlabel metal2 29400 25872 29400 25872 0 _037_
rlabel metal2 28056 28224 28056 28224 0 _038_
rlabel metal3 27104 26936 27104 26936 0 _039_
rlabel metal2 26600 19656 26600 19656 0 _040_
rlabel metal2 25256 18704 25256 18704 0 _041_
rlabel metal2 21896 20552 21896 20552 0 _042_
rlabel metal2 22120 19712 22120 19712 0 _043_
rlabel metal2 21448 18872 21448 18872 0 _044_
rlabel metal2 16408 22624 16408 22624 0 _045_
rlabel metal2 23128 21840 23128 21840 0 _046_
rlabel metal2 23464 23968 23464 23968 0 _047_
rlabel metal2 21336 20552 21336 20552 0 _048_
rlabel metal2 19992 19768 19992 19768 0 _049_
rlabel metal2 29624 21196 29624 21196 0 _050_
rlabel metal2 28392 20356 28392 20356 0 _051_
rlabel metal3 33040 23352 33040 23352 0 _052_
rlabel metal2 33096 21896 33096 21896 0 _053_
rlabel metal2 32200 23464 32200 23464 0 _054_
rlabel metal2 29960 23296 29960 23296 0 _055_
rlabel metal2 28952 22400 28952 22400 0 _056_
rlabel metal2 28168 23072 28168 23072 0 _057_
rlabel metal3 43120 21448 43120 21448 0 _058_
rlabel metal2 40936 21336 40936 21336 0 _059_
rlabel metal2 43960 22624 43960 22624 0 _060_
rlabel metal2 39704 22344 39704 22344 0 _061_
rlabel metal2 37408 21784 37408 21784 0 _062_
rlabel metal2 37016 21504 37016 21504 0 _063_
rlabel metal2 41272 23744 41272 23744 0 _064_
rlabel metal2 40712 26096 40712 26096 0 _065_
rlabel metal2 40152 27440 40152 27440 0 _066_
rlabel metal2 40040 25816 40040 25816 0 _067_
rlabel metal2 39368 26376 39368 26376 0 _068_
rlabel metal2 36960 24024 36960 24024 0 _069_
rlabel metal2 43960 17080 43960 17080 0 _070_
rlabel metal2 39984 17080 39984 17080 0 _071_
rlabel metal2 39816 17696 39816 17696 0 _072_
rlabel metal2 36232 19264 36232 19264 0 _073_
rlabel metal2 36120 18032 36120 18032 0 _074_
rlabel metal3 36232 20776 36232 20776 0 _075_
rlabel metal2 44072 15568 44072 15568 0 _076_
rlabel metal2 38136 15456 38136 15456 0 _077_
rlabel metal2 36064 14616 36064 14616 0 _078_
rlabel metal2 34440 16408 34440 16408 0 _079_
rlabel metal2 31864 16240 31864 16240 0 _080_
rlabel metal2 29624 17472 29624 17472 0 _081_
rlabel metal3 24976 13384 24976 13384 0 _082_
rlabel metal2 26376 15400 26376 15400 0 _083_
rlabel metal2 24248 15456 24248 15456 0 _084_
rlabel metal2 30184 14784 30184 14784 0 _085_
rlabel metal2 32088 15624 32088 15624 0 _086_
rlabel metal2 30296 15456 30296 15456 0 _087_
rlabel metal2 25928 16576 25928 16576 0 _088_
rlabel metal2 27384 15512 27384 15512 0 _089_
rlabel metal2 17528 16352 17528 16352 0 _090_
rlabel metal2 17752 15456 17752 15456 0 _091_
rlabel metal3 21000 17752 21000 17752 0 _092_
rlabel metal3 19600 16296 19600 16296 0 _093_
rlabel metal2 12600 18088 12600 18088 0 _094_
rlabel metal2 22120 16128 22120 16128 0 _095_
rlabel metal2 14728 15176 14728 15176 0 _096_
rlabel metal3 13272 14616 13272 14616 0 _097_
rlabel metal2 14168 17920 14168 17920 0 _098_
rlabel metal2 15624 17024 15624 17024 0 _099_
rlabel metal2 11144 16408 11144 16408 0 _100_
rlabel metal2 6216 18088 6216 18088 0 _101_
rlabel metal2 9912 15624 9912 15624 0 _102_
rlabel metal2 10136 19488 10136 19488 0 _103_
rlabel metal2 5432 14952 5432 14952 0 _104_
rlabel metal2 2072 16912 2072 16912 0 _105_
rlabel metal2 2184 17416 2184 17416 0 _106_
rlabel metal2 4984 16072 4984 16072 0 _107_
rlabel metal2 6328 19712 6328 19712 0 _108_
rlabel metal2 5656 20412 5656 20412 0 _109_
rlabel metal2 21000 27328 21000 27328 0 _110_
rlabel metal2 8344 26096 8344 26096 0 _111_
rlabel metal2 6776 24080 6776 24080 0 _112_
rlabel metal2 21672 29792 21672 29792 0 _113_
rlabel metal2 31416 25424 31416 25424 0 _114_
rlabel metal3 21672 24584 21672 24584 0 _115_
rlabel metal2 31640 23856 31640 23856 0 _116_
rlabel metal2 43736 23380 43736 23380 0 _117_
rlabel metal2 43736 17360 43736 17360 0 _118_
rlabel metal2 31584 15400 31584 15400 0 _119_
rlabel metal2 21672 14448 21672 14448 0 _120_
rlabel metal2 5992 20412 5992 20412 0 _121_
rlabel metal2 1736 27720 1736 27720 0 ccff_head
rlabel metal3 44520 22288 44520 22288 0 ccff_tail
rlabel metal2 44408 3192 44408 3192 0 chanx_left_in[0]
rlabel metal2 14168 44478 14168 44478 0 chanx_left_in[10]
rlabel metal2 43176 3080 43176 3080 0 chanx_left_in[12]
rlabel metal2 24864 4200 24864 4200 0 chanx_left_in[13]
rlabel metal2 38584 4256 38584 4256 0 chanx_left_in[14]
rlabel metal2 20440 41216 20440 41216 0 chanx_left_in[16]
rlabel metal2 33208 4088 33208 4088 0 chanx_left_in[17]
rlabel metal2 31080 3416 31080 3416 0 chanx_left_in[18]
rlabel metal2 20216 2422 20216 2422 0 chanx_left_in[1]
rlabel metal3 26824 4200 26824 4200 0 chanx_left_in[2]
rlabel metal2 44184 8904 44184 8904 0 chanx_left_in[3]
rlabel metal2 22008 41216 22008 41216 0 chanx_left_in[4]
rlabel metal2 27608 44478 27608 44478 0 chanx_left_in[5]
rlabel metal2 36120 3920 36120 3920 0 chanx_left_in[6]
rlabel metal2 35616 41944 35616 41944 0 chanx_left_in[8]
rlabel metal2 17528 44478 17528 44478 0 chanx_left_in[9]
rlabel metal2 32984 44478 32984 44478 0 chanx_left_out[10]
rlabel metal2 24248 44478 24248 44478 0 chanx_left_out[11]
rlabel metal2 19544 44478 19544 44478 0 chanx_left_out[13]
rlabel metal2 23576 2030 23576 2030 0 chanx_left_out[14]
rlabel metal3 44674 8120 44674 8120 0 chanx_left_out[15]
rlabel metal2 39704 44478 39704 44478 0 chanx_left_out[17]
rlabel metal2 38360 44478 38360 44478 0 chanx_left_out[18]
rlabel metal2 26936 41888 26936 41888 0 chanx_left_out[19]
rlabel metal2 16184 44478 16184 44478 0 chanx_left_out[1]
rlabel metal3 43610 45752 43610 45752 0 chanx_left_out[2]
rlabel metal2 18872 2030 18872 2030 0 chanx_left_out[3]
rlabel metal2 44072 41496 44072 41496 0 chanx_left_out[5]
rlabel metal2 36456 2464 36456 2464 0 chanx_left_out[6]
rlabel metal3 44674 31640 44674 31640 0 chanx_left_out[7]
rlabel metal2 41720 2198 41720 2198 0 chanx_left_out[9]
rlabel metal2 14840 44478 14840 44478 0 chanx_right_in[0]
rlabel metal2 23800 41216 23800 41216 0 chanx_right_in[10]
rlabel metal2 40376 44478 40376 44478 0 chanx_right_in[11]
rlabel metal2 20216 40656 20216 40656 0 chanx_right_in[12]
rlabel metal2 23800 3024 23800 3024 0 chanx_right_in[13]
rlabel metal3 44730 3416 44730 3416 0 chanx_right_in[14]
rlabel metal2 44520 41440 44520 41440 0 chanx_right_in[15]
rlabel metal2 37016 44478 37016 44478 0 chanx_right_in[16]
rlabel metal2 37912 41216 37912 41216 0 chanx_right_in[17]
rlabel metal2 25592 44478 25592 44478 0 chanx_right_in[18]
rlabel metal3 44618 44408 44618 44408 0 chanx_right_in[1]
rlabel metal2 19768 3808 19768 3808 0 chanx_right_in[2]
rlabel metal2 41272 3360 41272 3360 0 chanx_right_in[3]
rlabel metal2 43792 37464 43792 37464 0 chanx_right_in[4]
rlabel metal2 36568 4592 36568 4592 0 chanx_right_in[5]
rlabel metal3 44450 30968 44450 30968 0 chanx_right_in[6]
rlabel metal2 44408 40600 44408 40600 0 chanx_right_in[7]
rlabel metal2 41160 3864 41160 3864 0 chanx_right_in[8]
rlabel metal2 32312 44478 32312 44478 0 chanx_right_in[9]
rlabel metal2 19320 41328 19320 41328 0 chanx_right_out[10]
rlabel metal2 15512 44478 15512 44478 0 chanx_right_out[11]
rlabel metal2 44072 5600 44072 5600 0 chanx_right_out[13]
rlabel metal2 25592 2198 25592 2198 0 chanx_right_out[14]
rlabel metal2 38416 3304 38416 3304 0 chanx_right_out[15]
rlabel metal2 20888 44478 20888 44478 0 chanx_right_out[17]
rlabel metal2 34216 3640 34216 3640 0 chanx_right_out[18]
rlabel metal3 32144 3640 32144 3640 0 chanx_right_out[19]
rlabel metal3 44674 7448 44674 7448 0 chanx_right_out[1]
rlabel metal2 20888 1246 20888 1246 0 chanx_right_out[2]
rlabel metal3 28224 3640 28224 3640 0 chanx_right_out[3]
rlabel metal2 22736 45304 22736 45304 0 chanx_right_out[5]
rlabel metal2 26936 44478 26936 44478 0 chanx_right_out[6]
rlabel metal2 34888 4088 34888 4088 0 chanx_right_out[7]
rlabel metal2 40376 41888 40376 41888 0 chanx_right_out[9]
rlabel metal3 44786 45080 44786 45080 0 chany_bottom_out[15]
rlabel metal2 42392 43554 42392 43554 0 chany_bottom_out[16]
rlabel metal3 44506 43736 44506 43736 0 chany_bottom_out[17]
rlabel metal2 39032 2198 39032 2198 0 chany_bottom_out[18]
rlabel metal2 44072 6328 44072 6328 0 chany_bottom_out[19]
rlabel metal2 15680 27720 15680 27720 0 clknet_0_prog_clk
rlabel metal2 5320 21952 5320 21952 0 clknet_3_0__leaf_prog_clk
rlabel metal3 12320 16856 12320 16856 0 clknet_3_1__leaf_prog_clk
rlabel metal2 3976 27384 3976 27384 0 clknet_3_2__leaf_prog_clk
rlabel metal2 19712 28616 19712 28616 0 clknet_3_3__leaf_prog_clk
rlabel metal2 30296 19880 30296 19880 0 clknet_3_4__leaf_prog_clk
rlabel metal2 40376 15288 40376 15288 0 clknet_3_5__leaf_prog_clk
rlabel metal2 21336 28616 21336 28616 0 clknet_3_6__leaf_prog_clk
rlabel metal2 30072 23128 30072 23128 0 clknet_3_7__leaf_prog_clk
rlabel metal2 36568 29456 36568 29456 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal3 40264 26376 40264 26376 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal3 41720 27944 41720 27944 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 40656 27272 40656 27272 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 42840 27272 42840 27272 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal3 42504 25368 42504 25368 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal2 41720 23688 41720 23688 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal3 23072 16632 23072 16632 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal2 17248 12264 17248 12264 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal3 17640 14392 17640 14392 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal2 17528 12824 17528 12824 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal3 22344 18200 22344 18200 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal2 16632 13776 16632 13776 0 mem_bottom_track_15.DFFR_0_.Q
rlabel metal2 14224 12264 14224 12264 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal2 12488 13216 12488 13216 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal2 13048 16632 13048 16632 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 16016 14392 16016 14392 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal2 12824 14728 12824 14728 0 mem_bottom_track_19.DFFR_1_.Q
rlabel metal2 6104 15512 6104 15512 0 mem_bottom_track_21.DFFR_0_.Q
rlabel metal2 5544 18144 5544 18144 0 mem_bottom_track_21.DFFR_1_.Q
rlabel metal2 12432 14392 12432 14392 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal2 8008 15624 8008 15624 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal2 1680 16856 1680 16856 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 4984 13160 4984 13160 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal2 8456 14448 8456 14448 0 mem_bottom_track_27.DFFR_0_.Q
rlabel metal2 2408 15512 2408 15512 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal2 3080 17864 3080 17864 0 mem_bottom_track_29.DFFR_0_.Q
rlabel metal2 7280 18536 7280 18536 0 mem_bottom_track_29.DFFR_1_.Q
rlabel metal2 35784 16408 35784 16408 0 mem_bottom_track_3.DFFR_0_.Q
rlabel metal2 36680 17248 36680 17248 0 mem_bottom_track_3.DFFR_1_.Q
rlabel metal2 37072 19768 37072 19768 0 mem_bottom_track_3.DFFR_2_.Q
rlabel metal3 41720 15960 41720 15960 0 mem_bottom_track_3.DFFR_3_.Q
rlabel metal2 42952 14784 42952 14784 0 mem_bottom_track_3.DFFR_4_.Q
rlabel metal2 38248 14336 38248 14336 0 mem_bottom_track_3.DFFR_5_.Q
rlabel metal2 29176 16520 29176 16520 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal2 32648 17304 32648 17304 0 mem_bottom_track_5.DFFR_1_.Q
rlabel metal2 35672 13384 35672 13384 0 mem_bottom_track_5.DFFR_2_.Q
rlabel metal2 39032 13552 39032 13552 0 mem_bottom_track_5.DFFR_3_.Q
rlabel metal2 42056 13384 42056 13384 0 mem_bottom_track_5.DFFR_4_.Q
rlabel metal2 34888 11984 34888 11984 0 mem_bottom_track_5.DFFR_5_.Q
rlabel metal2 30856 14784 30856 14784 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal2 35504 12264 35504 12264 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal2 28056 11984 28056 11984 0 mem_bottom_track_7.DFFR_2_.Q
rlabel metal2 27272 12936 27272 12936 0 mem_bottom_track_7.DFFR_3_.Q
rlabel metal2 30408 14056 30408 14056 0 mem_bottom_track_7.DFFR_4_.Q
rlabel metal2 23016 11984 23016 11984 0 mem_bottom_track_7.DFFR_5_.Q
rlabel metal3 29064 12824 29064 12824 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal2 3080 21000 3080 21000 0 mem_left_track_1.DFFR_0_.Q
rlabel metal2 9240 23184 9240 23184 0 mem_left_track_1.DFFR_1_.Q
rlabel metal3 4984 22232 4984 22232 0 mem_left_track_1.DFFR_2_.Q
rlabel metal3 10864 20552 10864 20552 0 mem_left_track_1.DFFR_3_.Q
rlabel metal3 6776 23240 6776 23240 0 mem_left_track_1.DFFR_4_.Q
rlabel metal3 13720 21896 13720 21896 0 mem_left_track_1.DFFR_5_.Q
rlabel metal3 12208 21000 12208 21000 0 mem_left_track_1.DFFR_6_.Q
rlabel metal2 7000 23296 7000 23296 0 mem_left_track_1.DFFR_7_.Q
rlabel metal2 29288 15904 29288 15904 0 mem_left_track_17.DFFR_0_.D
rlabel metal2 39256 19936 39256 19936 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 29064 18872 29064 18872 0 mem_left_track_17.DFFR_1_.Q
rlabel metal3 15512 22232 15512 22232 0 mem_left_track_17.DFFR_2_.Q
rlabel metal3 20048 21784 20048 21784 0 mem_left_track_17.DFFR_3_.Q
rlabel metal2 22680 22288 22680 22288 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 22344 22400 22344 22400 0 mem_left_track_17.DFFR_5_.Q
rlabel metal2 31976 22680 31976 22680 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 31192 21000 31192 21000 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 30632 21784 30632 21784 0 mem_left_track_25.DFFR_2_.Q
rlabel metal3 34272 22232 34272 22232 0 mem_left_track_25.DFFR_3_.Q
rlabel metal3 38248 22568 38248 22568 0 mem_left_track_25.DFFR_4_.Q
rlabel metal2 32984 23408 32984 23408 0 mem_left_track_25.DFFR_5_.Q
rlabel metal2 42840 22960 42840 22960 0 mem_left_track_33.DFFR_0_.Q
rlabel metal3 40544 21336 40544 21336 0 mem_left_track_33.DFFR_1_.Q
rlabel metal3 41720 21672 41720 21672 0 mem_left_track_33.DFFR_2_.Q
rlabel metal2 40600 21392 40600 21392 0 mem_left_track_33.DFFR_3_.Q
rlabel metal3 42224 15400 42224 15400 0 mem_left_track_33.DFFR_4_.Q
rlabel metal2 14952 23184 14952 23184 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 20776 16688 20776 16688 0 mem_left_track_9.DFFR_1_.Q
rlabel metal2 21616 13832 21616 13832 0 mem_left_track_9.DFFR_2_.Q
rlabel metal2 22568 17696 22568 17696 0 mem_left_track_9.DFFR_3_.Q
rlabel metal2 31976 18984 31976 18984 0 mem_left_track_9.DFFR_4_.Q
rlabel metal2 5320 29848 5320 29848 0 mem_right_track_0.DFFR_0_.Q
rlabel metal2 2072 25144 2072 25144 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 2744 27272 2744 27272 0 mem_right_track_0.DFFR_2_.Q
rlabel metal2 7672 27104 7672 27104 0 mem_right_track_0.DFFR_3_.Q
rlabel metal2 9240 28672 9240 28672 0 mem_right_track_0.DFFR_4_.Q
rlabel metal2 7000 25032 7000 25032 0 mem_right_track_0.DFFR_5_.Q
rlabel metal2 13160 25704 13160 25704 0 mem_right_track_0.DFFR_6_.Q
rlabel metal2 13272 25144 13272 25144 0 mem_right_track_0.DFFR_7_.Q
rlabel metal2 15288 28280 15288 28280 0 mem_right_track_16.DFFR_0_.D
rlabel metal3 19096 30072 19096 30072 0 mem_right_track_16.DFFR_0_.Q
rlabel metal2 23576 27832 23576 27832 0 mem_right_track_16.DFFR_1_.Q
rlabel metal2 16408 28840 16408 28840 0 mem_right_track_16.DFFR_2_.Q
rlabel metal2 21224 29624 21224 29624 0 mem_right_track_16.DFFR_3_.Q
rlabel metal3 23744 30072 23744 30072 0 mem_right_track_16.DFFR_4_.Q
rlabel metal2 24808 29848 24808 29848 0 mem_right_track_16.DFFR_5_.Q
rlabel metal2 27832 28840 27832 28840 0 mem_right_track_24.DFFR_0_.Q
rlabel metal2 35336 29344 35336 29344 0 mem_right_track_24.DFFR_1_.Q
rlabel metal2 32760 29960 32760 29960 0 mem_right_track_24.DFFR_2_.Q
rlabel metal2 31528 26488 31528 26488 0 mem_right_track_24.DFFR_3_.Q
rlabel metal2 23352 25144 23352 25144 0 mem_right_track_24.DFFR_4_.Q
rlabel metal2 24808 26488 24808 26488 0 mem_right_track_24.DFFR_5_.Q
rlabel metal2 27384 28112 27384 28112 0 mem_right_track_32.DFFR_0_.Q
rlabel metal2 28840 26488 28840 26488 0 mem_right_track_32.DFFR_1_.Q
rlabel metal2 32088 27328 32088 27328 0 mem_right_track_32.DFFR_2_.Q
rlabel metal2 32648 29064 32648 29064 0 mem_right_track_32.DFFR_3_.Q
rlabel metal2 34216 28392 34216 28392 0 mem_right_track_32.DFFR_4_.Q
rlabel metal2 19880 26040 19880 26040 0 mem_right_track_8.DFFR_0_.Q
rlabel metal2 17248 31080 17248 31080 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 5488 25704 5488 25704 0 mem_right_track_8.DFFR_2_.Q
rlabel metal2 11592 30240 11592 30240 0 mem_right_track_8.DFFR_3_.Q
rlabel metal2 13048 28392 13048 28392 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 2072 28728 2072 28728 0 net1
rlabel metal2 20776 6468 20776 6468 0 net10
rlabel metal3 21784 15960 21784 15960 0 net100
rlabel metal2 19768 14868 19768 14868 0 net101
rlabel metal2 9912 22680 9912 22680 0 net102
rlabel metal2 19992 27720 19992 27720 0 net103
rlabel metal2 9912 16800 9912 16800 0 net104
rlabel metal2 15120 28728 15120 28728 0 net105
rlabel metal2 21784 29848 21784 29848 0 net106
rlabel metal2 19096 23072 19096 23072 0 net107
rlabel metal2 23688 21112 23688 21112 0 net108
rlabel metal2 8456 16520 8456 16520 0 net109
rlabel metal2 27160 6384 27160 6384 0 net11
rlabel metal2 8568 21616 8568 21616 0 net110
rlabel metal2 14952 29736 14952 29736 0 net111
rlabel metal2 32536 13272 32536 13272 0 net112
rlabel metal3 22344 25592 22344 25592 0 net113
rlabel metal2 31192 27888 31192 27888 0 net114
rlabel metal2 37464 23856 37464 23856 0 net115
rlabel metal2 12040 22288 12040 22288 0 net116
rlabel metal2 32200 19544 32200 19544 0 net117
rlabel metal2 38472 20832 38472 20832 0 net118
rlabel metal2 15960 23240 15960 23240 0 net119
rlabel metal2 43848 7112 43848 7112 0 net12
rlabel metal2 34888 21672 34888 21672 0 net120
rlabel metal2 36008 17696 36008 17696 0 net121
rlabel metal2 15400 22008 15400 22008 0 net122
rlabel metal3 31220 22344 31220 22344 0 net123
rlabel metal2 36008 29344 36008 29344 0 net124
rlabel metal2 12992 18424 12992 18424 0 net125
rlabel metal2 12376 23128 12376 23128 0 net126
rlabel metal3 18648 15848 18648 15848 0 net127
rlabel metal2 32200 17360 32200 17360 0 net128
rlabel metal3 5824 21560 5824 21560 0 net129
rlabel metal2 21448 36960 21448 36960 0 net13
rlabel metal3 6244 24024 6244 24024 0 net130
rlabel metal2 36008 19376 36008 19376 0 net131
rlabel metal2 10136 14952 10136 14952 0 net132
rlabel metal2 14840 14448 14840 14448 0 net133
rlabel metal2 10808 15344 10808 15344 0 net134
rlabel metal2 21840 14840 21840 14840 0 net135
rlabel metal2 24696 29456 24696 29456 0 net136
rlabel metal3 16856 25536 16856 25536 0 net137
rlabel metal2 29736 28952 29736 28952 0 net138
rlabel metal2 16800 16408 16800 16408 0 net139
rlabel metal2 26264 37128 26264 37128 0 net14
rlabel metal2 40040 15568 40040 15568 0 net140
rlabel metal3 25032 25592 25032 25592 0 net141
rlabel metal2 33544 24472 33544 24472 0 net142
rlabel metal2 29624 16576 29624 16576 0 net143
rlabel metal2 37464 16520 37464 16520 0 net144
rlabel metal2 18760 13580 18760 13580 0 net145
rlabel metal2 7448 15344 7448 15344 0 net146
rlabel metal2 4088 21392 4088 21392 0 net147
rlabel metal2 37576 21896 37576 21896 0 net148
rlabel metal2 37576 27384 37576 27384 0 net149
rlabel metal2 36456 4816 36456 4816 0 net15
rlabel metal2 26992 29400 26992 29400 0 net150
rlabel metal2 38808 24752 38808 24752 0 net151
rlabel metal2 28392 15288 28392 15288 0 net152
rlabel metal3 21252 28728 21252 28728 0 net153
rlabel metal2 35672 14728 35672 14728 0 net154
rlabel metal2 29736 23240 29736 23240 0 net155
rlabel metal2 12264 28560 12264 28560 0 net156
rlabel metal2 2744 14728 2744 14728 0 net157
rlabel metal2 29736 15344 29736 15344 0 net158
rlabel metal2 40040 13776 40040 13776 0 net159
rlabel metal3 37576 40488 37576 40488 0 net16
rlabel metal2 33544 15176 33544 15176 0 net160
rlabel metal2 37576 28672 37576 28672 0 net161
rlabel metal3 24752 14056 24752 14056 0 net162
rlabel metal2 8008 22960 8008 22960 0 net163
rlabel metal2 33544 28728 33544 28728 0 net164
rlabel metal2 20328 31416 20328 31416 0 net165
rlabel metal2 6216 28168 6216 28168 0 net166
rlabel metal2 25816 28560 25816 28560 0 net167
rlabel metal2 27832 13384 27832 13384 0 net168
rlabel metal2 18032 29400 18032 29400 0 net169
rlabel metal2 18536 40712 18536 40712 0 net17
rlabel metal2 15512 18480 15512 18480 0 net170
rlabel metal3 11704 30296 11704 30296 0 net171
rlabel metal2 2744 17472 2744 17472 0 net172
rlabel metal2 8008 18704 8008 18704 0 net173
rlabel metal2 4760 16912 4760 16912 0 net174
rlabel metal2 23912 12992 23912 12992 0 net175
rlabel metal3 4144 17752 4144 17752 0 net176
rlabel metal2 3976 19264 3976 19264 0 net177
rlabel metal2 4088 26712 4088 26712 0 net178
rlabel metal2 33656 15904 33656 15904 0 net179
rlabel metal2 14840 41272 14840 41272 0 net18
rlabel metal2 10024 28224 10024 28224 0 net180
rlabel metal2 39816 18872 39816 18872 0 net181
rlabel metal2 24360 19544 24360 19544 0 net182
rlabel metal2 36120 23072 36120 23072 0 net183
rlabel metal2 27608 22008 27608 22008 0 net184
rlabel metal2 29512 28448 29512 28448 0 net185
rlabel metal3 29176 16856 29176 16856 0 net186
rlabel metal2 8008 24640 8008 24640 0 net187
rlabel metal2 17976 18816 17976 18816 0 net188
rlabel metal2 37464 26992 37464 26992 0 net189
rlabel metal2 24136 38360 24136 38360 0 net19
rlabel metal3 24304 24024 24304 24024 0 net190
rlabel metal2 25704 12488 25704 12488 0 net191
rlabel metal2 3864 26712 3864 26712 0 net192
rlabel metal2 8008 28168 8008 28168 0 net193
rlabel metal2 23016 17192 23016 17192 0 net194
rlabel metal3 28812 21448 28812 21448 0 net195
rlabel metal2 34552 26544 34552 26544 0 net196
rlabel metal2 38248 26320 38248 26320 0 net197
rlabel metal2 16408 27776 16408 27776 0 net198
rlabel metal2 27048 24920 27048 24920 0 net199
rlabel metal2 43848 4592 43848 4592 0 net2
rlabel metal3 40432 39592 40432 39592 0 net20
rlabel metal2 5208 27496 5208 27496 0 net200
rlabel metal2 37576 17192 37576 17192 0 net201
rlabel metal2 33992 19544 33992 19544 0 net202
rlabel metal2 2968 14952 2968 14952 0 net203
rlabel metal2 13944 16912 13944 16912 0 net204
rlabel metal2 8680 25760 8680 25760 0 net205
rlabel metal2 19768 22288 19768 22288 0 net206
rlabel metal2 29960 25312 29960 25312 0 net207
rlabel metal2 19824 40376 19824 40376 0 net21
rlabel metal2 24024 4984 24024 4984 0 net22
rlabel metal2 43848 3808 43848 3808 0 net23
rlabel metal2 43848 41328 43848 41328 0 net24
rlabel metal3 38360 39592 38360 39592 0 net25
rlabel metal2 39816 40712 39816 40712 0 net26
rlabel metal2 25592 38304 25592 38304 0 net27
rlabel metal2 43848 39256 43848 39256 0 net28
rlabel metal2 19880 4536 19880 4536 0 net29
rlabel metal3 15008 40488 15008 40488 0 net3
rlabel metal2 38024 4368 38024 4368 0 net30
rlabel metal2 43176 39144 43176 39144 0 net31
rlabel metal2 37128 4816 37128 4816 0 net32
rlabel metal2 42504 31024 42504 31024 0 net33
rlabel metal2 43792 37912 43792 37912 0 net34
rlabel metal2 40936 4760 40936 4760 0 net35
rlabel metal2 32984 40488 32984 40488 0 net36
rlabel metal2 11536 16072 11536 16072 0 net37
rlabel metal2 42952 21896 42952 21896 0 net38
rlabel metal2 33432 41272 33432 41272 0 net39
rlabel metal2 43120 4424 43120 4424 0 net4
rlabel metal2 24528 35896 24528 35896 0 net40
rlabel metal2 19656 40600 19656 40600 0 net41
rlabel metal2 25256 3920 25256 3920 0 net42
rlabel metal2 42504 6608 42504 6608 0 net43
rlabel metal2 39480 39816 39480 39816 0 net44
rlabel metal2 39480 41272 39480 41272 0 net45
rlabel metal2 25816 37408 25816 37408 0 net46
rlabel metal2 15176 40880 15176 40880 0 net47
rlabel metal2 42504 40320 42504 40320 0 net48
rlabel metal2 20216 4592 20216 4592 0 net49
rlabel metal2 25200 4536 25200 4536 0 net5
rlabel metal2 42616 40880 42616 40880 0 net50
rlabel metal2 37240 4200 37240 4200 0 net51
rlabel metal2 42728 31472 42728 31472 0 net52
rlabel metal3 40712 3416 40712 3416 0 net53
rlabel metal2 18872 40768 18872 40768 0 net54
rlabel metal2 15848 41272 15848 41272 0 net55
rlabel metal2 41832 5432 41832 5432 0 net56
rlabel metal2 26152 4200 26152 4200 0 net57
rlabel metal2 39144 4200 39144 4200 0 net58
rlabel metal2 20832 35896 20832 35896 0 net59
rlabel metal2 38864 4536 38864 4536 0 net6
rlabel metal2 33880 4200 33880 4200 0 net60
rlabel metal2 32144 3528 32144 3528 0 net61
rlabel metal2 42840 6216 42840 6216 0 net62
rlabel metal2 21112 5964 21112 5964 0 net63
rlabel metal2 28392 5768 28392 5768 0 net64
rlabel metal3 22064 35896 22064 35896 0 net65
rlabel metal3 26824 35896 26824 35896 0 net66
rlabel metal2 37912 5096 37912 5096 0 net67
rlabel metal2 39144 40432 39144 40432 0 net68
rlabel metal2 42168 39424 42168 39424 0 net69
rlabel metal2 20552 38304 20552 38304 0 net7
rlabel metal2 40152 40152 40152 40152 0 net70
rlabel metal3 42448 40488 42448 40488 0 net71
rlabel metal3 39032 3528 39032 3528 0 net72
rlabel metal2 43512 5824 43512 5824 0 net73
rlabel metal2 24920 44478 24920 44478 0 net74
rlabel metal2 21560 2030 21560 2030 0 net75
rlabel metal3 44478 37688 44478 37688 0 net76
rlabel metal3 44506 36344 44506 36344 0 net77
rlabel metal2 26264 910 26264 910 0 net78
rlabel metal2 16856 44478 16856 44478 0 net79
rlabel metal2 33544 4816 33544 4816 0 net8
rlabel metal2 31640 44478 31640 44478 0 net80
rlabel metal2 42896 4536 42896 4536 0 net81
rlabel metal3 44478 38360 44478 38360 0 net82
rlabel metal3 43834 39032 43834 39032 0 net83
rlabel metal2 40376 40096 40376 40096 0 net84
rlabel metal3 44478 40376 44478 40376 0 net85
rlabel metal2 39704 2590 39704 2590 0 net86
rlabel metal2 44240 36232 44240 36232 0 net87
rlabel metal2 36344 44478 36344 44478 0 net88
rlabel metal2 41048 44478 41048 44478 0 net89
rlabel metal2 31528 4200 31528 4200 0 net9
rlabel metal2 30968 44478 30968 44478 0 net90
rlabel metal2 37016 2030 37016 2030 0 net91
rlabel metal2 42392 4256 42392 4256 0 net92
rlabel metal2 44184 37184 44184 37184 0 net93
rlabel metal2 41720 44478 41720 44478 0 net94
rlabel metal2 32368 4424 32368 4424 0 net95
rlabel metal2 42616 7168 42616 7168 0 net96
rlabel metal2 34328 44478 34328 44478 0 net97
rlabel metal3 44478 35000 44478 35000 0 net98
rlabel metal3 23576 13608 23576 13608 0 net99
rlabel metal2 1736 18928 1736 18928 0 pReset
rlabel metal3 2198 28952 2198 28952 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
