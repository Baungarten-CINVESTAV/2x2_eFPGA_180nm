magic
tech gf180mcuD
magscale 1 10
timestamp 1702149601
<< metal1 >>
rect 22194 37214 22206 37266
rect 22258 37263 22270 37266
rect 23090 37263 23102 37266
rect 22258 37217 23102 37263
rect 22258 37214 22270 37217
rect 23090 37214 23102 37217
rect 23154 37214 23166 37266
rect 1344 36874 38640 36908
rect 1344 36822 5876 36874
rect 5928 36822 5980 36874
rect 6032 36822 6084 36874
rect 6136 36822 15200 36874
rect 15252 36822 15304 36874
rect 15356 36822 15408 36874
rect 15460 36822 24524 36874
rect 24576 36822 24628 36874
rect 24680 36822 24732 36874
rect 24784 36822 33848 36874
rect 33900 36822 33952 36874
rect 34004 36822 34056 36874
rect 34108 36822 38640 36874
rect 1344 36788 38640 36822
rect 37774 36706 37826 36718
rect 29362 36654 29374 36706
rect 29426 36703 29438 36706
rect 29698 36703 29710 36706
rect 29426 36657 29710 36703
rect 29426 36654 29438 36657
rect 29698 36654 29710 36657
rect 29762 36654 29774 36706
rect 37774 36642 37826 36654
rect 19506 36542 19518 36594
rect 19570 36542 19582 36594
rect 21298 36542 21310 36594
rect 21362 36542 21374 36594
rect 23090 36542 23102 36594
rect 23154 36542 23166 36594
rect 26114 36542 26126 36594
rect 26178 36542 26190 36594
rect 28802 36542 28814 36594
rect 28866 36542 28878 36594
rect 32610 36542 32622 36594
rect 32674 36542 32686 36594
rect 34402 36542 34414 36594
rect 34466 36542 34478 36594
rect 29710 36482 29762 36494
rect 17714 36430 17726 36482
rect 17778 36430 17790 36482
rect 18386 36430 18398 36482
rect 18450 36430 18462 36482
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 22194 36430 22206 36482
rect 22258 36430 22270 36482
rect 25666 36430 25678 36482
rect 25730 36430 25742 36482
rect 30706 36430 30718 36482
rect 30770 36430 30782 36482
rect 29710 36418 29762 36430
rect 26686 36370 26738 36382
rect 26686 36306 26738 36318
rect 27134 36370 27186 36382
rect 27134 36306 27186 36318
rect 29934 36370 29986 36382
rect 29934 36306 29986 36318
rect 31614 36370 31666 36382
rect 31614 36306 31666 36318
rect 35310 36370 35362 36382
rect 35310 36306 35362 36318
rect 36206 36370 36258 36382
rect 36206 36306 36258 36318
rect 17950 36258 18002 36270
rect 17950 36194 18002 36206
rect 18622 36258 18674 36270
rect 18622 36194 18674 36206
rect 22654 36258 22706 36270
rect 22654 36194 22706 36206
rect 27470 36258 27522 36270
rect 27470 36194 27522 36206
rect 28366 36258 28418 36270
rect 28366 36194 28418 36206
rect 30494 36258 30546 36270
rect 30494 36194 30546 36206
rect 32174 36258 32226 36270
rect 32174 36194 32226 36206
rect 33742 36258 33794 36270
rect 33742 36194 33794 36206
rect 36542 36258 36594 36270
rect 36542 36194 36594 36206
rect 36990 36258 37042 36270
rect 36990 36194 37042 36206
rect 1344 36090 38800 36124
rect 1344 36038 10538 36090
rect 10590 36038 10642 36090
rect 10694 36038 10746 36090
rect 10798 36038 19862 36090
rect 19914 36038 19966 36090
rect 20018 36038 20070 36090
rect 20122 36038 29186 36090
rect 29238 36038 29290 36090
rect 29342 36038 29394 36090
rect 29446 36038 38510 36090
rect 38562 36038 38614 36090
rect 38666 36038 38718 36090
rect 38770 36038 38800 36090
rect 1344 36004 38800 36038
rect 18174 35922 18226 35934
rect 18174 35858 18226 35870
rect 18846 35922 18898 35934
rect 18846 35858 18898 35870
rect 20190 35922 20242 35934
rect 20190 35858 20242 35870
rect 20526 35922 20578 35934
rect 20526 35858 20578 35870
rect 21534 35922 21586 35934
rect 21534 35858 21586 35870
rect 22206 35922 22258 35934
rect 22206 35858 22258 35870
rect 22542 35922 22594 35934
rect 22542 35858 22594 35870
rect 28702 35922 28754 35934
rect 28702 35858 28754 35870
rect 28926 35922 28978 35934
rect 28926 35858 28978 35870
rect 29822 35922 29874 35934
rect 29822 35858 29874 35870
rect 30718 35922 30770 35934
rect 30718 35858 30770 35870
rect 31950 35922 32002 35934
rect 31950 35858 32002 35870
rect 19854 35810 19906 35822
rect 19854 35746 19906 35758
rect 21198 35810 21250 35822
rect 21198 35746 21250 35758
rect 21870 35810 21922 35822
rect 21870 35746 21922 35758
rect 23102 35810 23154 35822
rect 23102 35746 23154 35758
rect 23438 35810 23490 35822
rect 23438 35746 23490 35758
rect 23774 35810 23826 35822
rect 23774 35746 23826 35758
rect 24110 35810 24162 35822
rect 24110 35746 24162 35758
rect 34750 35810 34802 35822
rect 34750 35746 34802 35758
rect 35086 35810 35138 35822
rect 35086 35746 35138 35758
rect 27358 35698 27410 35710
rect 31614 35698 31666 35710
rect 20738 35646 20750 35698
rect 20802 35646 20814 35698
rect 26786 35646 26798 35698
rect 26850 35646 26862 35698
rect 29138 35646 29150 35698
rect 29202 35646 29214 35698
rect 30482 35646 30494 35698
rect 30546 35646 30558 35698
rect 27358 35634 27410 35646
rect 31614 35634 31666 35646
rect 33182 35698 33234 35710
rect 33182 35634 33234 35646
rect 34526 35698 34578 35710
rect 35410 35646 35422 35698
rect 35474 35646 35486 35698
rect 37090 35646 37102 35698
rect 37154 35646 37166 35698
rect 34526 35634 34578 35646
rect 26002 35534 26014 35586
rect 26066 35534 26078 35586
rect 27794 35534 27806 35586
rect 27858 35534 27870 35586
rect 33618 35534 33630 35586
rect 33682 35534 33694 35586
rect 36418 35534 36430 35586
rect 36482 35534 36494 35586
rect 37774 35474 37826 35486
rect 37774 35410 37826 35422
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 35646 35138 35698 35150
rect 35646 35074 35698 35086
rect 20414 35026 20466 35038
rect 20414 34962 20466 34974
rect 22878 35026 22930 35038
rect 22878 34962 22930 34974
rect 23550 35026 23602 35038
rect 23550 34962 23602 34974
rect 24222 35026 24274 35038
rect 37650 34974 37662 35026
rect 37714 34974 37726 35026
rect 24222 34962 24274 34974
rect 24446 34914 24498 34926
rect 24446 34850 24498 34862
rect 25342 34914 25394 34926
rect 36990 34914 37042 34926
rect 26114 34862 26126 34914
rect 26178 34862 26190 34914
rect 32386 34862 32398 34914
rect 32450 34862 32462 34914
rect 25342 34850 25394 34862
rect 36990 34850 37042 34862
rect 24782 34802 24834 34814
rect 24782 34738 24834 34750
rect 25678 34802 25730 34814
rect 25678 34738 25730 34750
rect 26350 34802 26402 34814
rect 26350 34738 26402 34750
rect 26686 34802 26738 34814
rect 26686 34738 26738 34750
rect 27022 34802 27074 34814
rect 27022 34738 27074 34750
rect 32622 34802 32674 34814
rect 32622 34738 32674 34750
rect 33518 34802 33570 34814
rect 33518 34738 33570 34750
rect 33966 34802 34018 34814
rect 33966 34738 34018 34750
rect 34302 34802 34354 34814
rect 34302 34738 34354 34750
rect 34974 34802 35026 34814
rect 34974 34738 35026 34750
rect 35310 34802 35362 34814
rect 35310 34738 35362 34750
rect 34638 34690 34690 34702
rect 34638 34626 34690 34638
rect 36430 34690 36482 34702
rect 36430 34626 36482 34638
rect 1344 34522 38800 34556
rect 1344 34470 10538 34522
rect 10590 34470 10642 34522
rect 10694 34470 10746 34522
rect 10798 34470 19862 34522
rect 19914 34470 19966 34522
rect 20018 34470 20070 34522
rect 20122 34470 29186 34522
rect 29238 34470 29290 34522
rect 29342 34470 29394 34522
rect 29446 34470 38510 34522
rect 38562 34470 38614 34522
rect 38666 34470 38718 34522
rect 38770 34470 38800 34522
rect 1344 34436 38800 34470
rect 33630 34354 33682 34366
rect 33630 34290 33682 34302
rect 34750 34354 34802 34366
rect 34750 34290 34802 34302
rect 34078 34242 34130 34254
rect 34078 34178 34130 34190
rect 35422 34242 35474 34254
rect 36978 34190 36990 34242
rect 37042 34190 37054 34242
rect 35422 34178 35474 34190
rect 34414 34130 34466 34142
rect 34414 34066 34466 34078
rect 35086 34130 35138 34142
rect 35086 34066 35138 34078
rect 35970 33966 35982 34018
rect 36034 33966 36046 34018
rect 1344 33738 38640 33772
rect 1344 33686 5876 33738
rect 5928 33686 5980 33738
rect 6032 33686 6084 33738
rect 6136 33686 15200 33738
rect 15252 33686 15304 33738
rect 15356 33686 15408 33738
rect 15460 33686 24524 33738
rect 24576 33686 24628 33738
rect 24680 33686 24732 33738
rect 24784 33686 33848 33738
rect 33900 33686 33952 33738
rect 34004 33686 34056 33738
rect 34108 33686 38640 33738
rect 1344 33652 38640 33686
rect 38222 33458 38274 33470
rect 35298 33406 35310 33458
rect 35362 33406 35374 33458
rect 37538 33406 37550 33458
rect 37602 33406 37614 33458
rect 38222 33394 38274 33406
rect 37090 33294 37102 33346
rect 37154 33294 37166 33346
rect 34066 33182 34078 33234
rect 34130 33182 34142 33234
rect 1344 32954 38800 32988
rect 1344 32902 10538 32954
rect 10590 32902 10642 32954
rect 10694 32902 10746 32954
rect 10798 32902 19862 32954
rect 19914 32902 19966 32954
rect 20018 32902 20070 32954
rect 20122 32902 29186 32954
rect 29238 32902 29290 32954
rect 29342 32902 29394 32954
rect 29446 32902 38510 32954
rect 38562 32902 38614 32954
rect 38666 32902 38718 32954
rect 38770 32902 38800 32954
rect 1344 32868 38800 32902
rect 34974 32786 35026 32798
rect 34974 32722 35026 32734
rect 37662 32786 37714 32798
rect 37662 32722 37714 32734
rect 38222 32786 38274 32798
rect 38222 32722 38274 32734
rect 35422 32674 35474 32686
rect 36978 32622 36990 32674
rect 37042 32622 37054 32674
rect 35422 32610 35474 32622
rect 35746 32398 35758 32450
rect 35810 32398 35822 32450
rect 1344 32170 38640 32204
rect 1344 32118 5876 32170
rect 5928 32118 5980 32170
rect 6032 32118 6084 32170
rect 6136 32118 15200 32170
rect 15252 32118 15304 32170
rect 15356 32118 15408 32170
rect 15460 32118 24524 32170
rect 24576 32118 24628 32170
rect 24680 32118 24732 32170
rect 24784 32118 33848 32170
rect 33900 32118 33952 32170
rect 34004 32118 34056 32170
rect 34108 32118 38640 32170
rect 1344 32084 38640 32118
rect 34290 31838 34302 31890
rect 34354 31838 34366 31890
rect 36194 31726 36206 31778
rect 36258 31726 36270 31778
rect 37314 31726 37326 31778
rect 37378 31726 37390 31778
rect 36430 31666 36482 31678
rect 35298 31614 35310 31666
rect 35362 31614 35374 31666
rect 36430 31602 36482 31614
rect 37886 31666 37938 31678
rect 37886 31602 37938 31614
rect 38222 31666 38274 31678
rect 38222 31602 38274 31614
rect 37550 31554 37602 31566
rect 37550 31490 37602 31502
rect 1344 31386 38800 31420
rect 1344 31334 10538 31386
rect 10590 31334 10642 31386
rect 10694 31334 10746 31386
rect 10798 31334 19862 31386
rect 19914 31334 19966 31386
rect 20018 31334 20070 31386
rect 20122 31334 29186 31386
rect 29238 31334 29290 31386
rect 29342 31334 29394 31386
rect 29446 31334 38510 31386
rect 38562 31334 38614 31386
rect 38666 31334 38718 31386
rect 38770 31334 38800 31386
rect 1344 31300 38800 31334
rect 36430 31218 36482 31230
rect 36430 31154 36482 31166
rect 36878 31218 36930 31230
rect 36878 31154 36930 31166
rect 37214 31218 37266 31230
rect 37214 31154 37266 31166
rect 37886 31218 37938 31230
rect 37886 31154 37938 31166
rect 38222 31106 38274 31118
rect 35410 31054 35422 31106
rect 35474 31054 35486 31106
rect 38222 31042 38274 31054
rect 37426 30942 37438 30994
rect 37490 30942 37502 30994
rect 34402 30830 34414 30882
rect 34466 30830 34478 30882
rect 1344 30602 38640 30636
rect 1344 30550 5876 30602
rect 5928 30550 5980 30602
rect 6032 30550 6084 30602
rect 6136 30550 15200 30602
rect 15252 30550 15304 30602
rect 15356 30550 15408 30602
rect 15460 30550 24524 30602
rect 24576 30550 24628 30602
rect 24680 30550 24732 30602
rect 24784 30550 33848 30602
rect 33900 30550 33952 30602
rect 34004 30550 34056 30602
rect 34108 30550 38640 30602
rect 1344 30516 38640 30550
rect 10434 30270 10446 30322
rect 10498 30270 10510 30322
rect 14466 30270 14478 30322
rect 14530 30270 14542 30322
rect 31042 30270 31054 30322
rect 31106 30270 31118 30322
rect 34962 30270 34974 30322
rect 35026 30270 35038 30322
rect 37102 30098 37154 30110
rect 11442 30046 11454 30098
rect 11506 30046 11518 30098
rect 15698 30046 15710 30098
rect 15762 30046 15774 30098
rect 32050 30046 32062 30098
rect 32114 30046 32126 30098
rect 36194 30046 36206 30098
rect 36258 30046 36270 30098
rect 37102 30034 37154 30046
rect 37550 30098 37602 30110
rect 37550 30034 37602 30046
rect 37886 30098 37938 30110
rect 37886 30034 37938 30046
rect 38222 30098 38274 30110
rect 38222 30034 38274 30046
rect 1344 29818 38800 29852
rect 1344 29766 10538 29818
rect 10590 29766 10642 29818
rect 10694 29766 10746 29818
rect 10798 29766 19862 29818
rect 19914 29766 19966 29818
rect 20018 29766 20070 29818
rect 20122 29766 29186 29818
rect 29238 29766 29290 29818
rect 29342 29766 29394 29818
rect 29446 29766 38510 29818
rect 38562 29766 38614 29818
rect 38666 29766 38718 29818
rect 38770 29766 38800 29818
rect 1344 29732 38800 29766
rect 36766 29650 36818 29662
rect 36766 29586 36818 29598
rect 37550 29650 37602 29662
rect 37550 29586 37602 29598
rect 37886 29650 37938 29662
rect 37886 29586 37938 29598
rect 13346 29486 13358 29538
rect 13410 29486 13422 29538
rect 16258 29486 16270 29538
rect 16322 29486 16334 29538
rect 29810 29486 29822 29538
rect 29874 29486 29886 29538
rect 35186 29486 35198 29538
rect 35250 29486 35262 29538
rect 38222 29426 38274 29438
rect 38222 29362 38274 29374
rect 37214 29314 37266 29326
rect 12338 29262 12350 29314
rect 12402 29262 12414 29314
rect 15250 29262 15262 29314
rect 15314 29262 15326 29314
rect 28466 29262 28478 29314
rect 28530 29262 28542 29314
rect 34066 29262 34078 29314
rect 34130 29262 34142 29314
rect 37214 29250 37266 29262
rect 1344 29034 38640 29068
rect 1344 28982 5876 29034
rect 5928 28982 5980 29034
rect 6032 28982 6084 29034
rect 6136 28982 15200 29034
rect 15252 28982 15304 29034
rect 15356 28982 15408 29034
rect 15460 28982 24524 29034
rect 24576 28982 24628 29034
rect 24680 28982 24732 29034
rect 24784 28982 33848 29034
rect 33900 28982 33952 29034
rect 34004 28982 34056 29034
rect 34108 28982 38640 29034
rect 1344 28948 38640 28982
rect 9650 28702 9662 28754
rect 9714 28702 9726 28754
rect 15250 28702 15262 28754
rect 15314 28702 15326 28754
rect 18050 28702 18062 28754
rect 18114 28702 18126 28754
rect 27010 28702 27022 28754
rect 27074 28702 27086 28754
rect 30146 28702 30158 28754
rect 30210 28702 30222 28754
rect 32946 28702 32958 28754
rect 33010 28702 33022 28754
rect 37662 28642 37714 28654
rect 38098 28590 38110 28642
rect 38162 28590 38174 28642
rect 37662 28578 37714 28590
rect 37886 28530 37938 28542
rect 10882 28478 10894 28530
rect 10946 28478 10958 28530
rect 16594 28478 16606 28530
rect 16658 28478 16670 28530
rect 19058 28478 19070 28530
rect 19122 28478 19134 28530
rect 28018 28478 28030 28530
rect 28082 28478 28094 28530
rect 31154 28478 31166 28530
rect 31218 28478 31230 28530
rect 34178 28478 34190 28530
rect 34242 28478 34254 28530
rect 37886 28466 37938 28478
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 37886 28082 37938 28094
rect 14690 28030 14702 28082
rect 14754 28030 14766 28082
rect 37886 28018 37938 28030
rect 15262 27970 15314 27982
rect 29374 27970 29426 27982
rect 7970 27918 7982 27970
rect 8034 27918 8046 27970
rect 19618 27918 19630 27970
rect 19682 27918 19694 27970
rect 22306 27918 22318 27970
rect 22370 27918 22382 27970
rect 15262 27906 15314 27918
rect 29374 27906 29426 27918
rect 30158 27970 30210 27982
rect 35298 27918 35310 27970
rect 35362 27918 35374 27970
rect 30158 27906 30210 27918
rect 11790 27858 11842 27870
rect 26686 27858 26738 27870
rect 38222 27858 38274 27870
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 27122 27806 27134 27858
rect 27186 27806 27198 27858
rect 32274 27806 32286 27858
rect 32338 27806 32350 27858
rect 11790 27794 11842 27806
rect 26686 27794 26738 27806
rect 38222 27794 38274 27806
rect 11006 27746 11058 27758
rect 37662 27746 37714 27758
rect 6962 27694 6974 27746
rect 7026 27694 7038 27746
rect 10658 27694 10670 27746
rect 10722 27694 10734 27746
rect 18610 27694 18622 27746
rect 18674 27694 18686 27746
rect 23426 27694 23438 27746
rect 23490 27694 23502 27746
rect 32050 27694 32062 27746
rect 32114 27694 32126 27746
rect 34290 27694 34302 27746
rect 34354 27694 34366 27746
rect 11006 27682 11058 27694
rect 37662 27682 37714 27694
rect 1344 27466 38640 27500
rect 1344 27414 5876 27466
rect 5928 27414 5980 27466
rect 6032 27414 6084 27466
rect 6136 27414 15200 27466
rect 15252 27414 15304 27466
rect 15356 27414 15408 27466
rect 15460 27414 24524 27466
rect 24576 27414 24628 27466
rect 24680 27414 24732 27466
rect 24784 27414 33848 27466
rect 33900 27414 33952 27466
rect 34004 27414 34056 27466
rect 34108 27414 38640 27466
rect 1344 27380 38640 27414
rect 12462 27298 12514 27310
rect 12462 27234 12514 27246
rect 18286 27298 18338 27310
rect 18286 27234 18338 27246
rect 26014 27298 26066 27310
rect 26014 27234 26066 27246
rect 30382 27298 30434 27310
rect 30382 27234 30434 27246
rect 7074 27134 7086 27186
rect 7138 27134 7150 27186
rect 29362 27134 29374 27186
rect 29426 27134 29438 27186
rect 8990 27074 9042 27086
rect 14590 27074 14642 27086
rect 22318 27074 22370 27086
rect 34078 27074 34130 27086
rect 9426 27022 9438 27074
rect 9490 27022 9502 27074
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 15250 27022 15262 27074
rect 15314 27022 15326 27074
rect 22978 27022 22990 27074
rect 23042 27022 23054 27074
rect 33506 27022 33518 27074
rect 33570 27022 33582 27074
rect 8990 27010 9042 27022
rect 14590 27010 14642 27022
rect 22318 27010 22370 27022
rect 34078 27010 34130 27022
rect 11678 26962 11730 26974
rect 18846 26962 18898 26974
rect 8082 26910 8094 26962
rect 8146 26910 8158 26962
rect 13458 26910 13470 26962
rect 13522 26910 13534 26962
rect 11678 26898 11730 26910
rect 18846 26898 18898 26910
rect 29150 26962 29202 26974
rect 29150 26898 29202 26910
rect 37774 26962 37826 26974
rect 37774 26898 37826 26910
rect 18958 26850 19010 26862
rect 36990 26850 37042 26862
rect 17490 26798 17502 26850
rect 17554 26798 17566 26850
rect 25442 26798 25454 26850
rect 25506 26798 25518 26850
rect 31154 26798 31166 26850
rect 31218 26798 31230 26850
rect 18958 26786 19010 26798
rect 36990 26786 37042 26798
rect 1344 26682 38800 26716
rect 1344 26630 10538 26682
rect 10590 26630 10642 26682
rect 10694 26630 10746 26682
rect 10798 26630 19862 26682
rect 19914 26630 19966 26682
rect 20018 26630 20070 26682
rect 20122 26630 29186 26682
rect 29238 26630 29290 26682
rect 29342 26630 29394 26682
rect 29446 26630 38510 26682
rect 38562 26630 38614 26682
rect 38666 26630 38718 26682
rect 38770 26630 38800 26682
rect 1344 26596 38800 26630
rect 9102 26514 9154 26526
rect 8306 26462 8318 26514
rect 8370 26462 8382 26514
rect 9102 26450 9154 26462
rect 16046 26514 16098 26526
rect 16046 26450 16098 26462
rect 16382 26514 16434 26526
rect 16382 26450 16434 26462
rect 21086 26514 21138 26526
rect 21086 26450 21138 26462
rect 28814 26514 28866 26526
rect 32622 26514 32674 26526
rect 31826 26462 31838 26514
rect 31890 26462 31902 26514
rect 28814 26450 28866 26462
rect 32622 26450 32674 26462
rect 32958 26514 33010 26526
rect 37886 26514 37938 26526
rect 33618 26462 33630 26514
rect 33682 26462 33694 26514
rect 32958 26450 33010 26462
rect 37886 26450 37938 26462
rect 2382 26402 2434 26414
rect 15262 26402 15314 26414
rect 21870 26402 21922 26414
rect 9762 26350 9774 26402
rect 9826 26350 9838 26402
rect 20402 26350 20414 26402
rect 20466 26350 20478 26402
rect 2382 26338 2434 26350
rect 15262 26338 15314 26350
rect 21870 26338 21922 26350
rect 28030 26402 28082 26414
rect 28030 26338 28082 26350
rect 37550 26402 37602 26414
rect 37550 26338 37602 26350
rect 38222 26402 38274 26414
rect 38222 26338 38274 26350
rect 5294 26290 5346 26302
rect 4610 26238 4622 26290
rect 4674 26238 4686 26290
rect 5294 26226 5346 26238
rect 5630 26290 5682 26302
rect 12574 26290 12626 26302
rect 25342 26290 25394 26302
rect 29150 26290 29202 26302
rect 36430 26290 36482 26302
rect 6066 26238 6078 26290
rect 6130 26238 6142 26290
rect 13010 26238 13022 26290
rect 13074 26238 13086 26290
rect 24210 26238 24222 26290
rect 24274 26238 24286 26290
rect 24658 26238 24670 26290
rect 24722 26238 24734 26290
rect 25778 26238 25790 26290
rect 25842 26238 25854 26290
rect 29586 26238 29598 26290
rect 29650 26238 29662 26290
rect 35970 26238 35982 26290
rect 36034 26238 36046 26290
rect 5630 26226 5682 26238
rect 12574 26226 12626 26238
rect 25342 26226 25394 26238
rect 29150 26226 29202 26238
rect 36430 26226 36482 26238
rect 16270 26178 16322 26190
rect 11106 26126 11118 26178
rect 11170 26126 11182 26178
rect 19394 26126 19406 26178
rect 19458 26126 19470 26178
rect 16270 26114 16322 26126
rect 1598 26066 1650 26078
rect 1598 26002 1650 26014
rect 1344 25898 38640 25932
rect 1344 25846 5876 25898
rect 5928 25846 5980 25898
rect 6032 25846 6084 25898
rect 6136 25846 15200 25898
rect 15252 25846 15304 25898
rect 15356 25846 15408 25898
rect 15460 25846 24524 25898
rect 24576 25846 24628 25898
rect 24680 25846 24732 25898
rect 24784 25846 33848 25898
rect 33900 25846 33952 25898
rect 34004 25846 34056 25898
rect 34108 25846 38640 25898
rect 1344 25812 38640 25846
rect 5518 25730 5570 25742
rect 5518 25666 5570 25678
rect 13022 25730 13074 25742
rect 13022 25666 13074 25678
rect 32734 25730 32786 25742
rect 32734 25666 32786 25678
rect 36542 25730 36594 25742
rect 36542 25666 36594 25678
rect 38334 25618 38386 25630
rect 3490 25566 3502 25618
rect 3554 25566 3566 25618
rect 14130 25566 14142 25618
rect 14194 25566 14206 25618
rect 15922 25566 15934 25618
rect 15986 25566 15998 25618
rect 22418 25566 22430 25618
rect 22482 25566 22494 25618
rect 25554 25566 25566 25618
rect 25618 25566 25630 25618
rect 27682 25566 27694 25618
rect 27746 25566 27758 25618
rect 38334 25554 38386 25566
rect 8990 25506 9042 25518
rect 8642 25454 8654 25506
rect 8706 25454 8718 25506
rect 8990 25442 9042 25454
rect 9326 25506 9378 25518
rect 17166 25506 17218 25518
rect 29262 25506 29314 25518
rect 33070 25506 33122 25518
rect 9986 25454 9998 25506
rect 10050 25454 10062 25506
rect 17826 25454 17838 25506
rect 17890 25454 17902 25506
rect 27458 25454 27470 25506
rect 27522 25454 27534 25506
rect 29698 25454 29710 25506
rect 29762 25454 29774 25506
rect 33394 25454 33406 25506
rect 33458 25454 33470 25506
rect 37202 25454 37214 25506
rect 37266 25454 37278 25506
rect 9326 25442 9378 25454
rect 17166 25442 17218 25454
rect 29262 25442 29314 25454
rect 33070 25442 33122 25454
rect 6302 25394 6354 25406
rect 2146 25342 2158 25394
rect 2210 25342 2222 25394
rect 6302 25330 6354 25342
rect 13806 25394 13858 25406
rect 20862 25394 20914 25406
rect 14914 25342 14926 25394
rect 14978 25342 14990 25394
rect 23538 25342 23550 25394
rect 23602 25342 23614 25394
rect 26562 25342 26574 25394
rect 26626 25342 26638 25394
rect 36978 25342 36990 25394
rect 37042 25342 37054 25394
rect 13806 25330 13858 25342
rect 20862 25330 20914 25342
rect 12450 25230 12462 25282
rect 12514 25230 12526 25282
rect 20178 25230 20190 25282
rect 20242 25230 20254 25282
rect 32050 25230 32062 25282
rect 32114 25230 32126 25282
rect 35970 25230 35982 25282
rect 36034 25230 36046 25282
rect 1344 25114 38800 25148
rect 1344 25062 10538 25114
rect 10590 25062 10642 25114
rect 10694 25062 10746 25114
rect 10798 25062 19862 25114
rect 19914 25062 19966 25114
rect 20018 25062 20070 25114
rect 20122 25062 29186 25114
rect 29238 25062 29290 25114
rect 29342 25062 29394 25114
rect 29446 25062 38510 25114
rect 38562 25062 38614 25114
rect 38666 25062 38718 25114
rect 38770 25062 38800 25114
rect 1344 25028 38800 25062
rect 8430 24946 8482 24958
rect 7858 24894 7870 24946
rect 7922 24894 7934 24946
rect 8430 24882 8482 24894
rect 15038 24946 15090 24958
rect 15038 24882 15090 24894
rect 18510 24946 18562 24958
rect 30158 24946 30210 24958
rect 29586 24894 29598 24946
rect 29650 24894 29662 24946
rect 18510 24882 18562 24894
rect 30158 24882 30210 24894
rect 30494 24946 30546 24958
rect 30494 24882 30546 24894
rect 38222 24946 38274 24958
rect 38222 24882 38274 24894
rect 14254 24834 14306 24846
rect 19294 24834 19346 24846
rect 37438 24834 37490 24846
rect 2258 24782 2270 24834
rect 2322 24782 2334 24834
rect 10098 24782 10110 24834
rect 10162 24782 10174 24834
rect 17490 24782 17502 24834
rect 17554 24782 17566 24834
rect 25218 24782 25230 24834
rect 25282 24782 25294 24834
rect 25890 24782 25902 24834
rect 25954 24782 25966 24834
rect 32050 24782 32062 24834
rect 32114 24782 32126 24834
rect 33170 24782 33182 24834
rect 33234 24782 33246 24834
rect 33954 24782 33966 24834
rect 34018 24782 34030 24834
rect 14254 24770 14306 24782
rect 19294 24770 19346 24782
rect 37438 24770 37490 24782
rect 4958 24722 5010 24734
rect 22206 24722 22258 24734
rect 5282 24670 5294 24722
rect 5346 24670 5358 24722
rect 10322 24670 10334 24722
rect 10386 24670 10398 24722
rect 10994 24670 11006 24722
rect 11058 24670 11070 24722
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 11890 24670 11902 24722
rect 11954 24670 11966 24722
rect 17714 24670 17726 24722
rect 17778 24670 17790 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 4958 24658 5010 24670
rect 22206 24658 22258 24670
rect 26686 24722 26738 24734
rect 34526 24722 34578 24734
rect 27122 24670 27134 24722
rect 27186 24670 27198 24722
rect 31826 24670 31838 24722
rect 31890 24670 31902 24722
rect 33394 24670 33406 24722
rect 33458 24670 33470 24722
rect 34178 24670 34190 24722
rect 34242 24670 34254 24722
rect 35186 24670 35198 24722
rect 35250 24670 35262 24722
rect 26686 24658 26738 24670
rect 34526 24658 34578 24670
rect 25566 24610 25618 24622
rect 3490 24558 3502 24610
rect 3554 24558 3566 24610
rect 10882 24558 10894 24610
rect 10946 24558 10958 24610
rect 25566 24546 25618 24558
rect 26238 24610 26290 24622
rect 26238 24546 26290 24558
rect 30382 24610 30434 24622
rect 30382 24546 30434 24558
rect 1344 24330 38640 24364
rect 1344 24278 5876 24330
rect 5928 24278 5980 24330
rect 6032 24278 6084 24330
rect 6136 24278 15200 24330
rect 15252 24278 15304 24330
rect 15356 24278 15408 24330
rect 15460 24278 24524 24330
rect 24576 24278 24628 24330
rect 24680 24278 24732 24330
rect 24784 24278 33848 24330
rect 33900 24278 33952 24330
rect 34004 24278 34056 24330
rect 34108 24278 38640 24330
rect 1344 24244 38640 24278
rect 9102 24162 9154 24174
rect 9102 24098 9154 24110
rect 19742 24162 19794 24174
rect 19742 24098 19794 24110
rect 36990 24050 37042 24062
rect 2258 23998 2270 24050
rect 2322 23998 2334 24050
rect 4050 23998 4062 24050
rect 4114 23998 4126 24050
rect 7634 23998 7646 24050
rect 7698 23998 7710 24050
rect 13458 23998 13470 24050
rect 13522 23998 13534 24050
rect 20178 23998 20190 24050
rect 20242 23998 20254 24050
rect 21298 23998 21310 24050
rect 21362 23998 21374 24050
rect 30146 23998 30158 24050
rect 30210 23998 30222 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 37314 23998 37326 24050
rect 37378 23998 37390 24050
rect 36990 23986 37042 23998
rect 12574 23938 12626 23950
rect 16046 23938 16098 23950
rect 12114 23886 12126 23938
rect 12178 23886 12190 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 16706 23886 16718 23938
rect 16770 23886 16782 23938
rect 20290 23886 20302 23938
rect 20354 23886 20366 23938
rect 21522 23886 21534 23938
rect 21586 23886 21598 23938
rect 23426 23886 23438 23938
rect 23490 23886 23502 23938
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 28242 23886 28254 23938
rect 28306 23886 28318 23938
rect 12574 23874 12626 23886
rect 16046 23874 16098 23886
rect 1934 23826 1986 23838
rect 5742 23826 5794 23838
rect 18958 23826 19010 23838
rect 27582 23826 27634 23838
rect 2930 23774 2942 23826
rect 2994 23774 3006 23826
rect 6626 23774 6638 23826
rect 6690 23774 6702 23826
rect 27234 23774 27246 23826
rect 27298 23774 27310 23826
rect 31154 23774 31166 23826
rect 31218 23774 31230 23826
rect 33954 23774 33966 23826
rect 34018 23774 34030 23826
rect 1934 23762 1986 23774
rect 5742 23762 5794 23774
rect 18958 23762 19010 23774
rect 27582 23762 27634 23774
rect 5854 23714 5906 23726
rect 27022 23714 27074 23726
rect 9874 23662 9886 23714
rect 9938 23662 9950 23714
rect 26450 23662 26462 23714
rect 26514 23662 26526 23714
rect 5854 23650 5906 23662
rect 27022 23650 27074 23662
rect 28254 23714 28306 23726
rect 28254 23650 28306 23662
rect 1344 23546 38800 23580
rect 1344 23494 10538 23546
rect 10590 23494 10642 23546
rect 10694 23494 10746 23546
rect 10798 23494 19862 23546
rect 19914 23494 19966 23546
rect 20018 23494 20070 23546
rect 20122 23494 29186 23546
rect 29238 23494 29290 23546
rect 29342 23494 29394 23546
rect 29446 23494 38510 23546
rect 38562 23494 38614 23546
rect 38666 23494 38718 23546
rect 38770 23494 38800 23546
rect 1344 23460 38800 23494
rect 2942 23378 2994 23390
rect 24782 23378 24834 23390
rect 36654 23378 36706 23390
rect 3714 23326 3726 23378
rect 3778 23326 3790 23378
rect 24210 23326 24222 23378
rect 24274 23326 24286 23378
rect 36082 23326 36094 23378
rect 36146 23326 36158 23378
rect 2942 23314 2994 23326
rect 24782 23314 24834 23326
rect 36654 23314 36706 23326
rect 6862 23266 6914 23278
rect 6862 23202 6914 23214
rect 7534 23266 7586 23278
rect 17726 23266 17778 23278
rect 7858 23214 7870 23266
rect 7922 23214 7934 23266
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 7534 23202 7586 23214
rect 17726 23202 17778 23214
rect 6414 23154 6466 23166
rect 21310 23154 21362 23166
rect 33182 23154 33234 23166
rect 5954 23102 5966 23154
rect 6018 23102 6030 23154
rect 14690 23102 14702 23154
rect 14754 23102 14766 23154
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 29362 23102 29374 23154
rect 29426 23102 29438 23154
rect 33618 23102 33630 23154
rect 33682 23102 33694 23154
rect 6414 23090 6466 23102
rect 21310 23090 21362 23102
rect 33182 23090 33234 23102
rect 15374 23042 15426 23054
rect 31390 23042 31442 23054
rect 7074 22990 7086 23042
rect 7138 22990 7150 23042
rect 10322 22990 10334 23042
rect 10386 22990 10398 23042
rect 17378 22990 17390 23042
rect 17442 22990 17454 23042
rect 19394 22990 19406 23042
rect 19458 22990 19470 23042
rect 26898 22990 26910 23042
rect 26962 22990 26974 23042
rect 15374 22978 15426 22990
rect 31390 22978 31442 22990
rect 1344 22762 38640 22796
rect 1344 22710 5876 22762
rect 5928 22710 5980 22762
rect 6032 22710 6084 22762
rect 6136 22710 15200 22762
rect 15252 22710 15304 22762
rect 15356 22710 15408 22762
rect 15460 22710 24524 22762
rect 24576 22710 24628 22762
rect 24680 22710 24732 22762
rect 24784 22710 33848 22762
rect 33900 22710 33952 22762
rect 34004 22710 34056 22762
rect 34108 22710 38640 22762
rect 1344 22676 38640 22710
rect 9326 22594 9378 22606
rect 9326 22530 9378 22542
rect 1934 22482 1986 22494
rect 29710 22482 29762 22494
rect 37662 22482 37714 22494
rect 4050 22430 4062 22482
rect 4114 22430 4126 22482
rect 16034 22430 16046 22482
rect 16098 22430 16110 22482
rect 26450 22430 26462 22482
rect 26514 22430 26526 22482
rect 28354 22430 28366 22482
rect 28418 22430 28430 22482
rect 33170 22430 33182 22482
rect 33234 22430 33246 22482
rect 36978 22430 36990 22482
rect 37042 22430 37054 22482
rect 1934 22418 1986 22430
rect 29710 22418 29762 22430
rect 37662 22418 37714 22430
rect 9214 22370 9266 22382
rect 12798 22370 12850 22382
rect 21758 22370 21810 22382
rect 8642 22318 8654 22370
rect 8706 22318 8718 22370
rect 12338 22318 12350 22370
rect 12402 22318 12414 22370
rect 15474 22318 15486 22370
rect 15538 22318 15550 22370
rect 20626 22318 20638 22370
rect 20690 22318 20702 22370
rect 22194 22318 22206 22370
rect 22258 22318 22270 22370
rect 29250 22318 29262 22370
rect 29314 22318 29326 22370
rect 31154 22318 31166 22370
rect 31218 22318 31230 22370
rect 37202 22318 37214 22370
rect 37266 22318 37278 22370
rect 9214 22306 9266 22318
rect 12798 22306 12850 22318
rect 21758 22306 21810 22318
rect 28590 22258 28642 22270
rect 2258 22206 2270 22258
rect 2322 22206 2334 22258
rect 3042 22206 3054 22258
rect 3106 22206 3118 22258
rect 20402 22206 20414 22258
rect 20466 22206 20478 22258
rect 27458 22206 27470 22258
rect 27522 22206 27534 22258
rect 28590 22194 28642 22206
rect 30830 22258 30882 22270
rect 30830 22194 30882 22206
rect 5518 22146 5570 22158
rect 19742 22146 19794 22158
rect 25230 22146 25282 22158
rect 6066 22094 6078 22146
rect 6130 22094 6142 22146
rect 10098 22094 10110 22146
rect 10162 22094 10174 22146
rect 24546 22094 24558 22146
rect 24610 22094 24622 22146
rect 5518 22082 5570 22094
rect 19742 22082 19794 22094
rect 25230 22082 25282 22094
rect 25566 22146 25618 22158
rect 25566 22082 25618 22094
rect 37774 22146 37826 22158
rect 37774 22082 37826 22094
rect 1344 21978 38800 22012
rect 1344 21926 10538 21978
rect 10590 21926 10642 21978
rect 10694 21926 10746 21978
rect 10798 21926 19862 21978
rect 19914 21926 19966 21978
rect 20018 21926 20070 21978
rect 20122 21926 29186 21978
rect 29238 21926 29290 21978
rect 29342 21926 29394 21978
rect 29446 21926 38510 21978
rect 38562 21926 38614 21978
rect 38666 21926 38718 21978
rect 38770 21926 38800 21978
rect 1344 21892 38800 21926
rect 1598 21810 1650 21822
rect 9662 21810 9714 21822
rect 22766 21810 22818 21822
rect 2258 21758 2270 21810
rect 2322 21758 2334 21810
rect 8530 21758 8542 21810
rect 8594 21758 8606 21810
rect 14018 21758 14030 21810
rect 14082 21758 14094 21810
rect 1598 21746 1650 21758
rect 9662 21746 9714 21758
rect 22766 21746 22818 21758
rect 24558 21810 24610 21822
rect 28814 21810 28866 21822
rect 38222 21810 38274 21822
rect 28242 21758 28254 21810
rect 28306 21758 28318 21810
rect 32050 21758 32062 21810
rect 32114 21758 32126 21810
rect 37650 21758 37662 21810
rect 37714 21758 37726 21810
rect 24558 21746 24610 21758
rect 28814 21746 28866 21758
rect 38222 21746 38274 21758
rect 9102 21698 9154 21710
rect 18510 21698 18562 21710
rect 12898 21646 12910 21698
rect 12962 21646 12974 21698
rect 9102 21634 9154 21646
rect 18510 21634 18562 21646
rect 21982 21698 22034 21710
rect 33406 21698 33458 21710
rect 33058 21646 33070 21698
rect 33122 21646 33134 21698
rect 21982 21634 22034 21646
rect 33406 21634 33458 21646
rect 33854 21698 33906 21710
rect 33854 21634 33906 21646
rect 5070 21586 5122 21598
rect 4722 21534 4734 21586
rect 4786 21534 4798 21586
rect 5070 21522 5122 21534
rect 5406 21586 5458 21598
rect 16718 21586 16770 21598
rect 19294 21586 19346 21598
rect 25342 21586 25394 21598
rect 28926 21586 28978 21598
rect 34526 21586 34578 21598
rect 5954 21534 5966 21586
rect 6018 21534 6030 21586
rect 16258 21534 16270 21586
rect 16322 21534 16334 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 19618 21534 19630 21586
rect 19682 21534 19694 21586
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 29586 21534 29598 21586
rect 29650 21534 29662 21586
rect 35186 21534 35198 21586
rect 35250 21534 35262 21586
rect 5406 21522 5458 21534
rect 16718 21522 16770 21534
rect 19294 21522 19346 21534
rect 25342 21522 25394 21534
rect 28926 21522 28978 21534
rect 34526 21522 34578 21534
rect 9550 21474 9602 21486
rect 24670 21474 24722 21486
rect 11554 21422 11566 21474
rect 11618 21422 11630 21474
rect 17602 21422 17614 21474
rect 17666 21422 17678 21474
rect 18722 21422 18734 21474
rect 18786 21422 18798 21474
rect 34178 21422 34190 21474
rect 34242 21422 34254 21474
rect 9550 21410 9602 21422
rect 24670 21410 24722 21422
rect 13246 21362 13298 21374
rect 13246 21298 13298 21310
rect 32622 21362 32674 21374
rect 32622 21298 32674 21310
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 6974 21026 7026 21038
rect 6974 20962 7026 20974
rect 11454 21026 11506 21038
rect 11454 20962 11506 20974
rect 12686 21026 12738 21038
rect 12686 20962 12738 20974
rect 19518 21026 19570 21038
rect 19518 20962 19570 20974
rect 34750 21026 34802 21038
rect 34750 20962 34802 20974
rect 13918 20914 13970 20926
rect 3826 20862 3838 20914
rect 3890 20862 3902 20914
rect 14242 20862 14254 20914
rect 14306 20862 14318 20914
rect 14578 20862 14590 20914
rect 14642 20862 14654 20914
rect 21746 20862 21758 20914
rect 21810 20862 21822 20914
rect 13918 20850 13970 20862
rect 5966 20802 6018 20814
rect 5966 20738 6018 20750
rect 7758 20802 7810 20814
rect 16046 20802 16098 20814
rect 26910 20802 26962 20814
rect 31054 20802 31106 20814
rect 8418 20750 8430 20802
rect 8482 20750 8494 20802
rect 11890 20750 11902 20802
rect 11954 20750 11966 20802
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 16370 20750 16382 20802
rect 16434 20750 16446 20802
rect 22306 20750 22318 20802
rect 22370 20750 22382 20802
rect 26562 20750 26574 20802
rect 26626 20750 26638 20802
rect 27570 20750 27582 20802
rect 27634 20750 27646 20802
rect 29810 20750 29822 20802
rect 29874 20750 29886 20802
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 7758 20738 7810 20750
rect 16046 20738 16098 20750
rect 26910 20738 26962 20750
rect 31054 20738 31106 20750
rect 18734 20690 18786 20702
rect 28590 20690 28642 20702
rect 34974 20690 35026 20702
rect 3042 20638 3054 20690
rect 3106 20638 3118 20690
rect 5618 20638 5630 20690
rect 5682 20638 5694 20690
rect 7522 20638 7534 20690
rect 7586 20638 7598 20690
rect 27346 20638 27358 20690
rect 27410 20638 27422 20690
rect 28242 20638 28254 20690
rect 28306 20638 28318 20690
rect 30370 20638 30382 20690
rect 30434 20638 30446 20690
rect 18734 20626 18786 20638
rect 28590 20626 28642 20638
rect 34974 20626 35026 20638
rect 13582 20578 13634 20590
rect 10882 20526 10894 20578
rect 10946 20526 10958 20578
rect 13582 20514 13634 20526
rect 22990 20578 23042 20590
rect 22990 20514 23042 20526
rect 23438 20578 23490 20590
rect 35086 20578 35138 20590
rect 24210 20526 24222 20578
rect 24274 20526 24286 20578
rect 34178 20526 34190 20578
rect 34242 20526 34254 20578
rect 23438 20514 23490 20526
rect 35086 20514 35138 20526
rect 38334 20578 38386 20590
rect 38334 20514 38386 20526
rect 1344 20410 38800 20444
rect 1344 20358 10538 20410
rect 10590 20358 10642 20410
rect 10694 20358 10746 20410
rect 10798 20358 19862 20410
rect 19914 20358 19966 20410
rect 20018 20358 20070 20410
rect 20122 20358 29186 20410
rect 29238 20358 29290 20410
rect 29342 20358 29394 20410
rect 29446 20358 38510 20410
rect 38562 20358 38614 20410
rect 38666 20358 38718 20410
rect 38770 20358 38800 20410
rect 1344 20324 38800 20358
rect 7074 20190 7086 20242
rect 7138 20190 7150 20242
rect 16370 20190 16382 20242
rect 16434 20190 16446 20242
rect 20402 20190 20414 20242
rect 20466 20190 20478 20242
rect 36754 20190 36766 20242
rect 36818 20190 36830 20242
rect 21310 20130 21362 20142
rect 26798 20130 26850 20142
rect 3826 20078 3838 20130
rect 3890 20078 3902 20130
rect 10994 20078 11006 20130
rect 11058 20078 11070 20130
rect 21634 20078 21646 20130
rect 21698 20078 21710 20130
rect 24210 20078 24222 20130
rect 24274 20078 24286 20130
rect 21310 20066 21362 20078
rect 26798 20066 26850 20078
rect 30606 20130 30658 20142
rect 38222 20130 38274 20142
rect 31938 20078 31950 20130
rect 32002 20078 32014 20130
rect 37874 20078 37886 20130
rect 37938 20078 37950 20130
rect 30606 20066 30658 20078
rect 38222 20066 38274 20078
rect 17278 20018 17330 20030
rect 29486 20018 29538 20030
rect 3602 19966 3614 20018
rect 3666 19966 3678 20018
rect 4162 19966 4174 20018
rect 4226 19966 4238 20018
rect 4722 19966 4734 20018
rect 4786 19966 4798 20018
rect 8082 19966 8094 20018
rect 8146 19966 8158 20018
rect 13346 19966 13358 20018
rect 13410 19966 13422 20018
rect 13794 19966 13806 20018
rect 13858 19966 13870 20018
rect 17938 19966 17950 20018
rect 18002 19966 18014 20018
rect 29138 19966 29150 20018
rect 29202 19966 29214 20018
rect 33282 19966 33294 20018
rect 33346 19966 33358 20018
rect 33730 19966 33742 20018
rect 33794 19966 33806 20018
rect 34290 19966 34302 20018
rect 34354 19966 34366 20018
rect 17278 19954 17330 19966
rect 29486 19954 29538 19966
rect 8766 19906 8818 19918
rect 22094 19906 22146 19918
rect 8306 19854 8318 19906
rect 8370 19854 8382 19906
rect 12002 19854 12014 19906
rect 12066 19854 12078 19906
rect 23202 19854 23214 19906
rect 23266 19854 23278 19906
rect 30930 19854 30942 19906
rect 30994 19854 31006 19906
rect 33058 19854 33070 19906
rect 33122 19854 33134 19906
rect 8766 19842 8818 19854
rect 22094 19842 22146 19854
rect 7758 19794 7810 19806
rect 7758 19730 7810 19742
rect 16942 19794 16994 19806
rect 16942 19730 16994 19742
rect 20974 19794 21026 19806
rect 20974 19730 21026 19742
rect 26014 19794 26066 19806
rect 26014 19730 26066 19742
rect 37326 19794 37378 19806
rect 37326 19730 37378 19742
rect 1344 19626 38640 19660
rect 1344 19574 5876 19626
rect 5928 19574 5980 19626
rect 6032 19574 6084 19626
rect 6136 19574 15200 19626
rect 15252 19574 15304 19626
rect 15356 19574 15408 19626
rect 15460 19574 24524 19626
rect 24576 19574 24628 19626
rect 24680 19574 24732 19626
rect 24784 19574 33848 19626
rect 33900 19574 33952 19626
rect 34004 19574 34056 19626
rect 34108 19574 38640 19626
rect 1344 19540 38640 19574
rect 13358 19458 13410 19470
rect 13358 19394 13410 19406
rect 17726 19346 17778 19358
rect 37326 19346 37378 19358
rect 4050 19294 4062 19346
rect 4114 19294 4126 19346
rect 12450 19294 12462 19346
rect 12514 19294 12526 19346
rect 19506 19294 19518 19346
rect 19570 19294 19582 19346
rect 36978 19294 36990 19346
rect 37042 19294 37054 19346
rect 17726 19282 17778 19294
rect 37326 19282 37378 19294
rect 37662 19346 37714 19358
rect 37662 19282 37714 19294
rect 10446 19234 10498 19246
rect 17054 19234 17106 19246
rect 28590 19234 28642 19246
rect 5842 19182 5854 19234
rect 5906 19182 5918 19234
rect 9986 19182 9998 19234
rect 10050 19182 10062 19234
rect 12674 19182 12686 19234
rect 12738 19182 12750 19234
rect 16370 19182 16382 19234
rect 16434 19182 16446 19234
rect 22082 19182 22094 19234
rect 22146 19182 22158 19234
rect 27906 19182 27918 19234
rect 27970 19182 27982 19234
rect 10446 19170 10498 19182
rect 17054 19170 17106 19182
rect 28590 19170 28642 19182
rect 29262 19234 29314 19246
rect 29698 19182 29710 19234
rect 29762 19182 29774 19234
rect 32946 19182 32958 19234
rect 33010 19182 33022 19234
rect 33506 19182 33518 19234
rect 33570 19182 33582 19234
rect 29262 19170 29314 19182
rect 11118 19122 11170 19134
rect 11790 19122 11842 19134
rect 35758 19122 35810 19134
rect 3042 19070 3054 19122
rect 3106 19070 3118 19122
rect 11442 19070 11454 19122
rect 11506 19070 11518 19122
rect 12114 19070 12126 19122
rect 12178 19070 12190 19122
rect 17378 19070 17390 19122
rect 17442 19070 17454 19122
rect 20626 19070 20638 19122
rect 20690 19070 20702 19122
rect 23762 19070 23774 19122
rect 23826 19070 23838 19122
rect 11118 19058 11170 19070
rect 11790 19058 11842 19070
rect 35758 19058 35810 19070
rect 5854 19010 5906 19022
rect 5854 18946 5906 18958
rect 6974 19010 7026 19022
rect 27582 19010 27634 19022
rect 32734 19010 32786 19022
rect 7746 18958 7758 19010
rect 7810 18958 7822 19010
rect 14130 18958 14142 19010
rect 14194 18958 14206 19010
rect 32162 18958 32174 19010
rect 32226 18958 32238 19010
rect 6974 18946 7026 18958
rect 27582 18946 27634 18958
rect 32734 18946 32786 18958
rect 36542 19010 36594 19022
rect 36542 18946 36594 18958
rect 37774 19010 37826 19022
rect 37774 18946 37826 18958
rect 1344 18842 38800 18876
rect 1344 18790 10538 18842
rect 10590 18790 10642 18842
rect 10694 18790 10746 18842
rect 10798 18790 19862 18842
rect 19914 18790 19966 18842
rect 20018 18790 20070 18842
rect 20122 18790 29186 18842
rect 29238 18790 29290 18842
rect 29342 18790 29394 18842
rect 29446 18790 38510 18842
rect 38562 18790 38614 18842
rect 38666 18790 38718 18842
rect 38770 18790 38800 18842
rect 1344 18756 38800 18790
rect 30382 18674 30434 18686
rect 8306 18622 8318 18674
rect 8370 18622 8382 18674
rect 12338 18622 12350 18674
rect 12402 18622 12414 18674
rect 36082 18622 36094 18674
rect 36146 18622 36158 18674
rect 30382 18610 30434 18622
rect 11006 18562 11058 18574
rect 3042 18510 3054 18562
rect 3106 18510 3118 18562
rect 11006 18498 11058 18510
rect 21870 18562 21922 18574
rect 21870 18498 21922 18510
rect 29150 18562 29202 18574
rect 37214 18562 37266 18574
rect 30706 18510 30718 18562
rect 30770 18510 30782 18562
rect 29150 18498 29202 18510
rect 37214 18498 37266 18510
rect 37550 18562 37602 18574
rect 37550 18498 37602 18510
rect 5294 18450 5346 18462
rect 15486 18450 15538 18462
rect 5842 18398 5854 18450
rect 5906 18398 5918 18450
rect 14914 18398 14926 18450
rect 14978 18398 14990 18450
rect 5294 18386 5346 18398
rect 15486 18386 15538 18398
rect 18958 18450 19010 18462
rect 32958 18450 33010 18462
rect 19506 18398 19518 18450
rect 19570 18398 19582 18450
rect 26338 18398 26350 18450
rect 26402 18398 26414 18450
rect 26898 18398 26910 18450
rect 26962 18398 26974 18450
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 36866 18398 36878 18450
rect 36930 18398 36942 18450
rect 18958 18386 19010 18398
rect 32958 18386 33010 18398
rect 8990 18338 9042 18350
rect 4050 18286 4062 18338
rect 4114 18286 4126 18338
rect 8990 18274 9042 18286
rect 9774 18338 9826 18350
rect 10334 18338 10386 18350
rect 11566 18338 11618 18350
rect 10098 18286 10110 18338
rect 10162 18286 10174 18338
rect 10770 18286 10782 18338
rect 10834 18286 10846 18338
rect 9774 18274 9826 18286
rect 10334 18274 10386 18286
rect 11566 18274 11618 18286
rect 15710 18338 15762 18350
rect 17614 18338 17666 18350
rect 16034 18286 16046 18338
rect 16098 18286 16110 18338
rect 15710 18274 15762 18286
rect 17614 18274 17666 18286
rect 18062 18338 18114 18350
rect 23214 18338 23266 18350
rect 23886 18338 23938 18350
rect 22866 18286 22878 18338
rect 22930 18286 22942 18338
rect 23538 18286 23550 18338
rect 23602 18286 23614 18338
rect 18062 18274 18114 18286
rect 23214 18274 23266 18286
rect 23886 18274 23938 18286
rect 31726 18338 31778 18350
rect 37874 18286 37886 18338
rect 37938 18286 37950 18338
rect 31726 18274 31778 18286
rect 11790 18226 11842 18238
rect 11790 18162 11842 18174
rect 22654 18226 22706 18238
rect 22654 18162 22706 18174
rect 29934 18226 29986 18238
rect 29934 18162 29986 18174
rect 36654 18226 36706 18238
rect 36654 18162 36706 18174
rect 1344 18058 38640 18092
rect 1344 18006 5876 18058
rect 5928 18006 5980 18058
rect 6032 18006 6084 18058
rect 6136 18006 15200 18058
rect 15252 18006 15304 18058
rect 15356 18006 15408 18058
rect 15460 18006 24524 18058
rect 24576 18006 24628 18058
rect 24680 18006 24732 18058
rect 24784 18006 33848 18058
rect 33900 18006 33952 18058
rect 34004 18006 34056 18058
rect 34108 18006 38640 18058
rect 1344 17972 38640 18006
rect 3938 17726 3950 17778
rect 4002 17726 4014 17778
rect 21746 17726 21758 17778
rect 21810 17726 21822 17778
rect 27346 17726 27358 17778
rect 27410 17726 27422 17778
rect 37538 17726 37550 17778
rect 37602 17726 37614 17778
rect 9326 17666 9378 17678
rect 13582 17666 13634 17678
rect 20638 17666 20690 17678
rect 8642 17614 8654 17666
rect 8706 17614 8718 17666
rect 9090 17614 9102 17666
rect 9154 17614 9166 17666
rect 9874 17614 9886 17666
rect 9938 17614 9950 17666
rect 13906 17614 13918 17666
rect 13970 17614 13982 17666
rect 20178 17614 20190 17666
rect 20242 17614 20254 17666
rect 9326 17602 9378 17614
rect 13582 17602 13634 17614
rect 20638 17602 20690 17614
rect 22206 17666 22258 17678
rect 32734 17666 32786 17678
rect 22866 17614 22878 17666
rect 22930 17614 22942 17666
rect 32162 17614 32174 17666
rect 32226 17614 32238 17666
rect 22206 17602 22258 17614
rect 32734 17602 32786 17614
rect 32846 17666 32898 17678
rect 33506 17614 33518 17666
rect 33570 17614 33582 17666
rect 38210 17614 38222 17666
rect 38274 17614 38286 17666
rect 32846 17602 32898 17614
rect 5518 17554 5570 17566
rect 3042 17502 3054 17554
rect 3106 17502 3118 17554
rect 5518 17490 5570 17502
rect 16270 17554 16322 17566
rect 16270 17490 16322 17502
rect 17950 17554 18002 17566
rect 17950 17490 18002 17502
rect 21982 17554 22034 17566
rect 26226 17502 26238 17554
rect 26290 17502 26302 17554
rect 21982 17490 22034 17502
rect 1822 17442 1874 17454
rect 13022 17442 13074 17454
rect 6178 17390 6190 17442
rect 6242 17390 6254 17442
rect 12450 17390 12462 17442
rect 12514 17390 12526 17442
rect 1822 17378 1874 17390
rect 13022 17378 13074 17390
rect 17054 17442 17106 17454
rect 17054 17378 17106 17390
rect 17166 17442 17218 17454
rect 25902 17442 25954 17454
rect 25218 17390 25230 17442
rect 25282 17390 25294 17442
rect 17166 17378 17218 17390
rect 25902 17378 25954 17390
rect 29038 17442 29090 17454
rect 36542 17442 36594 17454
rect 29810 17390 29822 17442
rect 29874 17390 29886 17442
rect 35970 17390 35982 17442
rect 36034 17390 36046 17442
rect 29038 17378 29090 17390
rect 36542 17378 36594 17390
rect 1344 17274 38800 17308
rect 1344 17222 10538 17274
rect 10590 17222 10642 17274
rect 10694 17222 10746 17274
rect 10798 17222 19862 17274
rect 19914 17222 19966 17274
rect 20018 17222 20070 17274
rect 20122 17222 29186 17274
rect 29238 17222 29290 17274
rect 29342 17222 29394 17274
rect 29446 17222 38510 17274
rect 38562 17222 38614 17274
rect 38666 17222 38718 17274
rect 38770 17222 38800 17274
rect 1344 17188 38800 17222
rect 8990 17106 9042 17118
rect 15262 17106 15314 17118
rect 4946 17054 4958 17106
rect 5010 17054 5022 17106
rect 14018 17054 14030 17106
rect 14082 17054 14094 17106
rect 23538 17054 23550 17106
rect 23602 17054 23614 17106
rect 37202 17054 37214 17106
rect 37266 17054 37278 17106
rect 8990 17042 9042 17054
rect 15262 17042 15314 17054
rect 24110 16994 24162 17006
rect 6178 16942 6190 16994
rect 6242 16942 6254 16994
rect 6962 16942 6974 16994
rect 7026 16942 7038 16994
rect 10770 16942 10782 16994
rect 10834 16942 10846 16994
rect 17826 16942 17838 16994
rect 17890 16942 17902 16994
rect 24110 16930 24162 16942
rect 24670 16994 24722 17006
rect 25566 16994 25618 17006
rect 25218 16942 25230 16994
rect 25282 16942 25294 16994
rect 24670 16930 24722 16942
rect 25566 16930 25618 16942
rect 28926 16994 28978 17006
rect 31938 16942 31950 16994
rect 32002 16942 32014 16994
rect 33058 16942 33070 16994
rect 33122 16942 33134 16994
rect 28926 16930 28978 16942
rect 2158 16882 2210 16894
rect 11342 16882 11394 16894
rect 20638 16882 20690 16894
rect 26014 16882 26066 16894
rect 34302 16882 34354 16894
rect 2594 16830 2606 16882
rect 2658 16830 2670 16882
rect 5954 16830 5966 16882
rect 6018 16830 6030 16882
rect 9986 16830 9998 16882
rect 10050 16830 10062 16882
rect 11778 16830 11790 16882
rect 11842 16830 11854 16882
rect 16706 16830 16718 16882
rect 16770 16830 16782 16882
rect 21074 16830 21086 16882
rect 21138 16830 21150 16882
rect 26562 16830 26574 16882
rect 26626 16830 26638 16882
rect 33282 16830 33294 16882
rect 33346 16830 33358 16882
rect 34738 16830 34750 16882
rect 34802 16830 34814 16882
rect 2158 16818 2210 16830
rect 11342 16818 11394 16830
rect 20638 16818 20690 16830
rect 26014 16818 26066 16830
rect 34302 16818 34354 16830
rect 8542 16770 8594 16782
rect 30606 16770 30658 16782
rect 7970 16718 7982 16770
rect 8034 16718 8046 16770
rect 16034 16718 16046 16770
rect 16098 16718 16110 16770
rect 19170 16718 19182 16770
rect 19234 16718 19246 16770
rect 24322 16718 24334 16770
rect 24386 16718 24398 16770
rect 30930 16718 30942 16770
rect 30994 16718 31006 16770
rect 8542 16706 8594 16718
rect 30606 16706 30658 16718
rect 5630 16658 5682 16670
rect 5630 16594 5682 16606
rect 14814 16658 14866 16670
rect 14814 16594 14866 16606
rect 29710 16658 29762 16670
rect 29710 16594 29762 16606
rect 37774 16658 37826 16670
rect 37774 16594 37826 16606
rect 1344 16490 38640 16524
rect 1344 16438 5876 16490
rect 5928 16438 5980 16490
rect 6032 16438 6084 16490
rect 6136 16438 15200 16490
rect 15252 16438 15304 16490
rect 15356 16438 15408 16490
rect 15460 16438 24524 16490
rect 24576 16438 24628 16490
rect 24680 16438 24732 16490
rect 24784 16438 33848 16490
rect 33900 16438 33952 16490
rect 34004 16438 34056 16490
rect 34108 16438 38640 16490
rect 1344 16404 38640 16438
rect 23438 16322 23490 16334
rect 23438 16258 23490 16270
rect 7534 16210 7586 16222
rect 21982 16210 22034 16222
rect 4050 16158 4062 16210
rect 4114 16158 4126 16210
rect 15922 16158 15934 16210
rect 15986 16158 15998 16210
rect 21634 16158 21646 16210
rect 21698 16158 21710 16210
rect 7534 16146 7586 16158
rect 21982 16146 22034 16158
rect 27582 16210 27634 16222
rect 28466 16158 28478 16210
rect 28530 16158 28542 16210
rect 30146 16158 30158 16210
rect 30210 16158 30222 16210
rect 27582 16146 27634 16158
rect 7758 16098 7810 16110
rect 14142 16098 14194 16110
rect 5842 16046 5854 16098
rect 5906 16046 5918 16098
rect 8306 16046 8318 16098
rect 8370 16046 8382 16098
rect 12786 16046 12798 16098
rect 12850 16046 12862 16098
rect 7758 16034 7810 16046
rect 14142 16034 14194 16046
rect 16382 16098 16434 16110
rect 26910 16098 26962 16110
rect 16706 16046 16718 16098
rect 16770 16046 16782 16098
rect 26562 16046 26574 16098
rect 26626 16046 26638 16098
rect 28354 16046 28366 16098
rect 28418 16046 28430 16098
rect 30818 16046 30830 16098
rect 30882 16046 30894 16098
rect 31266 16046 31278 16098
rect 31330 16046 31342 16098
rect 37202 16046 37214 16098
rect 37266 16046 37278 16098
rect 16382 16034 16434 16046
rect 26910 16034 26962 16046
rect 1710 15986 1762 15998
rect 20414 15986 20466 15998
rect 37662 15986 37714 15998
rect 3042 15934 3054 15986
rect 3106 15934 3118 15986
rect 5618 15934 5630 15986
rect 5682 15934 5694 15986
rect 12114 15934 12126 15986
rect 12178 15934 12190 15986
rect 14690 15934 14702 15986
rect 14754 15934 14766 15986
rect 20066 15934 20078 15986
rect 20130 15934 20142 15986
rect 34626 15934 34638 15986
rect 34690 15934 34702 15986
rect 36978 15934 36990 15986
rect 37042 15934 37054 15986
rect 1710 15922 1762 15934
rect 20414 15922 20466 15934
rect 37662 15922 37714 15934
rect 2046 15874 2098 15886
rect 2046 15810 2098 15822
rect 5070 15874 5122 15886
rect 5070 15810 5122 15822
rect 6414 15874 6466 15886
rect 6414 15810 6466 15822
rect 7422 15874 7474 15886
rect 11454 15874 11506 15886
rect 10882 15822 10894 15874
rect 10946 15822 10958 15874
rect 7422 15810 7474 15822
rect 11454 15810 11506 15822
rect 13582 15874 13634 15886
rect 19854 15874 19906 15886
rect 27694 15874 27746 15886
rect 19282 15822 19294 15874
rect 19346 15822 19358 15874
rect 24210 15822 24222 15874
rect 24274 15822 24286 15874
rect 13582 15810 13634 15822
rect 19854 15810 19906 15822
rect 27694 15810 27746 15822
rect 37774 15874 37826 15886
rect 37774 15810 37826 15822
rect 1344 15706 38800 15740
rect 1344 15654 10538 15706
rect 10590 15654 10642 15706
rect 10694 15654 10746 15706
rect 10798 15654 19862 15706
rect 19914 15654 19966 15706
rect 20018 15654 20070 15706
rect 20122 15654 29186 15706
rect 29238 15654 29290 15706
rect 29342 15654 29394 15706
rect 29446 15654 38510 15706
rect 38562 15654 38614 15706
rect 38666 15654 38718 15706
rect 38770 15654 38800 15706
rect 1344 15620 38800 15654
rect 16718 15538 16770 15550
rect 22766 15538 22818 15550
rect 2370 15486 2382 15538
rect 2434 15486 2446 15538
rect 5954 15486 5966 15538
rect 6018 15486 6030 15538
rect 18946 15486 18958 15538
rect 19010 15486 19022 15538
rect 33730 15486 33742 15538
rect 33794 15486 33806 15538
rect 16718 15474 16770 15486
rect 22766 15474 22818 15486
rect 12786 15374 12798 15426
rect 12850 15374 12862 15426
rect 24098 15374 24110 15426
rect 24162 15374 24174 15426
rect 5294 15314 5346 15326
rect 9102 15314 9154 15326
rect 21646 15314 21698 15326
rect 36430 15314 36482 15326
rect 4610 15262 4622 15314
rect 4674 15262 4686 15314
rect 8530 15262 8542 15314
rect 8594 15262 8606 15314
rect 14802 15262 14814 15314
rect 14866 15262 14878 15314
rect 15362 15262 15374 15314
rect 15426 15262 15438 15314
rect 16034 15262 16046 15314
rect 16098 15262 16110 15314
rect 21298 15262 21310 15314
rect 21362 15262 21374 15314
rect 29362 15262 29374 15314
rect 29426 15262 29438 15314
rect 31490 15262 31502 15314
rect 31554 15262 31566 15314
rect 35970 15262 35982 15314
rect 36034 15262 36046 15314
rect 5294 15250 5346 15262
rect 9102 15250 9154 15262
rect 21646 15250 21698 15262
rect 36430 15250 36482 15262
rect 17838 15202 17890 15214
rect 32958 15202 33010 15214
rect 15138 15150 15150 15202
rect 15202 15150 15214 15202
rect 16258 15150 16270 15202
rect 16322 15150 16334 15202
rect 17490 15150 17502 15202
rect 17554 15150 17566 15202
rect 23090 15150 23102 15202
rect 23154 15150 23166 15202
rect 25778 15150 25790 15202
rect 25842 15150 25854 15202
rect 17838 15138 17890 15150
rect 32958 15138 33010 15150
rect 1598 15090 1650 15102
rect 1598 15026 1650 15038
rect 5406 15090 5458 15102
rect 5406 15026 5458 15038
rect 18174 15090 18226 15102
rect 18174 15026 18226 15038
rect 32286 15090 32338 15102
rect 32286 15026 32338 15038
rect 1344 14922 38640 14956
rect 1344 14870 5876 14922
rect 5928 14870 5980 14922
rect 6032 14870 6084 14922
rect 6136 14870 15200 14922
rect 15252 14870 15304 14922
rect 15356 14870 15408 14922
rect 15460 14870 24524 14922
rect 24576 14870 24628 14922
rect 24680 14870 24732 14922
rect 24784 14870 33848 14922
rect 33900 14870 33952 14922
rect 34004 14870 34056 14922
rect 34108 14870 38640 14922
rect 1344 14836 38640 14870
rect 19518 14642 19570 14654
rect 3602 14590 3614 14642
rect 3666 14590 3678 14642
rect 5842 14590 5854 14642
rect 5906 14590 5918 14642
rect 8082 14590 8094 14642
rect 8146 14590 8158 14642
rect 16818 14590 16830 14642
rect 16882 14590 16894 14642
rect 19518 14578 19570 14590
rect 19966 14642 20018 14654
rect 28466 14590 28478 14642
rect 28530 14590 28542 14642
rect 19966 14578 20018 14590
rect 27134 14530 27186 14542
rect 29038 14530 29090 14542
rect 32846 14530 32898 14542
rect 12338 14478 12350 14530
rect 12402 14478 12414 14530
rect 12898 14478 12910 14530
rect 12962 14478 12974 14530
rect 13794 14478 13806 14530
rect 13858 14478 13870 14530
rect 26786 14478 26798 14530
rect 26850 14478 26862 14530
rect 28354 14478 28366 14530
rect 28418 14478 28430 14530
rect 29698 14478 29710 14530
rect 29762 14478 29774 14530
rect 33394 14478 33406 14530
rect 33458 14478 33470 14530
rect 37202 14478 37214 14530
rect 37266 14478 37278 14530
rect 27134 14466 27186 14478
rect 29038 14466 29090 14478
rect 32846 14466 32898 14478
rect 1934 14418 1986 14430
rect 5630 14418 5682 14430
rect 10110 14418 10162 14430
rect 4946 14366 4958 14418
rect 5010 14366 5022 14418
rect 7074 14366 7086 14418
rect 7138 14366 7150 14418
rect 1934 14354 1986 14366
rect 5630 14354 5682 14366
rect 10110 14354 10162 14366
rect 27582 14418 27634 14430
rect 27906 14366 27918 14418
rect 27970 14366 27982 14418
rect 36978 14366 36990 14418
rect 37042 14366 37054 14418
rect 27582 14354 27634 14366
rect 2046 14306 2098 14318
rect 2046 14242 2098 14254
rect 8654 14306 8706 14318
rect 8654 14242 8706 14254
rect 9102 14306 9154 14318
rect 9102 14242 9154 14254
rect 9326 14306 9378 14318
rect 9326 14242 9378 14254
rect 23662 14306 23714 14318
rect 32734 14306 32786 14318
rect 36542 14306 36594 14318
rect 24322 14254 24334 14306
rect 24386 14254 24398 14306
rect 32162 14254 32174 14306
rect 32226 14254 32238 14306
rect 35970 14254 35982 14306
rect 36034 14254 36046 14306
rect 23662 14242 23714 14254
rect 32734 14242 32786 14254
rect 36542 14242 36594 14254
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 38334 13970 38386 13982
rect 4722 13918 4734 13970
rect 4786 13918 4798 13970
rect 8306 13918 8318 13970
rect 8370 13918 8382 13970
rect 16370 13918 16382 13970
rect 16434 13918 16446 13970
rect 20402 13918 20414 13970
rect 20466 13918 20478 13970
rect 24210 13918 24222 13970
rect 24274 13918 24286 13970
rect 28018 13918 28030 13970
rect 28082 13918 28094 13970
rect 37762 13918 37774 13970
rect 37826 13918 37838 13970
rect 38334 13906 38386 13918
rect 12350 13858 12402 13870
rect 12350 13794 12402 13806
rect 31838 13858 31890 13870
rect 33058 13806 33070 13858
rect 33122 13806 33134 13858
rect 33730 13806 33742 13858
rect 33794 13806 33806 13858
rect 31838 13794 31890 13806
rect 1822 13746 1874 13758
rect 5630 13746 5682 13758
rect 9438 13746 9490 13758
rect 17278 13746 17330 13758
rect 21086 13746 21138 13758
rect 34638 13746 34690 13758
rect 2258 13694 2270 13746
rect 2322 13694 2334 13746
rect 6066 13694 6078 13746
rect 6130 13694 6142 13746
rect 10098 13694 10110 13746
rect 10162 13694 10174 13746
rect 13346 13694 13358 13746
rect 13410 13694 13422 13746
rect 13906 13694 13918 13746
rect 13970 13694 13982 13746
rect 17938 13694 17950 13746
rect 18002 13694 18014 13746
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 25218 13694 25230 13746
rect 25282 13694 25294 13746
rect 25666 13694 25678 13746
rect 25730 13694 25742 13746
rect 29026 13694 29038 13746
rect 29090 13694 29102 13746
rect 29586 13694 29598 13746
rect 29650 13694 29662 13746
rect 33282 13694 33294 13746
rect 33346 13694 33358 13746
rect 33954 13694 33966 13746
rect 34018 13694 34030 13746
rect 35186 13694 35198 13746
rect 35250 13694 35262 13746
rect 1822 13682 1874 13694
rect 5630 13682 5682 13694
rect 9438 13682 9490 13694
rect 17278 13682 17330 13694
rect 21086 13682 21138 13694
rect 34638 13682 34690 13694
rect 5294 13522 5346 13534
rect 5294 13458 5346 13470
rect 9102 13522 9154 13534
rect 9102 13458 9154 13470
rect 13134 13522 13186 13534
rect 13134 13458 13186 13470
rect 16942 13522 16994 13534
rect 16942 13458 16994 13470
rect 20974 13522 21026 13534
rect 20974 13458 21026 13470
rect 24782 13522 24834 13534
rect 24782 13458 24834 13470
rect 28814 13522 28866 13534
rect 28814 13458 28866 13470
rect 32622 13522 32674 13534
rect 32622 13458 32674 13470
rect 1344 13354 38640 13388
rect 1344 13302 5876 13354
rect 5928 13302 5980 13354
rect 6032 13302 6084 13354
rect 6136 13302 15200 13354
rect 15252 13302 15304 13354
rect 15356 13302 15408 13354
rect 15460 13302 24524 13354
rect 24576 13302 24628 13354
rect 24680 13302 24732 13354
rect 24784 13302 33848 13354
rect 33900 13302 33952 13354
rect 34004 13302 34056 13354
rect 34108 13302 38640 13354
rect 1344 13268 38640 13302
rect 1934 13074 1986 13086
rect 13022 13074 13074 13086
rect 37662 13074 37714 13086
rect 3826 13022 3838 13074
rect 3890 13022 3902 13074
rect 12450 13022 12462 13074
rect 12514 13022 12526 13074
rect 22194 13022 22206 13074
rect 22258 13022 22270 13074
rect 34514 13022 34526 13074
rect 34578 13022 34590 13074
rect 1934 13010 1986 13022
rect 13022 13010 13074 13022
rect 37662 13010 37714 13022
rect 7646 12962 7698 12974
rect 20862 12962 20914 12974
rect 23214 12962 23266 12974
rect 33070 12962 33122 12974
rect 5954 12910 5966 12962
rect 6018 12910 6030 12962
rect 8194 12910 8206 12962
rect 8258 12910 8270 12962
rect 13458 12910 13470 12962
rect 13522 12910 13534 12962
rect 13906 12910 13918 12962
rect 13970 12910 13982 12962
rect 20178 12910 20190 12962
rect 20242 12910 20254 12962
rect 22418 12910 22430 12962
rect 22482 12910 22494 12962
rect 23874 12910 23886 12962
rect 23938 12910 23950 12962
rect 32610 12910 32622 12962
rect 32674 12910 32686 12962
rect 37202 12910 37214 12962
rect 37266 12910 37278 12962
rect 7646 12898 7698 12910
rect 20862 12898 20914 12910
rect 23214 12898 23266 12910
rect 33070 12898 33122 12910
rect 6862 12850 6914 12862
rect 2258 12798 2270 12850
rect 2322 12798 2334 12850
rect 4946 12798 4958 12850
rect 5010 12798 5022 12850
rect 6178 12798 6190 12850
rect 6242 12798 6254 12850
rect 6514 12798 6526 12850
rect 6578 12798 6590 12850
rect 6862 12786 6914 12798
rect 12126 12850 12178 12862
rect 12126 12786 12178 12798
rect 16270 12850 16322 12862
rect 16270 12786 16322 12798
rect 17950 12850 18002 12862
rect 17950 12786 18002 12798
rect 21534 12850 21586 12862
rect 21858 12798 21870 12850
rect 21922 12798 21934 12850
rect 35522 12798 35534 12850
rect 35586 12798 35598 12850
rect 21534 12786 21586 12798
rect 7310 12738 7362 12750
rect 11342 12738 11394 12750
rect 10546 12686 10558 12738
rect 10610 12686 10622 12738
rect 7310 12674 7362 12686
rect 11342 12674 11394 12686
rect 11678 12738 11730 12750
rect 11678 12674 11730 12686
rect 17054 12738 17106 12750
rect 17054 12674 17106 12686
rect 17166 12738 17218 12750
rect 26910 12738 26962 12750
rect 26114 12686 26126 12738
rect 26178 12686 26190 12738
rect 17166 12674 17218 12686
rect 26910 12674 26962 12686
rect 29598 12738 29650 12750
rect 37214 12738 37266 12750
rect 30370 12686 30382 12738
rect 30434 12686 30446 12738
rect 29598 12674 29650 12686
rect 37214 12674 37266 12686
rect 37774 12738 37826 12750
rect 37774 12674 37826 12686
rect 1344 12570 38800 12604
rect 1344 12518 10538 12570
rect 10590 12518 10642 12570
rect 10694 12518 10746 12570
rect 10798 12518 19862 12570
rect 19914 12518 19966 12570
rect 20018 12518 20070 12570
rect 20122 12518 29186 12570
rect 29238 12518 29290 12570
rect 29342 12518 29394 12570
rect 29446 12518 38510 12570
rect 38562 12518 38614 12570
rect 38666 12518 38718 12570
rect 38770 12518 38800 12570
rect 1344 12484 38800 12518
rect 37886 12402 37938 12414
rect 4498 12350 4510 12402
rect 4562 12350 4574 12402
rect 16370 12350 16382 12402
rect 16434 12350 16446 12402
rect 22194 12350 22206 12402
rect 22258 12350 22270 12402
rect 36978 12350 36990 12402
rect 37042 12350 37054 12402
rect 37886 12338 37938 12350
rect 8318 12290 8370 12302
rect 24558 12290 24610 12302
rect 33630 12290 33682 12302
rect 12786 12238 12798 12290
rect 12850 12238 12862 12290
rect 17714 12238 17726 12290
rect 17778 12238 17790 12290
rect 24210 12238 24222 12290
rect 24274 12238 24286 12290
rect 26002 12238 26014 12290
rect 26066 12238 26078 12290
rect 28578 12238 28590 12290
rect 28642 12238 28654 12290
rect 31714 12238 31726 12290
rect 31778 12238 31790 12290
rect 33282 12238 33294 12290
rect 33346 12238 33358 12290
rect 8318 12226 8370 12238
rect 24558 12226 24610 12238
rect 33630 12226 33682 12238
rect 37774 12290 37826 12302
rect 37774 12226 37826 12238
rect 1822 12178 1874 12190
rect 5630 12178 5682 12190
rect 13470 12178 13522 12190
rect 19294 12178 19346 12190
rect 33854 12178 33906 12190
rect 2146 12126 2158 12178
rect 2210 12126 2222 12178
rect 5954 12126 5966 12178
rect 6018 12126 6030 12178
rect 13906 12126 13918 12178
rect 13970 12126 13982 12178
rect 17938 12126 17950 12178
rect 18002 12126 18014 12178
rect 19954 12126 19966 12178
rect 20018 12126 20030 12178
rect 23314 12126 23326 12178
rect 23378 12126 23390 12178
rect 34514 12126 34526 12178
rect 34578 12126 34590 12178
rect 1822 12114 1874 12126
rect 5630 12114 5682 12126
rect 13470 12114 13522 12126
rect 19294 12114 19346 12126
rect 33854 12114 33906 12126
rect 9886 12066 9938 12078
rect 10670 12066 10722 12078
rect 10098 12014 10110 12066
rect 10162 12014 10174 12066
rect 9886 12002 9938 12014
rect 10670 12002 10722 12014
rect 11230 12066 11282 12078
rect 18734 12066 18786 12078
rect 25678 12066 25730 12078
rect 11778 12014 11790 12066
rect 11842 12014 11854 12066
rect 19058 12014 19070 12066
rect 19122 12014 19134 12066
rect 23426 12014 23438 12066
rect 23490 12014 23502 12066
rect 27346 12014 27358 12066
rect 27410 12014 27422 12066
rect 30482 12014 30494 12066
rect 30546 12014 30558 12066
rect 11230 12002 11282 12014
rect 18734 12002 18786 12014
rect 25678 12002 25730 12014
rect 5294 11954 5346 11966
rect 5294 11890 5346 11902
rect 9102 11954 9154 11966
rect 16942 11954 16994 11966
rect 10658 11902 10670 11954
rect 10722 11951 10734 11954
rect 11218 11951 11230 11954
rect 10722 11905 11230 11951
rect 10722 11902 10734 11905
rect 11218 11902 11230 11905
rect 11282 11902 11294 11954
rect 9102 11890 9154 11902
rect 16942 11890 16994 11902
rect 22990 11954 23042 11966
rect 22990 11890 23042 11902
rect 37550 11954 37602 11966
rect 37550 11890 37602 11902
rect 1344 11786 38640 11820
rect 1344 11734 5876 11786
rect 5928 11734 5980 11786
rect 6032 11734 6084 11786
rect 6136 11734 15200 11786
rect 15252 11734 15304 11786
rect 15356 11734 15408 11786
rect 15460 11734 24524 11786
rect 24576 11734 24628 11786
rect 24680 11734 24732 11786
rect 24784 11734 33848 11786
rect 33900 11734 33952 11786
rect 34004 11734 34056 11786
rect 34108 11734 38640 11786
rect 1344 11700 38640 11734
rect 7870 11506 7922 11518
rect 15934 11506 15986 11518
rect 4050 11454 4062 11506
rect 4114 11454 4126 11506
rect 12338 11454 12350 11506
rect 12402 11454 12414 11506
rect 15362 11454 15374 11506
rect 15426 11454 15438 11506
rect 7870 11442 7922 11454
rect 15934 11442 15986 11454
rect 16382 11506 16434 11518
rect 22306 11454 22318 11506
rect 22370 11454 22382 11506
rect 25106 11454 25118 11506
rect 25170 11454 25182 11506
rect 34290 11454 34302 11506
rect 34354 11454 34366 11506
rect 38098 11454 38110 11506
rect 38162 11454 38174 11506
rect 16382 11442 16434 11454
rect 8094 11394 8146 11406
rect 16830 11394 16882 11406
rect 33742 11394 33794 11406
rect 8642 11342 8654 11394
rect 8706 11342 8718 11394
rect 17154 11342 17166 11394
rect 17218 11342 17230 11394
rect 33282 11342 33294 11394
rect 33346 11342 33358 11394
rect 36978 11342 36990 11394
rect 37042 11342 37054 11394
rect 8094 11330 8146 11342
rect 16830 11330 16882 11342
rect 33742 11330 33794 11342
rect 12126 11282 12178 11294
rect 19518 11282 19570 11294
rect 34526 11282 34578 11294
rect 2930 11230 2942 11282
rect 2994 11230 3006 11282
rect 7522 11230 7534 11282
rect 7586 11230 7598 11282
rect 14354 11230 14366 11282
rect 14418 11230 14430 11282
rect 23538 11230 23550 11282
rect 23602 11230 23614 11282
rect 26114 11230 26126 11282
rect 26178 11230 26190 11282
rect 12126 11218 12178 11230
rect 19518 11218 19570 11230
rect 34526 11218 34578 11230
rect 35758 11282 35810 11294
rect 35758 11218 35810 11230
rect 36430 11282 36482 11294
rect 36430 11218 36482 11230
rect 5742 11170 5794 11182
rect 11790 11170 11842 11182
rect 10994 11118 11006 11170
rect 11058 11118 11070 11170
rect 5742 11106 5794 11118
rect 11790 11106 11842 11118
rect 12910 11170 12962 11182
rect 12910 11106 12962 11118
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 20302 11170 20354 11182
rect 20302 11106 20354 11118
rect 20638 11170 20690 11182
rect 20638 11106 20690 11118
rect 30270 11170 30322 11182
rect 35198 11170 35250 11182
rect 31042 11118 31054 11170
rect 31106 11118 31118 11170
rect 30270 11106 30322 11118
rect 35198 11106 35250 11118
rect 35422 11170 35474 11182
rect 35422 11106 35474 11118
rect 36094 11170 36146 11182
rect 36094 11106 36146 11118
rect 1344 11002 38800 11036
rect 1344 10950 10538 11002
rect 10590 10950 10642 11002
rect 10694 10950 10746 11002
rect 10798 10950 19862 11002
rect 19914 10950 19966 11002
rect 20018 10950 20070 11002
rect 20122 10950 29186 11002
rect 29238 10950 29290 11002
rect 29342 10950 29394 11002
rect 29446 10950 38510 11002
rect 38562 10950 38614 11002
rect 38666 10950 38718 11002
rect 38770 10950 38800 11002
rect 1344 10916 38800 10950
rect 8766 10834 8818 10846
rect 5506 10782 5518 10834
rect 5570 10782 5582 10834
rect 8766 10770 8818 10782
rect 9774 10834 9826 10846
rect 9774 10770 9826 10782
rect 12238 10834 12290 10846
rect 12238 10770 12290 10782
rect 18174 10834 18226 10846
rect 38334 10834 38386 10846
rect 35858 10782 35870 10834
rect 35922 10782 35934 10834
rect 18174 10770 18226 10782
rect 38334 10770 38386 10782
rect 4734 10722 4786 10734
rect 2482 10670 2494 10722
rect 2546 10670 2558 10722
rect 4734 10658 4786 10670
rect 9662 10722 9714 10734
rect 13806 10722 13858 10734
rect 10434 10670 10446 10722
rect 10498 10670 10510 10722
rect 17378 10670 17390 10722
rect 17442 10670 17454 10722
rect 20178 10670 20190 10722
rect 20242 10670 20254 10722
rect 22978 10670 22990 10722
rect 23042 10670 23054 10722
rect 27234 10670 27246 10722
rect 27298 10670 27310 10722
rect 30370 10670 30382 10722
rect 30434 10670 30446 10722
rect 9662 10658 9714 10670
rect 13806 10658 13858 10670
rect 8206 10610 8258 10622
rect 16494 10610 16546 10622
rect 33182 10610 33234 10622
rect 36990 10610 37042 10622
rect 7746 10558 7758 10610
rect 7810 10558 7822 10610
rect 16146 10558 16158 10610
rect 16210 10558 16222 10610
rect 17602 10558 17614 10610
rect 17666 10558 17678 10610
rect 33618 10558 33630 10610
rect 33682 10558 33694 10610
rect 8206 10546 8258 10558
rect 16494 10546 16546 10558
rect 33182 10546 33234 10558
rect 36990 10546 37042 10558
rect 3378 10446 3390 10498
rect 3442 10446 3454 10498
rect 11778 10446 11790 10498
rect 11842 10446 11854 10498
rect 19394 10446 19406 10498
rect 19458 10446 19470 10498
rect 21970 10446 21982 10498
rect 22034 10446 22046 10498
rect 26226 10446 26238 10498
rect 26290 10446 26302 10498
rect 29026 10446 29038 10498
rect 29090 10446 29102 10498
rect 37538 10446 37550 10498
rect 37602 10446 37614 10498
rect 13022 10386 13074 10398
rect 13022 10322 13074 10334
rect 36654 10386 36706 10398
rect 36654 10322 36706 10334
rect 1344 10218 38640 10252
rect 1344 10166 5876 10218
rect 5928 10166 5980 10218
rect 6032 10166 6084 10218
rect 6136 10166 15200 10218
rect 15252 10166 15304 10218
rect 15356 10166 15408 10218
rect 15460 10166 24524 10218
rect 24576 10166 24628 10218
rect 24680 10166 24732 10218
rect 24784 10166 33848 10218
rect 33900 10166 33952 10218
rect 34004 10166 34056 10218
rect 34108 10166 38640 10218
rect 1344 10132 38640 10166
rect 37774 10050 37826 10062
rect 37774 9986 37826 9998
rect 15150 9938 15202 9950
rect 17390 9938 17442 9950
rect 3490 9886 3502 9938
rect 3554 9886 3566 9938
rect 9986 9886 9998 9938
rect 10050 9886 10062 9938
rect 11442 9886 11454 9938
rect 11506 9886 11518 9938
rect 16930 9886 16942 9938
rect 16994 9886 17006 9938
rect 15150 9874 15202 9886
rect 17390 9874 17442 9886
rect 17838 9938 17890 9950
rect 19282 9886 19294 9938
rect 19346 9886 19358 9938
rect 22418 9886 22430 9938
rect 22482 9886 22494 9938
rect 27570 9886 27582 9938
rect 27634 9886 27646 9938
rect 30930 9886 30942 9938
rect 30994 9886 31006 9938
rect 33842 9886 33854 9938
rect 33906 9886 33918 9938
rect 17838 9874 17890 9886
rect 8990 9826 9042 9838
rect 8530 9774 8542 9826
rect 8594 9774 8606 9826
rect 9874 9774 9886 9826
rect 9938 9774 9950 9826
rect 35746 9774 35758 9826
rect 35810 9774 35822 9826
rect 8990 9762 9042 9774
rect 6302 9714 6354 9726
rect 2370 9662 2382 9714
rect 2434 9662 2446 9714
rect 12786 9662 12798 9714
rect 12850 9662 12862 9714
rect 14802 9662 14814 9714
rect 14866 9662 14878 9714
rect 15698 9662 15710 9714
rect 15762 9662 15774 9714
rect 20626 9662 20638 9714
rect 20690 9662 20702 9714
rect 23538 9662 23550 9714
rect 23602 9662 23614 9714
rect 26562 9662 26574 9714
rect 26626 9662 26638 9714
rect 31938 9662 31950 9714
rect 32002 9662 32014 9714
rect 34738 9662 34750 9714
rect 34802 9662 34814 9714
rect 6302 9650 6354 9662
rect 5518 9602 5570 9614
rect 5518 9538 5570 9550
rect 32958 9602 33010 9614
rect 32958 9538 33010 9550
rect 35534 9602 35586 9614
rect 35534 9538 35586 9550
rect 36318 9602 36370 9614
rect 36318 9538 36370 9550
rect 36990 9602 37042 9614
rect 36990 9538 37042 9550
rect 1344 9434 38800 9468
rect 1344 9382 10538 9434
rect 10590 9382 10642 9434
rect 10694 9382 10746 9434
rect 10798 9382 19862 9434
rect 19914 9382 19966 9434
rect 20018 9382 20070 9434
rect 20122 9382 29186 9434
rect 29238 9382 29290 9434
rect 29342 9382 29394 9434
rect 29446 9382 38510 9434
rect 38562 9382 38614 9434
rect 38666 9382 38718 9434
rect 38770 9382 38800 9434
rect 1344 9348 38800 9382
rect 9662 9266 9714 9278
rect 33966 9266 34018 9278
rect 6178 9214 6190 9266
rect 6242 9214 6254 9266
rect 14130 9214 14142 9266
rect 14194 9214 14206 9266
rect 37314 9214 37326 9266
rect 37378 9214 37390 9266
rect 9662 9202 9714 9214
rect 33966 9202 34018 9214
rect 31166 9154 31218 9166
rect 19394 9102 19406 9154
rect 19458 9102 19470 9154
rect 29922 9102 29934 9154
rect 29986 9102 29998 9154
rect 31166 9090 31218 9102
rect 31502 9154 31554 9166
rect 31502 9090 31554 9102
rect 31838 9154 31890 9166
rect 31838 9090 31890 9102
rect 32174 9154 32226 9166
rect 32174 9090 32226 9102
rect 33294 9154 33346 9166
rect 33294 9090 33346 9102
rect 33630 9154 33682 9166
rect 33630 9090 33682 9102
rect 3054 9042 3106 9054
rect 11230 9042 11282 9054
rect 15038 9042 15090 9054
rect 34190 9042 34242 9054
rect 3714 8990 3726 9042
rect 3778 8990 3790 9042
rect 11666 8990 11678 9042
rect 11730 8990 11742 9042
rect 30930 8990 30942 9042
rect 30994 8990 31006 9042
rect 32386 8990 32398 9042
rect 32450 8990 32462 9042
rect 34738 8990 34750 9042
rect 34802 8990 34814 9042
rect 3054 8978 3106 8990
rect 11230 8978 11282 8990
rect 15038 8978 15090 8990
rect 34190 8978 34242 8990
rect 7086 8930 7138 8942
rect 18386 8878 18398 8930
rect 18450 8878 18462 8930
rect 28914 8878 28926 8930
rect 28978 8878 28990 8930
rect 7086 8866 7138 8878
rect 6750 8818 6802 8830
rect 6750 8754 6802 8766
rect 14702 8818 14754 8830
rect 14702 8754 14754 8766
rect 37886 8818 37938 8830
rect 37886 8754 37938 8766
rect 1344 8650 38640 8684
rect 1344 8598 5876 8650
rect 5928 8598 5980 8650
rect 6032 8598 6084 8650
rect 6136 8598 15200 8650
rect 15252 8598 15304 8650
rect 15356 8598 15408 8650
rect 15460 8598 24524 8650
rect 24576 8598 24628 8650
rect 24680 8598 24732 8650
rect 24784 8598 33848 8650
rect 33900 8598 33952 8650
rect 34004 8598 34056 8650
rect 34108 8598 38640 8650
rect 1344 8564 38640 8598
rect 31166 8370 31218 8382
rect 3602 8318 3614 8370
rect 3666 8318 3678 8370
rect 7298 8318 7310 8370
rect 7362 8318 7374 8370
rect 11442 8318 11454 8370
rect 11506 8318 11518 8370
rect 15922 8318 15934 8370
rect 15986 8318 15998 8370
rect 18722 8318 18734 8370
rect 18786 8318 18798 8370
rect 27570 8318 27582 8370
rect 27634 8318 27646 8370
rect 31378 8318 31390 8370
rect 31442 8318 31454 8370
rect 34626 8318 34638 8370
rect 34690 8318 34702 8370
rect 37762 8318 37774 8370
rect 37826 8318 37838 8370
rect 31166 8306 31218 8318
rect 21970 8206 21982 8258
rect 22034 8206 22046 8258
rect 29810 8206 29822 8258
rect 29874 8206 29886 8258
rect 4946 8094 4958 8146
rect 5010 8094 5022 8146
rect 6066 8094 6078 8146
rect 6130 8094 6142 8146
rect 12450 8094 12462 8146
rect 12514 8094 12526 8146
rect 17154 8094 17166 8146
rect 17218 8094 17230 8146
rect 19730 8094 19742 8146
rect 19794 8094 19806 8146
rect 26562 8094 26574 8146
rect 26626 8094 26638 8146
rect 32498 8094 32510 8146
rect 32562 8094 32574 8146
rect 35634 8094 35646 8146
rect 35698 8094 35710 8146
rect 22206 8034 22258 8046
rect 22206 7970 22258 7982
rect 30046 8034 30098 8046
rect 30046 7970 30098 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 36990 8034 37042 8046
rect 36990 7970 37042 7982
rect 1344 7866 38800 7900
rect 1344 7814 10538 7866
rect 10590 7814 10642 7866
rect 10694 7814 10746 7866
rect 10798 7814 19862 7866
rect 19914 7814 19966 7866
rect 20018 7814 20070 7866
rect 20122 7814 29186 7866
rect 29238 7814 29290 7866
rect 29342 7814 29394 7866
rect 29446 7814 38510 7866
rect 38562 7814 38614 7866
rect 38666 7814 38718 7866
rect 38770 7814 38800 7866
rect 1344 7780 38800 7814
rect 5630 7698 5682 7710
rect 4722 7646 4734 7698
rect 4786 7646 4798 7698
rect 5630 7634 5682 7646
rect 33406 7698 33458 7710
rect 33406 7634 33458 7646
rect 36654 7586 36706 7598
rect 6850 7534 6862 7586
rect 6914 7534 6926 7586
rect 11890 7534 11902 7586
rect 11954 7534 11966 7586
rect 14354 7534 14366 7586
rect 14418 7534 14430 7586
rect 27682 7534 27694 7586
rect 27746 7534 27758 7586
rect 30482 7534 30494 7586
rect 30546 7534 30558 7586
rect 36082 7534 36094 7586
rect 36146 7534 36158 7586
rect 38098 7534 38110 7586
rect 38162 7534 38174 7586
rect 36654 7522 36706 7534
rect 1822 7474 1874 7486
rect 33070 7474 33122 7486
rect 2258 7422 2270 7474
rect 2322 7422 2334 7474
rect 36978 7422 36990 7474
rect 37042 7422 37054 7474
rect 1822 7410 1874 7422
rect 33070 7410 33122 7422
rect 29262 7362 29314 7374
rect 7858 7310 7870 7362
rect 7922 7310 7934 7362
rect 10546 7310 10558 7362
rect 10610 7310 10622 7362
rect 13346 7310 13358 7362
rect 13410 7310 13422 7362
rect 28690 7310 28702 7362
rect 28754 7310 28766 7362
rect 29262 7298 29314 7310
rect 29822 7362 29874 7374
rect 31490 7310 31502 7362
rect 31554 7310 31566 7362
rect 34962 7310 34974 7362
rect 35026 7310 35038 7362
rect 29822 7298 29874 7310
rect 5294 7250 5346 7262
rect 29138 7198 29150 7250
rect 29202 7247 29214 7250
rect 29810 7247 29822 7250
rect 29202 7201 29822 7247
rect 29202 7198 29214 7201
rect 29810 7198 29822 7201
rect 29874 7198 29886 7250
rect 5294 7186 5346 7198
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 7634 6750 7646 6802
rect 7698 6750 7710 6802
rect 10658 6750 10670 6802
rect 10722 6750 10734 6802
rect 16818 6750 16830 6802
rect 16882 6750 16894 6802
rect 32386 6750 32398 6802
rect 32450 6750 32462 6802
rect 34178 6750 34190 6802
rect 34242 6750 34254 6802
rect 27246 6690 27298 6702
rect 37774 6690 37826 6702
rect 27682 6638 27694 6690
rect 27746 6638 27758 6690
rect 30706 6638 30718 6690
rect 30770 6638 30782 6690
rect 27246 6626 27298 6638
rect 37774 6626 37826 6638
rect 27918 6578 27970 6590
rect 6626 6526 6638 6578
rect 6690 6526 6702 6578
rect 12002 6526 12014 6578
rect 12066 6526 12078 6578
rect 15698 6526 15710 6578
rect 15762 6526 15774 6578
rect 27918 6514 27970 6526
rect 28254 6578 28306 6590
rect 28254 6514 28306 6526
rect 28590 6578 28642 6590
rect 28590 6514 28642 6526
rect 29150 6578 29202 6590
rect 29150 6514 29202 6526
rect 29486 6578 29538 6590
rect 29486 6514 29538 6526
rect 30158 6578 30210 6590
rect 30158 6514 30210 6526
rect 30494 6578 30546 6590
rect 30494 6514 30546 6526
rect 31278 6578 31330 6590
rect 33170 6526 33182 6578
rect 33234 6526 33246 6578
rect 34962 6526 34974 6578
rect 35026 6526 35038 6578
rect 31278 6514 31330 6526
rect 29822 6466 29874 6478
rect 29822 6402 29874 6414
rect 36990 6466 37042 6478
rect 36990 6402 37042 6414
rect 1344 6298 38800 6332
rect 1344 6246 10538 6298
rect 10590 6246 10642 6298
rect 10694 6246 10746 6298
rect 10798 6246 19862 6298
rect 19914 6246 19966 6298
rect 20018 6246 20070 6298
rect 20122 6246 29186 6298
rect 29238 6246 29290 6298
rect 29342 6246 29394 6298
rect 29446 6246 38510 6298
rect 38562 6246 38614 6298
rect 38666 6246 38718 6298
rect 38770 6246 38800 6298
rect 1344 6212 38800 6246
rect 27694 6130 27746 6142
rect 27694 6066 27746 6078
rect 33406 6130 33458 6142
rect 33406 6066 33458 6078
rect 26686 6018 26738 6030
rect 5730 5966 5742 6018
rect 5794 5966 5806 6018
rect 6850 5966 6862 6018
rect 6914 5966 6926 6018
rect 11778 5966 11790 6018
rect 11842 5966 11854 6018
rect 26686 5954 26738 5966
rect 27022 6018 27074 6030
rect 27022 5954 27074 5966
rect 28030 6018 28082 6030
rect 28030 5954 28082 5966
rect 28366 6018 28418 6030
rect 28366 5954 28418 5966
rect 29038 6018 29090 6030
rect 29038 5954 29090 5966
rect 29374 6018 29426 6030
rect 33070 6018 33122 6030
rect 30258 5966 30270 6018
rect 30322 5966 30334 6018
rect 37986 5966 37998 6018
rect 38050 5966 38062 6018
rect 29374 5954 29426 5966
rect 33070 5954 33122 5966
rect 29710 5906 29762 5918
rect 27458 5854 27470 5906
rect 27522 5854 27534 5906
rect 28802 5854 28814 5906
rect 28866 5854 28878 5906
rect 29710 5842 29762 5854
rect 33854 5906 33906 5918
rect 33854 5842 33906 5854
rect 26462 5794 26514 5806
rect 31950 5794 32002 5806
rect 4722 5742 4734 5794
rect 4786 5742 4798 5794
rect 7970 5742 7982 5794
rect 8034 5742 8046 5794
rect 10546 5742 10558 5794
rect 10610 5742 10622 5794
rect 31378 5742 31390 5794
rect 31442 5742 31454 5794
rect 34402 5742 34414 5794
rect 34466 5742 34478 5794
rect 36754 5742 36766 5794
rect 36818 5742 36830 5794
rect 26462 5730 26514 5742
rect 31950 5730 32002 5742
rect 1344 5514 38640 5548
rect 1344 5462 5876 5514
rect 5928 5462 5980 5514
rect 6032 5462 6084 5514
rect 6136 5462 15200 5514
rect 15252 5462 15304 5514
rect 15356 5462 15408 5514
rect 15460 5462 24524 5514
rect 24576 5462 24628 5514
rect 24680 5462 24732 5514
rect 24784 5462 33848 5514
rect 33900 5462 33952 5514
rect 34004 5462 34056 5514
rect 34108 5462 38640 5514
rect 1344 5428 38640 5462
rect 29710 5234 29762 5246
rect 30370 5182 30382 5234
rect 30434 5182 30446 5234
rect 32386 5182 32398 5234
rect 32450 5182 32462 5234
rect 35186 5182 35198 5234
rect 35250 5182 35262 5234
rect 29710 5170 29762 5182
rect 30830 5122 30882 5134
rect 26786 5070 26798 5122
rect 26850 5070 26862 5122
rect 30830 5058 30882 5070
rect 36990 5122 37042 5134
rect 36990 5058 37042 5070
rect 27022 5010 27074 5022
rect 27022 4946 27074 4958
rect 27358 5010 27410 5022
rect 27358 4946 27410 4958
rect 27694 5010 27746 5022
rect 27694 4946 27746 4958
rect 28030 5010 28082 5022
rect 31602 4958 31614 5010
rect 31666 4958 31678 5010
rect 36082 4958 36094 5010
rect 36146 4958 36158 5010
rect 28030 4946 28082 4958
rect 28366 4898 28418 4910
rect 28366 4834 28418 4846
rect 29262 4898 29314 4910
rect 29262 4834 29314 4846
rect 37774 4898 37826 4910
rect 37774 4834 37826 4846
rect 1344 4730 38800 4764
rect 1344 4678 10538 4730
rect 10590 4678 10642 4730
rect 10694 4678 10746 4730
rect 10798 4678 19862 4730
rect 19914 4678 19966 4730
rect 20018 4678 20070 4730
rect 20122 4678 29186 4730
rect 29238 4678 29290 4730
rect 29342 4678 29394 4730
rect 29446 4678 38510 4730
rect 38562 4678 38614 4730
rect 38666 4678 38718 4730
rect 38770 4678 38800 4730
rect 1344 4644 38800 4678
rect 26686 4562 26738 4574
rect 26686 4498 26738 4510
rect 27358 4562 27410 4574
rect 27358 4498 27410 4510
rect 28702 4562 28754 4574
rect 28702 4498 28754 4510
rect 29038 4562 29090 4574
rect 29038 4498 29090 4510
rect 30494 4562 30546 4574
rect 30494 4498 30546 4510
rect 32510 4562 32562 4574
rect 32510 4498 32562 4510
rect 23102 4450 23154 4462
rect 23102 4386 23154 4398
rect 26126 4450 26178 4462
rect 26126 4386 26178 4398
rect 28030 4450 28082 4462
rect 28030 4386 28082 4398
rect 28366 4450 28418 4462
rect 37762 4398 37774 4450
rect 37826 4398 37838 4450
rect 28366 4386 28418 4398
rect 27694 4338 27746 4350
rect 26450 4286 26462 4338
rect 26514 4286 26526 4338
rect 27122 4286 27134 4338
rect 27186 4286 27198 4338
rect 27694 4274 27746 4286
rect 29374 4338 29426 4350
rect 30942 4338 30994 4350
rect 29810 4286 29822 4338
rect 29874 4286 29886 4338
rect 29374 4274 29426 4286
rect 30942 4274 30994 4286
rect 33070 4338 33122 4350
rect 33070 4274 33122 4286
rect 34638 4338 34690 4350
rect 34638 4274 34690 4286
rect 32050 4174 32062 4226
rect 32114 4174 32126 4226
rect 33506 4174 33518 4226
rect 33570 4174 33582 4226
rect 35186 4174 35198 4226
rect 35250 4174 35262 4226
rect 36754 4174 36766 4226
rect 36818 4174 36830 4226
rect 1344 3946 38640 3980
rect 1344 3894 5876 3946
rect 5928 3894 5980 3946
rect 6032 3894 6084 3946
rect 6136 3894 15200 3946
rect 15252 3894 15304 3946
rect 15356 3894 15408 3946
rect 15460 3894 24524 3946
rect 24576 3894 24628 3946
rect 24680 3894 24732 3946
rect 24784 3894 33848 3946
rect 33900 3894 33952 3946
rect 34004 3894 34056 3946
rect 34108 3894 38640 3946
rect 1344 3860 38640 3894
rect 29710 3666 29762 3678
rect 22866 3614 22878 3666
rect 22930 3614 22942 3666
rect 28914 3614 28926 3666
rect 28978 3614 28990 3666
rect 30482 3614 30494 3666
rect 30546 3614 30558 3666
rect 34290 3614 34302 3666
rect 34354 3614 34366 3666
rect 36418 3614 36430 3666
rect 36482 3614 36494 3666
rect 29710 3602 29762 3614
rect 22430 3554 22482 3566
rect 30046 3554 30098 3566
rect 26898 3502 26910 3554
rect 26962 3502 26974 3554
rect 27570 3502 27582 3554
rect 27634 3502 27646 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 22430 3490 22482 3502
rect 30046 3490 30098 3502
rect 32174 3554 32226 3566
rect 32174 3490 32226 3502
rect 35982 3554 36034 3566
rect 35982 3490 36034 3502
rect 37326 3554 37378 3566
rect 37326 3490 37378 3502
rect 21534 3442 21586 3454
rect 21534 3378 21586 3390
rect 21758 3442 21810 3454
rect 21758 3378 21810 3390
rect 22094 3442 22146 3454
rect 22094 3378 22146 3390
rect 26126 3442 26178 3454
rect 26126 3378 26178 3390
rect 27134 3442 27186 3454
rect 27134 3378 27186 3390
rect 27806 3442 27858 3454
rect 27806 3378 27858 3390
rect 32510 3442 32562 3454
rect 37550 3442 37602 3454
rect 33058 3390 33070 3442
rect 33122 3390 33134 3442
rect 32510 3378 32562 3390
rect 37550 3378 37602 3390
rect 37886 3442 37938 3454
rect 37886 3378 37938 3390
rect 24558 3330 24610 3342
rect 24558 3266 24610 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 1344 3162 38800 3196
rect 1344 3110 10538 3162
rect 10590 3110 10642 3162
rect 10694 3110 10746 3162
rect 10798 3110 19862 3162
rect 19914 3110 19966 3162
rect 20018 3110 20070 3162
rect 20122 3110 29186 3162
rect 29238 3110 29290 3162
rect 29342 3110 29394 3162
rect 29446 3110 38510 3162
rect 38562 3110 38614 3162
rect 38666 3110 38718 3162
rect 38770 3110 38800 3162
rect 1344 3076 38800 3110
<< via1 >>
rect 22206 37214 22258 37266
rect 23102 37214 23154 37266
rect 5876 36822 5928 36874
rect 5980 36822 6032 36874
rect 6084 36822 6136 36874
rect 15200 36822 15252 36874
rect 15304 36822 15356 36874
rect 15408 36822 15460 36874
rect 24524 36822 24576 36874
rect 24628 36822 24680 36874
rect 24732 36822 24784 36874
rect 33848 36822 33900 36874
rect 33952 36822 34004 36874
rect 34056 36822 34108 36874
rect 29374 36654 29426 36706
rect 29710 36654 29762 36706
rect 37774 36654 37826 36706
rect 19518 36542 19570 36594
rect 21310 36542 21362 36594
rect 23102 36542 23154 36594
rect 26126 36542 26178 36594
rect 28814 36542 28866 36594
rect 32622 36542 32674 36594
rect 34414 36542 34466 36594
rect 17726 36430 17778 36482
rect 18398 36430 18450 36482
rect 20190 36430 20242 36482
rect 22206 36430 22258 36482
rect 25678 36430 25730 36482
rect 29710 36430 29762 36482
rect 30718 36430 30770 36482
rect 26686 36318 26738 36370
rect 27134 36318 27186 36370
rect 29934 36318 29986 36370
rect 31614 36318 31666 36370
rect 35310 36318 35362 36370
rect 36206 36318 36258 36370
rect 17950 36206 18002 36258
rect 18622 36206 18674 36258
rect 22654 36206 22706 36258
rect 27470 36206 27522 36258
rect 28366 36206 28418 36258
rect 30494 36206 30546 36258
rect 32174 36206 32226 36258
rect 33742 36206 33794 36258
rect 36542 36206 36594 36258
rect 36990 36206 37042 36258
rect 10538 36038 10590 36090
rect 10642 36038 10694 36090
rect 10746 36038 10798 36090
rect 19862 36038 19914 36090
rect 19966 36038 20018 36090
rect 20070 36038 20122 36090
rect 29186 36038 29238 36090
rect 29290 36038 29342 36090
rect 29394 36038 29446 36090
rect 38510 36038 38562 36090
rect 38614 36038 38666 36090
rect 38718 36038 38770 36090
rect 18174 35870 18226 35922
rect 18846 35870 18898 35922
rect 20190 35870 20242 35922
rect 20526 35870 20578 35922
rect 21534 35870 21586 35922
rect 22206 35870 22258 35922
rect 22542 35870 22594 35922
rect 28702 35870 28754 35922
rect 28926 35870 28978 35922
rect 29822 35870 29874 35922
rect 30718 35870 30770 35922
rect 31950 35870 32002 35922
rect 19854 35758 19906 35810
rect 21198 35758 21250 35810
rect 21870 35758 21922 35810
rect 23102 35758 23154 35810
rect 23438 35758 23490 35810
rect 23774 35758 23826 35810
rect 24110 35758 24162 35810
rect 34750 35758 34802 35810
rect 35086 35758 35138 35810
rect 20750 35646 20802 35698
rect 26798 35646 26850 35698
rect 27358 35646 27410 35698
rect 29150 35646 29202 35698
rect 30494 35646 30546 35698
rect 31614 35646 31666 35698
rect 33182 35646 33234 35698
rect 34526 35646 34578 35698
rect 35422 35646 35474 35698
rect 37102 35646 37154 35698
rect 26014 35534 26066 35586
rect 27806 35534 27858 35586
rect 33630 35534 33682 35586
rect 36430 35534 36482 35586
rect 37774 35422 37826 35474
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 35646 35086 35698 35138
rect 20414 34974 20466 35026
rect 22878 34974 22930 35026
rect 23550 34974 23602 35026
rect 24222 34974 24274 35026
rect 37662 34974 37714 35026
rect 24446 34862 24498 34914
rect 25342 34862 25394 34914
rect 26126 34862 26178 34914
rect 32398 34862 32450 34914
rect 36990 34862 37042 34914
rect 24782 34750 24834 34802
rect 25678 34750 25730 34802
rect 26350 34750 26402 34802
rect 26686 34750 26738 34802
rect 27022 34750 27074 34802
rect 32622 34750 32674 34802
rect 33518 34750 33570 34802
rect 33966 34750 34018 34802
rect 34302 34750 34354 34802
rect 34974 34750 35026 34802
rect 35310 34750 35362 34802
rect 34638 34638 34690 34690
rect 36430 34638 36482 34690
rect 10538 34470 10590 34522
rect 10642 34470 10694 34522
rect 10746 34470 10798 34522
rect 19862 34470 19914 34522
rect 19966 34470 20018 34522
rect 20070 34470 20122 34522
rect 29186 34470 29238 34522
rect 29290 34470 29342 34522
rect 29394 34470 29446 34522
rect 38510 34470 38562 34522
rect 38614 34470 38666 34522
rect 38718 34470 38770 34522
rect 33630 34302 33682 34354
rect 34750 34302 34802 34354
rect 34078 34190 34130 34242
rect 35422 34190 35474 34242
rect 36990 34190 37042 34242
rect 34414 34078 34466 34130
rect 35086 34078 35138 34130
rect 35982 33966 36034 34018
rect 5876 33686 5928 33738
rect 5980 33686 6032 33738
rect 6084 33686 6136 33738
rect 15200 33686 15252 33738
rect 15304 33686 15356 33738
rect 15408 33686 15460 33738
rect 24524 33686 24576 33738
rect 24628 33686 24680 33738
rect 24732 33686 24784 33738
rect 33848 33686 33900 33738
rect 33952 33686 34004 33738
rect 34056 33686 34108 33738
rect 35310 33406 35362 33458
rect 37550 33406 37602 33458
rect 38222 33406 38274 33458
rect 37102 33294 37154 33346
rect 34078 33182 34130 33234
rect 10538 32902 10590 32954
rect 10642 32902 10694 32954
rect 10746 32902 10798 32954
rect 19862 32902 19914 32954
rect 19966 32902 20018 32954
rect 20070 32902 20122 32954
rect 29186 32902 29238 32954
rect 29290 32902 29342 32954
rect 29394 32902 29446 32954
rect 38510 32902 38562 32954
rect 38614 32902 38666 32954
rect 38718 32902 38770 32954
rect 34974 32734 35026 32786
rect 37662 32734 37714 32786
rect 38222 32734 38274 32786
rect 35422 32622 35474 32674
rect 36990 32622 37042 32674
rect 35758 32398 35810 32450
rect 5876 32118 5928 32170
rect 5980 32118 6032 32170
rect 6084 32118 6136 32170
rect 15200 32118 15252 32170
rect 15304 32118 15356 32170
rect 15408 32118 15460 32170
rect 24524 32118 24576 32170
rect 24628 32118 24680 32170
rect 24732 32118 24784 32170
rect 33848 32118 33900 32170
rect 33952 32118 34004 32170
rect 34056 32118 34108 32170
rect 34302 31838 34354 31890
rect 36206 31726 36258 31778
rect 37326 31726 37378 31778
rect 35310 31614 35362 31666
rect 36430 31614 36482 31666
rect 37886 31614 37938 31666
rect 38222 31614 38274 31666
rect 37550 31502 37602 31554
rect 10538 31334 10590 31386
rect 10642 31334 10694 31386
rect 10746 31334 10798 31386
rect 19862 31334 19914 31386
rect 19966 31334 20018 31386
rect 20070 31334 20122 31386
rect 29186 31334 29238 31386
rect 29290 31334 29342 31386
rect 29394 31334 29446 31386
rect 38510 31334 38562 31386
rect 38614 31334 38666 31386
rect 38718 31334 38770 31386
rect 36430 31166 36482 31218
rect 36878 31166 36930 31218
rect 37214 31166 37266 31218
rect 37886 31166 37938 31218
rect 35422 31054 35474 31106
rect 38222 31054 38274 31106
rect 37438 30942 37490 30994
rect 34414 30830 34466 30882
rect 5876 30550 5928 30602
rect 5980 30550 6032 30602
rect 6084 30550 6136 30602
rect 15200 30550 15252 30602
rect 15304 30550 15356 30602
rect 15408 30550 15460 30602
rect 24524 30550 24576 30602
rect 24628 30550 24680 30602
rect 24732 30550 24784 30602
rect 33848 30550 33900 30602
rect 33952 30550 34004 30602
rect 34056 30550 34108 30602
rect 10446 30270 10498 30322
rect 14478 30270 14530 30322
rect 31054 30270 31106 30322
rect 34974 30270 35026 30322
rect 11454 30046 11506 30098
rect 15710 30046 15762 30098
rect 32062 30046 32114 30098
rect 36206 30046 36258 30098
rect 37102 30046 37154 30098
rect 37550 30046 37602 30098
rect 37886 30046 37938 30098
rect 38222 30046 38274 30098
rect 10538 29766 10590 29818
rect 10642 29766 10694 29818
rect 10746 29766 10798 29818
rect 19862 29766 19914 29818
rect 19966 29766 20018 29818
rect 20070 29766 20122 29818
rect 29186 29766 29238 29818
rect 29290 29766 29342 29818
rect 29394 29766 29446 29818
rect 38510 29766 38562 29818
rect 38614 29766 38666 29818
rect 38718 29766 38770 29818
rect 36766 29598 36818 29650
rect 37550 29598 37602 29650
rect 37886 29598 37938 29650
rect 13358 29486 13410 29538
rect 16270 29486 16322 29538
rect 29822 29486 29874 29538
rect 35198 29486 35250 29538
rect 38222 29374 38274 29426
rect 12350 29262 12402 29314
rect 15262 29262 15314 29314
rect 28478 29262 28530 29314
rect 34078 29262 34130 29314
rect 37214 29262 37266 29314
rect 5876 28982 5928 29034
rect 5980 28982 6032 29034
rect 6084 28982 6136 29034
rect 15200 28982 15252 29034
rect 15304 28982 15356 29034
rect 15408 28982 15460 29034
rect 24524 28982 24576 29034
rect 24628 28982 24680 29034
rect 24732 28982 24784 29034
rect 33848 28982 33900 29034
rect 33952 28982 34004 29034
rect 34056 28982 34108 29034
rect 9662 28702 9714 28754
rect 15262 28702 15314 28754
rect 18062 28702 18114 28754
rect 27022 28702 27074 28754
rect 30158 28702 30210 28754
rect 32958 28702 33010 28754
rect 37662 28590 37714 28642
rect 38110 28590 38162 28642
rect 10894 28478 10946 28530
rect 16606 28478 16658 28530
rect 19070 28478 19122 28530
rect 28030 28478 28082 28530
rect 31166 28478 31218 28530
rect 34190 28478 34242 28530
rect 37886 28478 37938 28530
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 14702 28030 14754 28082
rect 37886 28030 37938 28082
rect 7982 27918 8034 27970
rect 15262 27918 15314 27970
rect 19630 27918 19682 27970
rect 22318 27918 22370 27970
rect 29374 27918 29426 27970
rect 30158 27918 30210 27970
rect 35310 27918 35362 27970
rect 11790 27806 11842 27858
rect 12238 27806 12290 27858
rect 26686 27806 26738 27858
rect 27134 27806 27186 27858
rect 32286 27806 32338 27858
rect 38222 27806 38274 27858
rect 6974 27694 7026 27746
rect 10670 27694 10722 27746
rect 11006 27694 11058 27746
rect 18622 27694 18674 27746
rect 23438 27694 23490 27746
rect 32062 27694 32114 27746
rect 34302 27694 34354 27746
rect 37662 27694 37714 27746
rect 5876 27414 5928 27466
rect 5980 27414 6032 27466
rect 6084 27414 6136 27466
rect 15200 27414 15252 27466
rect 15304 27414 15356 27466
rect 15408 27414 15460 27466
rect 24524 27414 24576 27466
rect 24628 27414 24680 27466
rect 24732 27414 24784 27466
rect 33848 27414 33900 27466
rect 33952 27414 34004 27466
rect 34056 27414 34108 27466
rect 12462 27246 12514 27298
rect 18286 27246 18338 27298
rect 26014 27246 26066 27298
rect 30382 27246 30434 27298
rect 7086 27134 7138 27186
rect 29374 27134 29426 27186
rect 8990 27022 9042 27074
rect 9438 27022 9490 27074
rect 13694 27022 13746 27074
rect 14590 27022 14642 27074
rect 15262 27022 15314 27074
rect 22318 27022 22370 27074
rect 22990 27022 23042 27074
rect 33518 27022 33570 27074
rect 34078 27022 34130 27074
rect 8094 26910 8146 26962
rect 11678 26910 11730 26962
rect 13470 26910 13522 26962
rect 18846 26910 18898 26962
rect 29150 26910 29202 26962
rect 37774 26910 37826 26962
rect 17502 26798 17554 26850
rect 18958 26798 19010 26850
rect 25454 26798 25506 26850
rect 31166 26798 31218 26850
rect 36990 26798 37042 26850
rect 10538 26630 10590 26682
rect 10642 26630 10694 26682
rect 10746 26630 10798 26682
rect 19862 26630 19914 26682
rect 19966 26630 20018 26682
rect 20070 26630 20122 26682
rect 29186 26630 29238 26682
rect 29290 26630 29342 26682
rect 29394 26630 29446 26682
rect 38510 26630 38562 26682
rect 38614 26630 38666 26682
rect 38718 26630 38770 26682
rect 8318 26462 8370 26514
rect 9102 26462 9154 26514
rect 16046 26462 16098 26514
rect 16382 26462 16434 26514
rect 21086 26462 21138 26514
rect 28814 26462 28866 26514
rect 31838 26462 31890 26514
rect 32622 26462 32674 26514
rect 32958 26462 33010 26514
rect 33630 26462 33682 26514
rect 37886 26462 37938 26514
rect 2382 26350 2434 26402
rect 9774 26350 9826 26402
rect 15262 26350 15314 26402
rect 20414 26350 20466 26402
rect 21870 26350 21922 26402
rect 28030 26350 28082 26402
rect 37550 26350 37602 26402
rect 38222 26350 38274 26402
rect 4622 26238 4674 26290
rect 5294 26238 5346 26290
rect 5630 26238 5682 26290
rect 6078 26238 6130 26290
rect 12574 26238 12626 26290
rect 13022 26238 13074 26290
rect 24222 26238 24274 26290
rect 24670 26238 24722 26290
rect 25342 26238 25394 26290
rect 25790 26238 25842 26290
rect 29150 26238 29202 26290
rect 29598 26238 29650 26290
rect 35982 26238 36034 26290
rect 36430 26238 36482 26290
rect 11118 26126 11170 26178
rect 16270 26126 16322 26178
rect 19406 26126 19458 26178
rect 1598 26014 1650 26066
rect 5876 25846 5928 25898
rect 5980 25846 6032 25898
rect 6084 25846 6136 25898
rect 15200 25846 15252 25898
rect 15304 25846 15356 25898
rect 15408 25846 15460 25898
rect 24524 25846 24576 25898
rect 24628 25846 24680 25898
rect 24732 25846 24784 25898
rect 33848 25846 33900 25898
rect 33952 25846 34004 25898
rect 34056 25846 34108 25898
rect 5518 25678 5570 25730
rect 13022 25678 13074 25730
rect 32734 25678 32786 25730
rect 36542 25678 36594 25730
rect 3502 25566 3554 25618
rect 14142 25566 14194 25618
rect 15934 25566 15986 25618
rect 22430 25566 22482 25618
rect 25566 25566 25618 25618
rect 27694 25566 27746 25618
rect 38334 25566 38386 25618
rect 8654 25454 8706 25506
rect 8990 25454 9042 25506
rect 9326 25454 9378 25506
rect 9998 25454 10050 25506
rect 17166 25454 17218 25506
rect 17838 25454 17890 25506
rect 27470 25454 27522 25506
rect 29262 25454 29314 25506
rect 29710 25454 29762 25506
rect 33070 25454 33122 25506
rect 33406 25454 33458 25506
rect 37214 25454 37266 25506
rect 2158 25342 2210 25394
rect 6302 25342 6354 25394
rect 13806 25342 13858 25394
rect 14926 25342 14978 25394
rect 20862 25342 20914 25394
rect 23550 25342 23602 25394
rect 26574 25342 26626 25394
rect 36990 25342 37042 25394
rect 12462 25230 12514 25282
rect 20190 25230 20242 25282
rect 32062 25230 32114 25282
rect 35982 25230 36034 25282
rect 10538 25062 10590 25114
rect 10642 25062 10694 25114
rect 10746 25062 10798 25114
rect 19862 25062 19914 25114
rect 19966 25062 20018 25114
rect 20070 25062 20122 25114
rect 29186 25062 29238 25114
rect 29290 25062 29342 25114
rect 29394 25062 29446 25114
rect 38510 25062 38562 25114
rect 38614 25062 38666 25114
rect 38718 25062 38770 25114
rect 7870 24894 7922 24946
rect 8430 24894 8482 24946
rect 15038 24894 15090 24946
rect 18510 24894 18562 24946
rect 29598 24894 29650 24946
rect 30158 24894 30210 24946
rect 30494 24894 30546 24946
rect 38222 24894 38274 24946
rect 2270 24782 2322 24834
rect 10110 24782 10162 24834
rect 14254 24782 14306 24834
rect 17502 24782 17554 24834
rect 19294 24782 19346 24834
rect 25230 24782 25282 24834
rect 25902 24782 25954 24834
rect 32062 24782 32114 24834
rect 33182 24782 33234 24834
rect 33966 24782 34018 24834
rect 37438 24782 37490 24834
rect 4958 24670 5010 24722
rect 5294 24670 5346 24722
rect 10334 24670 10386 24722
rect 11006 24670 11058 24722
rect 11454 24670 11506 24722
rect 11902 24670 11954 24722
rect 17726 24670 17778 24722
rect 21646 24670 21698 24722
rect 22206 24670 22258 24722
rect 26686 24670 26738 24722
rect 27134 24670 27186 24722
rect 31838 24670 31890 24722
rect 33406 24670 33458 24722
rect 34190 24670 34242 24722
rect 34526 24670 34578 24722
rect 35198 24670 35250 24722
rect 3502 24558 3554 24610
rect 10894 24558 10946 24610
rect 25566 24558 25618 24610
rect 26238 24558 26290 24610
rect 30382 24558 30434 24610
rect 5876 24278 5928 24330
rect 5980 24278 6032 24330
rect 6084 24278 6136 24330
rect 15200 24278 15252 24330
rect 15304 24278 15356 24330
rect 15408 24278 15460 24330
rect 24524 24278 24576 24330
rect 24628 24278 24680 24330
rect 24732 24278 24784 24330
rect 33848 24278 33900 24330
rect 33952 24278 34004 24330
rect 34056 24278 34108 24330
rect 9102 24110 9154 24162
rect 19742 24110 19794 24162
rect 2270 23998 2322 24050
rect 4062 23998 4114 24050
rect 7646 23998 7698 24050
rect 13470 23998 13522 24050
rect 20190 23998 20242 24050
rect 21310 23998 21362 24050
rect 30158 23998 30210 24050
rect 32958 23998 33010 24050
rect 36990 23998 37042 24050
rect 37326 23998 37378 24050
rect 12126 23886 12178 23938
rect 12574 23886 12626 23938
rect 13694 23886 13746 23938
rect 16046 23886 16098 23938
rect 16718 23886 16770 23938
rect 20302 23886 20354 23938
rect 21534 23886 21586 23938
rect 23438 23886 23490 23938
rect 23998 23886 24050 23938
rect 28254 23886 28306 23938
rect 1934 23774 1986 23826
rect 2942 23774 2994 23826
rect 5742 23774 5794 23826
rect 6638 23774 6690 23826
rect 18958 23774 19010 23826
rect 27246 23774 27298 23826
rect 27582 23774 27634 23826
rect 31166 23774 31218 23826
rect 33966 23774 34018 23826
rect 5854 23662 5906 23714
rect 9886 23662 9938 23714
rect 26462 23662 26514 23714
rect 27022 23662 27074 23714
rect 28254 23662 28306 23714
rect 10538 23494 10590 23546
rect 10642 23494 10694 23546
rect 10746 23494 10798 23546
rect 19862 23494 19914 23546
rect 19966 23494 20018 23546
rect 20070 23494 20122 23546
rect 29186 23494 29238 23546
rect 29290 23494 29342 23546
rect 29394 23494 29446 23546
rect 38510 23494 38562 23546
rect 38614 23494 38666 23546
rect 38718 23494 38770 23546
rect 2942 23326 2994 23378
rect 3726 23326 3778 23378
rect 24222 23326 24274 23378
rect 24782 23326 24834 23378
rect 36094 23326 36146 23378
rect 36654 23326 36706 23378
rect 6862 23214 6914 23266
rect 7534 23214 7586 23266
rect 7870 23214 7922 23266
rect 17726 23214 17778 23266
rect 20414 23214 20466 23266
rect 5966 23102 6018 23154
rect 6414 23102 6466 23154
rect 14702 23102 14754 23154
rect 21310 23102 21362 23154
rect 21758 23102 21810 23154
rect 29374 23102 29426 23154
rect 33182 23102 33234 23154
rect 33630 23102 33682 23154
rect 7086 22990 7138 23042
rect 10334 22990 10386 23042
rect 15374 22990 15426 23042
rect 17390 22990 17442 23042
rect 19406 22990 19458 23042
rect 26910 22990 26962 23042
rect 31390 22990 31442 23042
rect 5876 22710 5928 22762
rect 5980 22710 6032 22762
rect 6084 22710 6136 22762
rect 15200 22710 15252 22762
rect 15304 22710 15356 22762
rect 15408 22710 15460 22762
rect 24524 22710 24576 22762
rect 24628 22710 24680 22762
rect 24732 22710 24784 22762
rect 33848 22710 33900 22762
rect 33952 22710 34004 22762
rect 34056 22710 34108 22762
rect 9326 22542 9378 22594
rect 1934 22430 1986 22482
rect 4062 22430 4114 22482
rect 16046 22430 16098 22482
rect 26462 22430 26514 22482
rect 28366 22430 28418 22482
rect 29710 22430 29762 22482
rect 33182 22430 33234 22482
rect 36990 22430 37042 22482
rect 37662 22430 37714 22482
rect 8654 22318 8706 22370
rect 9214 22318 9266 22370
rect 12350 22318 12402 22370
rect 12798 22318 12850 22370
rect 15486 22318 15538 22370
rect 20638 22318 20690 22370
rect 21758 22318 21810 22370
rect 22206 22318 22258 22370
rect 29262 22318 29314 22370
rect 31166 22318 31218 22370
rect 37214 22318 37266 22370
rect 2270 22206 2322 22258
rect 3054 22206 3106 22258
rect 20414 22206 20466 22258
rect 27470 22206 27522 22258
rect 28590 22206 28642 22258
rect 30830 22206 30882 22258
rect 5518 22094 5570 22146
rect 6078 22094 6130 22146
rect 10110 22094 10162 22146
rect 19742 22094 19794 22146
rect 24558 22094 24610 22146
rect 25230 22094 25282 22146
rect 25566 22094 25618 22146
rect 37774 22094 37826 22146
rect 10538 21926 10590 21978
rect 10642 21926 10694 21978
rect 10746 21926 10798 21978
rect 19862 21926 19914 21978
rect 19966 21926 20018 21978
rect 20070 21926 20122 21978
rect 29186 21926 29238 21978
rect 29290 21926 29342 21978
rect 29394 21926 29446 21978
rect 38510 21926 38562 21978
rect 38614 21926 38666 21978
rect 38718 21926 38770 21978
rect 1598 21758 1650 21810
rect 2270 21758 2322 21810
rect 8542 21758 8594 21810
rect 9662 21758 9714 21810
rect 14030 21758 14082 21810
rect 22766 21758 22818 21810
rect 24558 21758 24610 21810
rect 28254 21758 28306 21810
rect 28814 21758 28866 21810
rect 32062 21758 32114 21810
rect 37662 21758 37714 21810
rect 38222 21758 38274 21810
rect 9102 21646 9154 21698
rect 12910 21646 12962 21698
rect 18510 21646 18562 21698
rect 21982 21646 22034 21698
rect 33070 21646 33122 21698
rect 33406 21646 33458 21698
rect 33854 21646 33906 21698
rect 4734 21534 4786 21586
rect 5070 21534 5122 21586
rect 5406 21534 5458 21586
rect 5966 21534 6018 21586
rect 16270 21534 16322 21586
rect 16718 21534 16770 21586
rect 17838 21534 17890 21586
rect 19294 21534 19346 21586
rect 19630 21534 19682 21586
rect 25342 21534 25394 21586
rect 25790 21534 25842 21586
rect 28926 21534 28978 21586
rect 29598 21534 29650 21586
rect 34526 21534 34578 21586
rect 35198 21534 35250 21586
rect 9550 21422 9602 21474
rect 11566 21422 11618 21474
rect 17614 21422 17666 21474
rect 18734 21422 18786 21474
rect 24670 21422 24722 21474
rect 34190 21422 34242 21474
rect 13246 21310 13298 21362
rect 32622 21310 32674 21362
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 6974 20974 7026 21026
rect 11454 20974 11506 21026
rect 12686 20974 12738 21026
rect 19518 20974 19570 21026
rect 34750 20974 34802 21026
rect 3838 20862 3890 20914
rect 13918 20862 13970 20914
rect 14254 20862 14306 20914
rect 14590 20862 14642 20914
rect 21758 20862 21810 20914
rect 5966 20750 6018 20802
rect 7758 20750 7810 20802
rect 8430 20750 8482 20802
rect 11902 20750 11954 20802
rect 14814 20750 14866 20802
rect 16046 20750 16098 20802
rect 16382 20750 16434 20802
rect 22318 20750 22370 20802
rect 26574 20750 26626 20802
rect 26910 20750 26962 20802
rect 27582 20750 27634 20802
rect 29822 20750 29874 20802
rect 31054 20750 31106 20802
rect 31614 20750 31666 20802
rect 3054 20638 3106 20690
rect 5630 20638 5682 20690
rect 7534 20638 7586 20690
rect 18734 20638 18786 20690
rect 27358 20638 27410 20690
rect 28254 20638 28306 20690
rect 28590 20638 28642 20690
rect 30382 20638 30434 20690
rect 34974 20638 35026 20690
rect 10894 20526 10946 20578
rect 13582 20526 13634 20578
rect 22990 20526 23042 20578
rect 23438 20526 23490 20578
rect 24222 20526 24274 20578
rect 34190 20526 34242 20578
rect 35086 20526 35138 20578
rect 38334 20526 38386 20578
rect 10538 20358 10590 20410
rect 10642 20358 10694 20410
rect 10746 20358 10798 20410
rect 19862 20358 19914 20410
rect 19966 20358 20018 20410
rect 20070 20358 20122 20410
rect 29186 20358 29238 20410
rect 29290 20358 29342 20410
rect 29394 20358 29446 20410
rect 38510 20358 38562 20410
rect 38614 20358 38666 20410
rect 38718 20358 38770 20410
rect 7086 20190 7138 20242
rect 16382 20190 16434 20242
rect 20414 20190 20466 20242
rect 36766 20190 36818 20242
rect 3838 20078 3890 20130
rect 11006 20078 11058 20130
rect 21310 20078 21362 20130
rect 21646 20078 21698 20130
rect 24222 20078 24274 20130
rect 26798 20078 26850 20130
rect 30606 20078 30658 20130
rect 31950 20078 32002 20130
rect 37886 20078 37938 20130
rect 38222 20078 38274 20130
rect 3614 19966 3666 20018
rect 4174 19966 4226 20018
rect 4734 19966 4786 20018
rect 8094 19966 8146 20018
rect 13358 19966 13410 20018
rect 13806 19966 13858 20018
rect 17278 19966 17330 20018
rect 17950 19966 18002 20018
rect 29150 19966 29202 20018
rect 29486 19966 29538 20018
rect 33294 19966 33346 20018
rect 33742 19966 33794 20018
rect 34302 19966 34354 20018
rect 8318 19854 8370 19906
rect 8766 19854 8818 19906
rect 12014 19854 12066 19906
rect 22094 19854 22146 19906
rect 23214 19854 23266 19906
rect 30942 19854 30994 19906
rect 33070 19854 33122 19906
rect 7758 19742 7810 19794
rect 16942 19742 16994 19794
rect 20974 19742 21026 19794
rect 26014 19742 26066 19794
rect 37326 19742 37378 19794
rect 5876 19574 5928 19626
rect 5980 19574 6032 19626
rect 6084 19574 6136 19626
rect 15200 19574 15252 19626
rect 15304 19574 15356 19626
rect 15408 19574 15460 19626
rect 24524 19574 24576 19626
rect 24628 19574 24680 19626
rect 24732 19574 24784 19626
rect 33848 19574 33900 19626
rect 33952 19574 34004 19626
rect 34056 19574 34108 19626
rect 13358 19406 13410 19458
rect 4062 19294 4114 19346
rect 12462 19294 12514 19346
rect 17726 19294 17778 19346
rect 19518 19294 19570 19346
rect 36990 19294 37042 19346
rect 37326 19294 37378 19346
rect 37662 19294 37714 19346
rect 5854 19182 5906 19234
rect 9998 19182 10050 19234
rect 10446 19182 10498 19234
rect 12686 19182 12738 19234
rect 16382 19182 16434 19234
rect 17054 19182 17106 19234
rect 22094 19182 22146 19234
rect 27918 19182 27970 19234
rect 28590 19182 28642 19234
rect 29262 19182 29314 19234
rect 29710 19182 29762 19234
rect 32958 19182 33010 19234
rect 33518 19182 33570 19234
rect 3054 19070 3106 19122
rect 11118 19070 11170 19122
rect 11454 19070 11506 19122
rect 11790 19070 11842 19122
rect 12126 19070 12178 19122
rect 17390 19070 17442 19122
rect 20638 19070 20690 19122
rect 23774 19070 23826 19122
rect 35758 19070 35810 19122
rect 5854 18958 5906 19010
rect 6974 18958 7026 19010
rect 7758 18958 7810 19010
rect 14142 18958 14194 19010
rect 27582 18958 27634 19010
rect 32174 18958 32226 19010
rect 32734 18958 32786 19010
rect 36542 18958 36594 19010
rect 37774 18958 37826 19010
rect 10538 18790 10590 18842
rect 10642 18790 10694 18842
rect 10746 18790 10798 18842
rect 19862 18790 19914 18842
rect 19966 18790 20018 18842
rect 20070 18790 20122 18842
rect 29186 18790 29238 18842
rect 29290 18790 29342 18842
rect 29394 18790 29446 18842
rect 38510 18790 38562 18842
rect 38614 18790 38666 18842
rect 38718 18790 38770 18842
rect 8318 18622 8370 18674
rect 12350 18622 12402 18674
rect 30382 18622 30434 18674
rect 36094 18622 36146 18674
rect 3054 18510 3106 18562
rect 11006 18510 11058 18562
rect 21870 18510 21922 18562
rect 29150 18510 29202 18562
rect 30718 18510 30770 18562
rect 37214 18510 37266 18562
rect 37550 18510 37602 18562
rect 5294 18398 5346 18450
rect 5854 18398 5906 18450
rect 14926 18398 14978 18450
rect 15486 18398 15538 18450
rect 18958 18398 19010 18450
rect 19518 18398 19570 18450
rect 26350 18398 26402 18450
rect 26910 18398 26962 18450
rect 32958 18398 33010 18450
rect 33630 18398 33682 18450
rect 36878 18398 36930 18450
rect 4062 18286 4114 18338
rect 8990 18286 9042 18338
rect 9774 18286 9826 18338
rect 10110 18286 10162 18338
rect 10334 18286 10386 18338
rect 10782 18286 10834 18338
rect 11566 18286 11618 18338
rect 15710 18286 15762 18338
rect 16046 18286 16098 18338
rect 17614 18286 17666 18338
rect 18062 18286 18114 18338
rect 22878 18286 22930 18338
rect 23214 18286 23266 18338
rect 23550 18286 23602 18338
rect 23886 18286 23938 18338
rect 31726 18286 31778 18338
rect 37886 18286 37938 18338
rect 11790 18174 11842 18226
rect 22654 18174 22706 18226
rect 29934 18174 29986 18226
rect 36654 18174 36706 18226
rect 5876 18006 5928 18058
rect 5980 18006 6032 18058
rect 6084 18006 6136 18058
rect 15200 18006 15252 18058
rect 15304 18006 15356 18058
rect 15408 18006 15460 18058
rect 24524 18006 24576 18058
rect 24628 18006 24680 18058
rect 24732 18006 24784 18058
rect 33848 18006 33900 18058
rect 33952 18006 34004 18058
rect 34056 18006 34108 18058
rect 3950 17726 4002 17778
rect 21758 17726 21810 17778
rect 27358 17726 27410 17778
rect 37550 17726 37602 17778
rect 8654 17614 8706 17666
rect 9102 17614 9154 17666
rect 9326 17614 9378 17666
rect 9886 17614 9938 17666
rect 13582 17614 13634 17666
rect 13918 17614 13970 17666
rect 20190 17614 20242 17666
rect 20638 17614 20690 17666
rect 22206 17614 22258 17666
rect 22878 17614 22930 17666
rect 32174 17614 32226 17666
rect 32734 17614 32786 17666
rect 32846 17614 32898 17666
rect 33518 17614 33570 17666
rect 38222 17614 38274 17666
rect 3054 17502 3106 17554
rect 5518 17502 5570 17554
rect 16270 17502 16322 17554
rect 17950 17502 18002 17554
rect 21982 17502 22034 17554
rect 26238 17502 26290 17554
rect 1822 17390 1874 17442
rect 6190 17390 6242 17442
rect 12462 17390 12514 17442
rect 13022 17390 13074 17442
rect 17054 17390 17106 17442
rect 17166 17390 17218 17442
rect 25230 17390 25282 17442
rect 25902 17390 25954 17442
rect 29038 17390 29090 17442
rect 29822 17390 29874 17442
rect 35982 17390 36034 17442
rect 36542 17390 36594 17442
rect 10538 17222 10590 17274
rect 10642 17222 10694 17274
rect 10746 17222 10798 17274
rect 19862 17222 19914 17274
rect 19966 17222 20018 17274
rect 20070 17222 20122 17274
rect 29186 17222 29238 17274
rect 29290 17222 29342 17274
rect 29394 17222 29446 17274
rect 38510 17222 38562 17274
rect 38614 17222 38666 17274
rect 38718 17222 38770 17274
rect 4958 17054 5010 17106
rect 8990 17054 9042 17106
rect 14030 17054 14082 17106
rect 15262 17054 15314 17106
rect 23550 17054 23602 17106
rect 37214 17054 37266 17106
rect 6190 16942 6242 16994
rect 6974 16942 7026 16994
rect 10782 16942 10834 16994
rect 17838 16942 17890 16994
rect 24110 16942 24162 16994
rect 24670 16942 24722 16994
rect 25230 16942 25282 16994
rect 25566 16942 25618 16994
rect 28926 16942 28978 16994
rect 31950 16942 32002 16994
rect 33070 16942 33122 16994
rect 2158 16830 2210 16882
rect 2606 16830 2658 16882
rect 5966 16830 6018 16882
rect 9998 16830 10050 16882
rect 11342 16830 11394 16882
rect 11790 16830 11842 16882
rect 16718 16830 16770 16882
rect 20638 16830 20690 16882
rect 21086 16830 21138 16882
rect 26014 16830 26066 16882
rect 26574 16830 26626 16882
rect 33294 16830 33346 16882
rect 34302 16830 34354 16882
rect 34750 16830 34802 16882
rect 7982 16718 8034 16770
rect 8542 16718 8594 16770
rect 16046 16718 16098 16770
rect 19182 16718 19234 16770
rect 24334 16718 24386 16770
rect 30606 16718 30658 16770
rect 30942 16718 30994 16770
rect 5630 16606 5682 16658
rect 14814 16606 14866 16658
rect 29710 16606 29762 16658
rect 37774 16606 37826 16658
rect 5876 16438 5928 16490
rect 5980 16438 6032 16490
rect 6084 16438 6136 16490
rect 15200 16438 15252 16490
rect 15304 16438 15356 16490
rect 15408 16438 15460 16490
rect 24524 16438 24576 16490
rect 24628 16438 24680 16490
rect 24732 16438 24784 16490
rect 33848 16438 33900 16490
rect 33952 16438 34004 16490
rect 34056 16438 34108 16490
rect 23438 16270 23490 16322
rect 4062 16158 4114 16210
rect 7534 16158 7586 16210
rect 15934 16158 15986 16210
rect 21646 16158 21698 16210
rect 21982 16158 22034 16210
rect 27582 16158 27634 16210
rect 28478 16158 28530 16210
rect 30158 16158 30210 16210
rect 5854 16046 5906 16098
rect 7758 16046 7810 16098
rect 8318 16046 8370 16098
rect 12798 16046 12850 16098
rect 14142 16046 14194 16098
rect 16382 16046 16434 16098
rect 16718 16046 16770 16098
rect 26574 16046 26626 16098
rect 26910 16046 26962 16098
rect 28366 16046 28418 16098
rect 30830 16046 30882 16098
rect 31278 16046 31330 16098
rect 37214 16046 37266 16098
rect 1710 15934 1762 15986
rect 3054 15934 3106 15986
rect 5630 15934 5682 15986
rect 12126 15934 12178 15986
rect 14702 15934 14754 15986
rect 20078 15934 20130 15986
rect 20414 15934 20466 15986
rect 34638 15934 34690 15986
rect 36990 15934 37042 15986
rect 37662 15934 37714 15986
rect 2046 15822 2098 15874
rect 5070 15822 5122 15874
rect 6414 15822 6466 15874
rect 7422 15822 7474 15874
rect 10894 15822 10946 15874
rect 11454 15822 11506 15874
rect 13582 15822 13634 15874
rect 19294 15822 19346 15874
rect 19854 15822 19906 15874
rect 24222 15822 24274 15874
rect 27694 15822 27746 15874
rect 37774 15822 37826 15874
rect 10538 15654 10590 15706
rect 10642 15654 10694 15706
rect 10746 15654 10798 15706
rect 19862 15654 19914 15706
rect 19966 15654 20018 15706
rect 20070 15654 20122 15706
rect 29186 15654 29238 15706
rect 29290 15654 29342 15706
rect 29394 15654 29446 15706
rect 38510 15654 38562 15706
rect 38614 15654 38666 15706
rect 38718 15654 38770 15706
rect 2382 15486 2434 15538
rect 5966 15486 6018 15538
rect 16718 15486 16770 15538
rect 18958 15486 19010 15538
rect 22766 15486 22818 15538
rect 33742 15486 33794 15538
rect 12798 15374 12850 15426
rect 24110 15374 24162 15426
rect 4622 15262 4674 15314
rect 5294 15262 5346 15314
rect 8542 15262 8594 15314
rect 9102 15262 9154 15314
rect 14814 15262 14866 15314
rect 15374 15262 15426 15314
rect 16046 15262 16098 15314
rect 21310 15262 21362 15314
rect 21646 15262 21698 15314
rect 29374 15262 29426 15314
rect 31502 15262 31554 15314
rect 35982 15262 36034 15314
rect 36430 15262 36482 15314
rect 15150 15150 15202 15202
rect 16270 15150 16322 15202
rect 17502 15150 17554 15202
rect 17838 15150 17890 15202
rect 23102 15150 23154 15202
rect 25790 15150 25842 15202
rect 32958 15150 33010 15202
rect 1598 15038 1650 15090
rect 5406 15038 5458 15090
rect 18174 15038 18226 15090
rect 32286 15038 32338 15090
rect 5876 14870 5928 14922
rect 5980 14870 6032 14922
rect 6084 14870 6136 14922
rect 15200 14870 15252 14922
rect 15304 14870 15356 14922
rect 15408 14870 15460 14922
rect 24524 14870 24576 14922
rect 24628 14870 24680 14922
rect 24732 14870 24784 14922
rect 33848 14870 33900 14922
rect 33952 14870 34004 14922
rect 34056 14870 34108 14922
rect 3614 14590 3666 14642
rect 5854 14590 5906 14642
rect 8094 14590 8146 14642
rect 16830 14590 16882 14642
rect 19518 14590 19570 14642
rect 19966 14590 20018 14642
rect 28478 14590 28530 14642
rect 12350 14478 12402 14530
rect 12910 14478 12962 14530
rect 13806 14478 13858 14530
rect 26798 14478 26850 14530
rect 27134 14478 27186 14530
rect 28366 14478 28418 14530
rect 29038 14478 29090 14530
rect 29710 14478 29762 14530
rect 32846 14478 32898 14530
rect 33406 14478 33458 14530
rect 37214 14478 37266 14530
rect 1934 14366 1986 14418
rect 4958 14366 5010 14418
rect 5630 14366 5682 14418
rect 7086 14366 7138 14418
rect 10110 14366 10162 14418
rect 27582 14366 27634 14418
rect 27918 14366 27970 14418
rect 36990 14366 37042 14418
rect 2046 14254 2098 14306
rect 8654 14254 8706 14306
rect 9102 14254 9154 14306
rect 9326 14254 9378 14306
rect 23662 14254 23714 14306
rect 24334 14254 24386 14306
rect 32174 14254 32226 14306
rect 32734 14254 32786 14306
rect 35982 14254 36034 14306
rect 36542 14254 36594 14306
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 4734 13918 4786 13970
rect 8318 13918 8370 13970
rect 16382 13918 16434 13970
rect 20414 13918 20466 13970
rect 24222 13918 24274 13970
rect 28030 13918 28082 13970
rect 37774 13918 37826 13970
rect 38334 13918 38386 13970
rect 12350 13806 12402 13858
rect 31838 13806 31890 13858
rect 33070 13806 33122 13858
rect 33742 13806 33794 13858
rect 1822 13694 1874 13746
rect 2270 13694 2322 13746
rect 5630 13694 5682 13746
rect 6078 13694 6130 13746
rect 9438 13694 9490 13746
rect 10110 13694 10162 13746
rect 13358 13694 13410 13746
rect 13918 13694 13970 13746
rect 17278 13694 17330 13746
rect 17950 13694 18002 13746
rect 21086 13694 21138 13746
rect 21758 13694 21810 13746
rect 25230 13694 25282 13746
rect 25678 13694 25730 13746
rect 29038 13694 29090 13746
rect 29598 13694 29650 13746
rect 33294 13694 33346 13746
rect 33966 13694 34018 13746
rect 34638 13694 34690 13746
rect 35198 13694 35250 13746
rect 5294 13470 5346 13522
rect 9102 13470 9154 13522
rect 13134 13470 13186 13522
rect 16942 13470 16994 13522
rect 20974 13470 21026 13522
rect 24782 13470 24834 13522
rect 28814 13470 28866 13522
rect 32622 13470 32674 13522
rect 5876 13302 5928 13354
rect 5980 13302 6032 13354
rect 6084 13302 6136 13354
rect 15200 13302 15252 13354
rect 15304 13302 15356 13354
rect 15408 13302 15460 13354
rect 24524 13302 24576 13354
rect 24628 13302 24680 13354
rect 24732 13302 24784 13354
rect 33848 13302 33900 13354
rect 33952 13302 34004 13354
rect 34056 13302 34108 13354
rect 1934 13022 1986 13074
rect 3838 13022 3890 13074
rect 12462 13022 12514 13074
rect 13022 13022 13074 13074
rect 22206 13022 22258 13074
rect 34526 13022 34578 13074
rect 37662 13022 37714 13074
rect 5966 12910 6018 12962
rect 7646 12910 7698 12962
rect 8206 12910 8258 12962
rect 13470 12910 13522 12962
rect 13918 12910 13970 12962
rect 20190 12910 20242 12962
rect 20862 12910 20914 12962
rect 22430 12910 22482 12962
rect 23214 12910 23266 12962
rect 23886 12910 23938 12962
rect 32622 12910 32674 12962
rect 33070 12910 33122 12962
rect 37214 12910 37266 12962
rect 2270 12798 2322 12850
rect 4958 12798 5010 12850
rect 6190 12798 6242 12850
rect 6526 12798 6578 12850
rect 6862 12798 6914 12850
rect 12126 12798 12178 12850
rect 16270 12798 16322 12850
rect 17950 12798 18002 12850
rect 21534 12798 21586 12850
rect 21870 12798 21922 12850
rect 35534 12798 35586 12850
rect 7310 12686 7362 12738
rect 10558 12686 10610 12738
rect 11342 12686 11394 12738
rect 11678 12686 11730 12738
rect 17054 12686 17106 12738
rect 17166 12686 17218 12738
rect 26126 12686 26178 12738
rect 26910 12686 26962 12738
rect 29598 12686 29650 12738
rect 30382 12686 30434 12738
rect 37214 12686 37266 12738
rect 37774 12686 37826 12738
rect 10538 12518 10590 12570
rect 10642 12518 10694 12570
rect 10746 12518 10798 12570
rect 19862 12518 19914 12570
rect 19966 12518 20018 12570
rect 20070 12518 20122 12570
rect 29186 12518 29238 12570
rect 29290 12518 29342 12570
rect 29394 12518 29446 12570
rect 38510 12518 38562 12570
rect 38614 12518 38666 12570
rect 38718 12518 38770 12570
rect 4510 12350 4562 12402
rect 16382 12350 16434 12402
rect 22206 12350 22258 12402
rect 36990 12350 37042 12402
rect 37886 12350 37938 12402
rect 8318 12238 8370 12290
rect 12798 12238 12850 12290
rect 17726 12238 17778 12290
rect 24222 12238 24274 12290
rect 24558 12238 24610 12290
rect 26014 12238 26066 12290
rect 28590 12238 28642 12290
rect 31726 12238 31778 12290
rect 33294 12238 33346 12290
rect 33630 12238 33682 12290
rect 37774 12238 37826 12290
rect 1822 12126 1874 12178
rect 2158 12126 2210 12178
rect 5630 12126 5682 12178
rect 5966 12126 6018 12178
rect 13470 12126 13522 12178
rect 13918 12126 13970 12178
rect 17950 12126 18002 12178
rect 19294 12126 19346 12178
rect 19966 12126 20018 12178
rect 23326 12126 23378 12178
rect 33854 12126 33906 12178
rect 34526 12126 34578 12178
rect 9886 12014 9938 12066
rect 10110 12014 10162 12066
rect 10670 12014 10722 12066
rect 11230 12014 11282 12066
rect 11790 12014 11842 12066
rect 18734 12014 18786 12066
rect 19070 12014 19122 12066
rect 23438 12014 23490 12066
rect 25678 12014 25730 12066
rect 27358 12014 27410 12066
rect 30494 12014 30546 12066
rect 5294 11902 5346 11954
rect 9102 11902 9154 11954
rect 10670 11902 10722 11954
rect 11230 11902 11282 11954
rect 16942 11902 16994 11954
rect 22990 11902 23042 11954
rect 37550 11902 37602 11954
rect 5876 11734 5928 11786
rect 5980 11734 6032 11786
rect 6084 11734 6136 11786
rect 15200 11734 15252 11786
rect 15304 11734 15356 11786
rect 15408 11734 15460 11786
rect 24524 11734 24576 11786
rect 24628 11734 24680 11786
rect 24732 11734 24784 11786
rect 33848 11734 33900 11786
rect 33952 11734 34004 11786
rect 34056 11734 34108 11786
rect 4062 11454 4114 11506
rect 7870 11454 7922 11506
rect 12350 11454 12402 11506
rect 15374 11454 15426 11506
rect 15934 11454 15986 11506
rect 16382 11454 16434 11506
rect 22318 11454 22370 11506
rect 25118 11454 25170 11506
rect 34302 11454 34354 11506
rect 38110 11454 38162 11506
rect 8094 11342 8146 11394
rect 8654 11342 8706 11394
rect 16830 11342 16882 11394
rect 17166 11342 17218 11394
rect 33294 11342 33346 11394
rect 33742 11342 33794 11394
rect 36990 11342 37042 11394
rect 2942 11230 2994 11282
rect 7534 11230 7586 11282
rect 12126 11230 12178 11282
rect 14366 11230 14418 11282
rect 19518 11230 19570 11282
rect 23550 11230 23602 11282
rect 26126 11230 26178 11282
rect 34526 11230 34578 11282
rect 35758 11230 35810 11282
rect 36430 11230 36482 11282
rect 5742 11118 5794 11170
rect 11006 11118 11058 11170
rect 11790 11118 11842 11170
rect 12910 11118 12962 11170
rect 13582 11118 13634 11170
rect 20302 11118 20354 11170
rect 20638 11118 20690 11170
rect 30270 11118 30322 11170
rect 31054 11118 31106 11170
rect 35198 11118 35250 11170
rect 35422 11118 35474 11170
rect 36094 11118 36146 11170
rect 10538 10950 10590 11002
rect 10642 10950 10694 11002
rect 10746 10950 10798 11002
rect 19862 10950 19914 11002
rect 19966 10950 20018 11002
rect 20070 10950 20122 11002
rect 29186 10950 29238 11002
rect 29290 10950 29342 11002
rect 29394 10950 29446 11002
rect 38510 10950 38562 11002
rect 38614 10950 38666 11002
rect 38718 10950 38770 11002
rect 5518 10782 5570 10834
rect 8766 10782 8818 10834
rect 9774 10782 9826 10834
rect 12238 10782 12290 10834
rect 18174 10782 18226 10834
rect 35870 10782 35922 10834
rect 38334 10782 38386 10834
rect 2494 10670 2546 10722
rect 4734 10670 4786 10722
rect 9662 10670 9714 10722
rect 10446 10670 10498 10722
rect 13806 10670 13858 10722
rect 17390 10670 17442 10722
rect 20190 10670 20242 10722
rect 22990 10670 23042 10722
rect 27246 10670 27298 10722
rect 30382 10670 30434 10722
rect 7758 10558 7810 10610
rect 8206 10558 8258 10610
rect 16158 10558 16210 10610
rect 16494 10558 16546 10610
rect 17614 10558 17666 10610
rect 33182 10558 33234 10610
rect 33630 10558 33682 10610
rect 36990 10558 37042 10610
rect 3390 10446 3442 10498
rect 11790 10446 11842 10498
rect 19406 10446 19458 10498
rect 21982 10446 22034 10498
rect 26238 10446 26290 10498
rect 29038 10446 29090 10498
rect 37550 10446 37602 10498
rect 13022 10334 13074 10386
rect 36654 10334 36706 10386
rect 5876 10166 5928 10218
rect 5980 10166 6032 10218
rect 6084 10166 6136 10218
rect 15200 10166 15252 10218
rect 15304 10166 15356 10218
rect 15408 10166 15460 10218
rect 24524 10166 24576 10218
rect 24628 10166 24680 10218
rect 24732 10166 24784 10218
rect 33848 10166 33900 10218
rect 33952 10166 34004 10218
rect 34056 10166 34108 10218
rect 37774 9998 37826 10050
rect 3502 9886 3554 9938
rect 9998 9886 10050 9938
rect 11454 9886 11506 9938
rect 15150 9886 15202 9938
rect 16942 9886 16994 9938
rect 17390 9886 17442 9938
rect 17838 9886 17890 9938
rect 19294 9886 19346 9938
rect 22430 9886 22482 9938
rect 27582 9886 27634 9938
rect 30942 9886 30994 9938
rect 33854 9886 33906 9938
rect 8542 9774 8594 9826
rect 8990 9774 9042 9826
rect 9886 9774 9938 9826
rect 35758 9774 35810 9826
rect 2382 9662 2434 9714
rect 6302 9662 6354 9714
rect 12798 9662 12850 9714
rect 14814 9662 14866 9714
rect 15710 9662 15762 9714
rect 20638 9662 20690 9714
rect 23550 9662 23602 9714
rect 26574 9662 26626 9714
rect 31950 9662 32002 9714
rect 34750 9662 34802 9714
rect 5518 9550 5570 9602
rect 32958 9550 33010 9602
rect 35534 9550 35586 9602
rect 36318 9550 36370 9602
rect 36990 9550 37042 9602
rect 10538 9382 10590 9434
rect 10642 9382 10694 9434
rect 10746 9382 10798 9434
rect 19862 9382 19914 9434
rect 19966 9382 20018 9434
rect 20070 9382 20122 9434
rect 29186 9382 29238 9434
rect 29290 9382 29342 9434
rect 29394 9382 29446 9434
rect 38510 9382 38562 9434
rect 38614 9382 38666 9434
rect 38718 9382 38770 9434
rect 6190 9214 6242 9266
rect 9662 9214 9714 9266
rect 14142 9214 14194 9266
rect 33966 9214 34018 9266
rect 37326 9214 37378 9266
rect 19406 9102 19458 9154
rect 29934 9102 29986 9154
rect 31166 9102 31218 9154
rect 31502 9102 31554 9154
rect 31838 9102 31890 9154
rect 32174 9102 32226 9154
rect 33294 9102 33346 9154
rect 33630 9102 33682 9154
rect 3054 8990 3106 9042
rect 3726 8990 3778 9042
rect 11230 8990 11282 9042
rect 11678 8990 11730 9042
rect 15038 8990 15090 9042
rect 30942 8990 30994 9042
rect 32398 8990 32450 9042
rect 34190 8990 34242 9042
rect 34750 8990 34802 9042
rect 7086 8878 7138 8930
rect 18398 8878 18450 8930
rect 28926 8878 28978 8930
rect 6750 8766 6802 8818
rect 14702 8766 14754 8818
rect 37886 8766 37938 8818
rect 5876 8598 5928 8650
rect 5980 8598 6032 8650
rect 6084 8598 6136 8650
rect 15200 8598 15252 8650
rect 15304 8598 15356 8650
rect 15408 8598 15460 8650
rect 24524 8598 24576 8650
rect 24628 8598 24680 8650
rect 24732 8598 24784 8650
rect 33848 8598 33900 8650
rect 33952 8598 34004 8650
rect 34056 8598 34108 8650
rect 3614 8318 3666 8370
rect 7310 8318 7362 8370
rect 11454 8318 11506 8370
rect 15934 8318 15986 8370
rect 18734 8318 18786 8370
rect 27582 8318 27634 8370
rect 31166 8318 31218 8370
rect 31390 8318 31442 8370
rect 34638 8318 34690 8370
rect 37774 8318 37826 8370
rect 21982 8206 22034 8258
rect 29822 8206 29874 8258
rect 4958 8094 5010 8146
rect 6078 8094 6130 8146
rect 12462 8094 12514 8146
rect 17166 8094 17218 8146
rect 19742 8094 19794 8146
rect 26574 8094 26626 8146
rect 32510 8094 32562 8146
rect 35646 8094 35698 8146
rect 22206 7982 22258 8034
rect 30046 7982 30098 8034
rect 36318 7982 36370 8034
rect 36990 7982 37042 8034
rect 10538 7814 10590 7866
rect 10642 7814 10694 7866
rect 10746 7814 10798 7866
rect 19862 7814 19914 7866
rect 19966 7814 20018 7866
rect 20070 7814 20122 7866
rect 29186 7814 29238 7866
rect 29290 7814 29342 7866
rect 29394 7814 29446 7866
rect 38510 7814 38562 7866
rect 38614 7814 38666 7866
rect 38718 7814 38770 7866
rect 4734 7646 4786 7698
rect 5630 7646 5682 7698
rect 33406 7646 33458 7698
rect 6862 7534 6914 7586
rect 11902 7534 11954 7586
rect 14366 7534 14418 7586
rect 27694 7534 27746 7586
rect 30494 7534 30546 7586
rect 36094 7534 36146 7586
rect 36654 7534 36706 7586
rect 38110 7534 38162 7586
rect 1822 7422 1874 7474
rect 2270 7422 2322 7474
rect 33070 7422 33122 7474
rect 36990 7422 37042 7474
rect 7870 7310 7922 7362
rect 10558 7310 10610 7362
rect 13358 7310 13410 7362
rect 28702 7310 28754 7362
rect 29262 7310 29314 7362
rect 29822 7310 29874 7362
rect 31502 7310 31554 7362
rect 34974 7310 35026 7362
rect 5294 7198 5346 7250
rect 29150 7198 29202 7250
rect 29822 7198 29874 7250
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 7646 6750 7698 6802
rect 10670 6750 10722 6802
rect 16830 6750 16882 6802
rect 32398 6750 32450 6802
rect 34190 6750 34242 6802
rect 27246 6638 27298 6690
rect 27694 6638 27746 6690
rect 30718 6638 30770 6690
rect 37774 6638 37826 6690
rect 6638 6526 6690 6578
rect 12014 6526 12066 6578
rect 15710 6526 15762 6578
rect 27918 6526 27970 6578
rect 28254 6526 28306 6578
rect 28590 6526 28642 6578
rect 29150 6526 29202 6578
rect 29486 6526 29538 6578
rect 30158 6526 30210 6578
rect 30494 6526 30546 6578
rect 31278 6526 31330 6578
rect 33182 6526 33234 6578
rect 34974 6526 35026 6578
rect 29822 6414 29874 6466
rect 36990 6414 37042 6466
rect 10538 6246 10590 6298
rect 10642 6246 10694 6298
rect 10746 6246 10798 6298
rect 19862 6246 19914 6298
rect 19966 6246 20018 6298
rect 20070 6246 20122 6298
rect 29186 6246 29238 6298
rect 29290 6246 29342 6298
rect 29394 6246 29446 6298
rect 38510 6246 38562 6298
rect 38614 6246 38666 6298
rect 38718 6246 38770 6298
rect 27694 6078 27746 6130
rect 33406 6078 33458 6130
rect 5742 5966 5794 6018
rect 6862 5966 6914 6018
rect 11790 5966 11842 6018
rect 26686 5966 26738 6018
rect 27022 5966 27074 6018
rect 28030 5966 28082 6018
rect 28366 5966 28418 6018
rect 29038 5966 29090 6018
rect 29374 5966 29426 6018
rect 30270 5966 30322 6018
rect 33070 5966 33122 6018
rect 37998 5966 38050 6018
rect 27470 5854 27522 5906
rect 28814 5854 28866 5906
rect 29710 5854 29762 5906
rect 33854 5854 33906 5906
rect 4734 5742 4786 5794
rect 7982 5742 8034 5794
rect 10558 5742 10610 5794
rect 26462 5742 26514 5794
rect 31390 5742 31442 5794
rect 31950 5742 32002 5794
rect 34414 5742 34466 5794
rect 36766 5742 36818 5794
rect 5876 5462 5928 5514
rect 5980 5462 6032 5514
rect 6084 5462 6136 5514
rect 15200 5462 15252 5514
rect 15304 5462 15356 5514
rect 15408 5462 15460 5514
rect 24524 5462 24576 5514
rect 24628 5462 24680 5514
rect 24732 5462 24784 5514
rect 33848 5462 33900 5514
rect 33952 5462 34004 5514
rect 34056 5462 34108 5514
rect 29710 5182 29762 5234
rect 30382 5182 30434 5234
rect 32398 5182 32450 5234
rect 35198 5182 35250 5234
rect 26798 5070 26850 5122
rect 30830 5070 30882 5122
rect 36990 5070 37042 5122
rect 27022 4958 27074 5010
rect 27358 4958 27410 5010
rect 27694 4958 27746 5010
rect 28030 4958 28082 5010
rect 31614 4958 31666 5010
rect 36094 4958 36146 5010
rect 28366 4846 28418 4898
rect 29262 4846 29314 4898
rect 37774 4846 37826 4898
rect 10538 4678 10590 4730
rect 10642 4678 10694 4730
rect 10746 4678 10798 4730
rect 19862 4678 19914 4730
rect 19966 4678 20018 4730
rect 20070 4678 20122 4730
rect 29186 4678 29238 4730
rect 29290 4678 29342 4730
rect 29394 4678 29446 4730
rect 38510 4678 38562 4730
rect 38614 4678 38666 4730
rect 38718 4678 38770 4730
rect 26686 4510 26738 4562
rect 27358 4510 27410 4562
rect 28702 4510 28754 4562
rect 29038 4510 29090 4562
rect 30494 4510 30546 4562
rect 32510 4510 32562 4562
rect 23102 4398 23154 4450
rect 26126 4398 26178 4450
rect 28030 4398 28082 4450
rect 28366 4398 28418 4450
rect 37774 4398 37826 4450
rect 26462 4286 26514 4338
rect 27134 4286 27186 4338
rect 27694 4286 27746 4338
rect 29374 4286 29426 4338
rect 29822 4286 29874 4338
rect 30942 4286 30994 4338
rect 33070 4286 33122 4338
rect 34638 4286 34690 4338
rect 32062 4174 32114 4226
rect 33518 4174 33570 4226
rect 35198 4174 35250 4226
rect 36766 4174 36818 4226
rect 5876 3894 5928 3946
rect 5980 3894 6032 3946
rect 6084 3894 6136 3946
rect 15200 3894 15252 3946
rect 15304 3894 15356 3946
rect 15408 3894 15460 3946
rect 24524 3894 24576 3946
rect 24628 3894 24680 3946
rect 24732 3894 24784 3946
rect 33848 3894 33900 3946
rect 33952 3894 34004 3946
rect 34056 3894 34108 3946
rect 22878 3614 22930 3666
rect 28926 3614 28978 3666
rect 29710 3614 29762 3666
rect 30494 3614 30546 3666
rect 34302 3614 34354 3666
rect 36430 3614 36482 3666
rect 22430 3502 22482 3554
rect 26910 3502 26962 3554
rect 27582 3502 27634 3554
rect 28590 3502 28642 3554
rect 30046 3502 30098 3554
rect 32174 3502 32226 3554
rect 35982 3502 36034 3554
rect 37326 3502 37378 3554
rect 21534 3390 21586 3442
rect 21758 3390 21810 3442
rect 22094 3390 22146 3442
rect 26126 3390 26178 3442
rect 27134 3390 27186 3442
rect 27806 3390 27858 3442
rect 32510 3390 32562 3442
rect 33070 3390 33122 3442
rect 37550 3390 37602 3442
rect 37886 3390 37938 3442
rect 24558 3278 24610 3330
rect 26462 3278 26514 3330
rect 10538 3110 10590 3162
rect 10642 3110 10694 3162
rect 10746 3110 10798 3162
rect 19862 3110 19914 3162
rect 19966 3110 20018 3162
rect 20070 3110 20122 3162
rect 29186 3110 29238 3162
rect 29290 3110 29342 3162
rect 29394 3110 29446 3162
rect 38510 3110 38562 3162
rect 38614 3110 38666 3162
rect 38718 3110 38770 3162
<< metal2 >>
rect 18144 39200 18256 40000
rect 18816 39200 18928 40000
rect 19488 39200 19600 40000
rect 20160 39200 20272 40000
rect 20832 39200 20944 40000
rect 21504 39200 21616 40000
rect 22176 39200 22288 40000
rect 22848 39200 22960 40000
rect 23520 39200 23632 40000
rect 24192 39200 24304 40000
rect 24864 39200 24976 40000
rect 25536 39200 25648 40000
rect 26208 39200 26320 40000
rect 26880 39200 26992 40000
rect 27552 39200 27664 40000
rect 28224 39200 28336 40000
rect 28896 39200 29008 40000
rect 29568 39200 29680 40000
rect 30240 39200 30352 40000
rect 30912 39200 31024 40000
rect 31584 39200 31696 40000
rect 32256 39200 32368 40000
rect 32928 39200 33040 40000
rect 33600 39200 33712 40000
rect 34272 39200 34384 40000
rect 34944 39200 35056 40000
rect 35196 39732 35252 39742
rect 5874 36876 6138 36886
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 5874 36810 6138 36820
rect 15198 36876 15462 36886
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15198 36810 15462 36820
rect 17724 36484 17780 36494
rect 18172 36484 18228 39200
rect 17724 36482 18228 36484
rect 17724 36430 17726 36482
rect 17778 36430 18228 36482
rect 17724 36428 18228 36430
rect 17724 36418 17780 36428
rect 17948 36260 18004 36270
rect 17948 36166 18004 36204
rect 10536 36092 10800 36102
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10536 36026 10800 36036
rect 18172 35922 18228 36428
rect 18396 36484 18452 36494
rect 18844 36484 18900 39200
rect 19516 36594 19572 39200
rect 20188 36708 20244 39200
rect 20860 37828 20916 39200
rect 20860 37772 21364 37828
rect 19516 36542 19518 36594
rect 19570 36542 19572 36594
rect 19516 36530 19572 36542
rect 19740 36652 20244 36708
rect 18396 36482 18900 36484
rect 18396 36430 18398 36482
rect 18450 36430 18900 36482
rect 18396 36428 18900 36430
rect 18396 36418 18452 36428
rect 18172 35870 18174 35922
rect 18226 35870 18228 35922
rect 18172 35858 18228 35870
rect 18620 36258 18676 36270
rect 18620 36206 18622 36258
rect 18674 36206 18676 36258
rect 18620 35812 18676 36206
rect 18844 35922 18900 36428
rect 18844 35870 18846 35922
rect 18898 35870 18900 35922
rect 18844 35858 18900 35870
rect 19740 35812 19796 36652
rect 21308 36594 21364 37772
rect 21532 36932 21588 39200
rect 22204 37266 22260 39200
rect 22204 37214 22206 37266
rect 22258 37214 22260 37266
rect 22204 37202 22260 37214
rect 21532 36866 21588 36876
rect 22540 36932 22596 36942
rect 21308 36542 21310 36594
rect 21362 36542 21364 36594
rect 21308 36530 21364 36542
rect 20188 36484 20244 36494
rect 20188 36482 20580 36484
rect 20188 36430 20190 36482
rect 20242 36430 20580 36482
rect 20188 36428 20580 36430
rect 20188 36418 20244 36428
rect 19860 36092 20124 36102
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 19860 36026 20124 36036
rect 20188 35924 20244 35934
rect 20188 35830 20244 35868
rect 20524 35922 20580 36428
rect 22204 36482 22260 36494
rect 22204 36430 22206 36482
rect 22258 36430 22260 36482
rect 20524 35870 20526 35922
rect 20578 35870 20580 35922
rect 20524 35858 20580 35870
rect 20748 36260 20804 36270
rect 19852 35812 19908 35822
rect 19740 35810 20132 35812
rect 19740 35758 19854 35810
rect 19906 35758 20132 35810
rect 19740 35756 20132 35758
rect 18620 35746 18676 35756
rect 19852 35746 19908 35756
rect 20076 35476 20132 35756
rect 20748 35698 20804 36204
rect 21532 36260 21588 36270
rect 21084 35924 21140 35934
rect 21140 35868 21252 35924
rect 21084 35858 21140 35868
rect 21196 35810 21252 35868
rect 21532 35922 21588 36204
rect 21532 35870 21534 35922
rect 21586 35870 21588 35922
rect 21532 35858 21588 35870
rect 22204 35922 22260 36430
rect 22204 35870 22206 35922
rect 22258 35870 22260 35922
rect 22204 35858 22260 35870
rect 22540 35922 22596 36876
rect 22652 36260 22708 36270
rect 22652 36166 22708 36204
rect 22540 35870 22542 35922
rect 22594 35870 22596 35922
rect 22540 35858 22596 35870
rect 21196 35758 21198 35810
rect 21250 35758 21252 35810
rect 21196 35746 21252 35758
rect 21868 35812 21924 35822
rect 21868 35718 21924 35756
rect 22876 35812 22932 39200
rect 23100 37266 23156 37278
rect 23100 37214 23102 37266
rect 23154 37214 23156 37266
rect 23100 36594 23156 37214
rect 23100 36542 23102 36594
rect 23154 36542 23156 36594
rect 23100 36530 23156 36542
rect 23100 35812 23156 35822
rect 22876 35810 23156 35812
rect 22876 35758 23102 35810
rect 23154 35758 23156 35810
rect 22876 35756 23156 35758
rect 20748 35646 20750 35698
rect 20802 35646 20804 35698
rect 20748 35634 20804 35646
rect 20076 35420 20468 35476
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 20412 35026 20468 35420
rect 20412 34974 20414 35026
rect 20466 34974 20468 35026
rect 20412 34962 20468 34974
rect 22876 35026 22932 35756
rect 23100 35746 23156 35756
rect 23436 35810 23492 35822
rect 23436 35758 23438 35810
rect 23490 35758 23492 35810
rect 22876 34974 22878 35026
rect 22930 34974 22932 35026
rect 22876 34962 22932 34974
rect 23436 34916 23492 35758
rect 23548 35812 23604 39200
rect 23772 35812 23828 35822
rect 23548 35810 23828 35812
rect 23548 35758 23774 35810
rect 23826 35758 23828 35810
rect 23548 35756 23828 35758
rect 23548 35026 23604 35756
rect 23772 35746 23828 35756
rect 24108 35812 24164 35822
rect 24108 35718 24164 35756
rect 23548 34974 23550 35026
rect 23602 34974 23604 35026
rect 23548 34962 23604 34974
rect 24220 35028 24276 39200
rect 24522 36876 24786 36886
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24522 36810 24786 36820
rect 24892 36708 24948 39200
rect 25564 37380 25620 39200
rect 26236 37828 26292 39200
rect 26236 37772 26740 37828
rect 25564 37324 26068 37380
rect 24892 36642 24948 36652
rect 25676 36482 25732 36494
rect 25676 36430 25678 36482
rect 25730 36430 25732 36482
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 24220 35026 24500 35028
rect 24220 34974 24222 35026
rect 24274 34974 24500 35026
rect 24220 34972 24500 34974
rect 24220 34962 24276 34972
rect 23436 34850 23492 34860
rect 24444 34914 24500 34972
rect 24444 34862 24446 34914
rect 24498 34862 24500 34914
rect 24444 34850 24500 34862
rect 25340 34916 25396 34926
rect 25340 34822 25396 34860
rect 24780 34804 24836 34814
rect 24780 34710 24836 34748
rect 25676 34802 25732 36430
rect 26012 35586 26068 37324
rect 26124 36708 26180 36718
rect 26124 36594 26180 36652
rect 26124 36542 26126 36594
rect 26178 36542 26180 36594
rect 26124 36530 26180 36542
rect 26684 36370 26740 37772
rect 26908 37380 26964 39200
rect 26908 37324 27412 37380
rect 26684 36318 26686 36370
rect 26738 36318 26740 36370
rect 26684 36306 26740 36318
rect 27132 36372 27188 36382
rect 27132 36278 27188 36316
rect 27356 36036 27412 37324
rect 27580 36708 27636 39200
rect 28252 36820 28308 39200
rect 28924 37828 28980 39200
rect 28924 37772 29428 37828
rect 28252 36764 28756 36820
rect 27580 36642 27636 36652
rect 27468 36260 27524 36270
rect 28364 36260 28420 36270
rect 27468 36258 28420 36260
rect 27468 36206 27470 36258
rect 27522 36206 28366 36258
rect 28418 36206 28420 36258
rect 27468 36204 28420 36206
rect 27468 36194 27524 36204
rect 28364 36194 28420 36204
rect 27356 35980 27860 36036
rect 26012 35534 26014 35586
rect 26066 35534 26068 35586
rect 26012 35522 26068 35534
rect 26124 35812 26180 35822
rect 26124 34914 26180 35756
rect 26796 35700 26852 35710
rect 27356 35700 27412 35710
rect 26124 34862 26126 34914
rect 26178 34862 26180 34914
rect 26124 34850 26180 34862
rect 26348 35698 26852 35700
rect 26348 35646 26798 35698
rect 26850 35646 26852 35698
rect 26348 35644 26852 35646
rect 25676 34750 25678 34802
rect 25730 34750 25732 34802
rect 25676 34738 25732 34750
rect 26348 34802 26404 35644
rect 26796 35634 26852 35644
rect 27020 35698 27412 35700
rect 27020 35646 27358 35698
rect 27410 35646 27412 35698
rect 27020 35644 27412 35646
rect 26348 34750 26350 34802
rect 26402 34750 26404 34802
rect 26348 34738 26404 34750
rect 26684 34804 26740 34814
rect 26684 34710 26740 34748
rect 27020 34802 27076 35644
rect 27356 35634 27412 35644
rect 27804 35586 27860 35980
rect 28700 35922 28756 36764
rect 28812 36708 28868 36718
rect 28812 36594 28868 36652
rect 29372 36706 29428 37772
rect 29372 36654 29374 36706
rect 29426 36654 29428 36706
rect 29372 36642 29428 36654
rect 28812 36542 28814 36594
rect 28866 36542 28868 36594
rect 28812 36530 28868 36542
rect 28700 35870 28702 35922
rect 28754 35870 28756 35922
rect 28700 35700 28756 35870
rect 28924 36372 28980 36382
rect 28924 35922 28980 36316
rect 29184 36092 29448 36102
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29184 36026 29448 36036
rect 28924 35870 28926 35922
rect 28978 35870 28980 35922
rect 28924 35858 28980 35870
rect 29596 35924 29652 39200
rect 29708 36708 29764 36718
rect 29708 36706 29988 36708
rect 29708 36654 29710 36706
rect 29762 36654 29988 36706
rect 29708 36652 29988 36654
rect 29708 36642 29764 36652
rect 29708 36484 29764 36494
rect 29708 36390 29764 36428
rect 29932 36370 29988 36652
rect 30268 36484 30324 39200
rect 30940 36708 30996 39200
rect 30940 36642 30996 36652
rect 30268 36418 30324 36428
rect 30716 36484 30772 36522
rect 30716 36418 30772 36428
rect 29932 36318 29934 36370
rect 29986 36318 29988 36370
rect 29932 36306 29988 36318
rect 31612 36370 31668 39200
rect 32284 36596 32340 39200
rect 32956 36932 33012 39200
rect 33628 37828 33684 39200
rect 33628 37772 34244 37828
rect 32956 36866 33012 36876
rect 33628 36932 33684 36942
rect 32284 36530 32340 36540
rect 32620 36708 32676 36718
rect 32620 36594 32676 36652
rect 32620 36542 32622 36594
rect 32674 36542 32676 36594
rect 32620 36530 32676 36542
rect 31612 36318 31614 36370
rect 31666 36318 31668 36370
rect 31612 36306 31668 36318
rect 30492 36258 30548 36270
rect 30492 36206 30494 36258
rect 30546 36206 30548 36258
rect 29820 35924 29876 35934
rect 29596 35922 29876 35924
rect 29596 35870 29822 35922
rect 29874 35870 29876 35922
rect 29596 35868 29876 35870
rect 29820 35858 29876 35868
rect 29148 35700 29204 35710
rect 28700 35698 29204 35700
rect 28700 35646 29150 35698
rect 29202 35646 29204 35698
rect 28700 35644 29204 35646
rect 29148 35634 29204 35644
rect 30492 35698 30548 36206
rect 30716 36260 30772 36270
rect 30716 35922 30772 36204
rect 32172 36260 32228 36270
rect 32172 36166 32228 36204
rect 30716 35870 30718 35922
rect 30770 35870 30772 35922
rect 30716 35858 30772 35870
rect 31948 35924 32004 35934
rect 31948 35830 32004 35868
rect 32396 35812 32452 35822
rect 30492 35646 30494 35698
rect 30546 35646 30548 35698
rect 30492 35634 30548 35646
rect 31612 35698 31668 35710
rect 31612 35646 31614 35698
rect 31666 35646 31668 35698
rect 27804 35534 27806 35586
rect 27858 35534 27860 35586
rect 27804 35522 27860 35534
rect 27020 34750 27022 34802
rect 27074 34750 27076 34802
rect 27020 34738 27076 34750
rect 10536 34524 10800 34534
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10536 34458 10800 34468
rect 19860 34524 20124 34534
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 19860 34458 20124 34468
rect 29184 34524 29448 34534
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29184 34458 29448 34468
rect 5874 33740 6138 33750
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 5874 33674 6138 33684
rect 15198 33740 15462 33750
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15198 33674 15462 33684
rect 24522 33740 24786 33750
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24522 33674 24786 33684
rect 10536 32956 10800 32966
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10536 32890 10800 32900
rect 19860 32956 20124 32966
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 19860 32890 20124 32900
rect 29184 32956 29448 32966
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29184 32890 29448 32900
rect 5874 32172 6138 32182
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 5874 32106 6138 32116
rect 15198 32172 15462 32182
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15198 32106 15462 32116
rect 24522 32172 24786 32182
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24522 32106 24786 32116
rect 10536 31388 10800 31398
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10536 31322 10800 31332
rect 19860 31388 20124 31398
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 19860 31322 20124 31332
rect 29184 31388 29448 31398
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29184 31322 29448 31332
rect 31612 31220 31668 35646
rect 32396 34914 32452 35756
rect 33180 35700 33236 35710
rect 32396 34862 32398 34914
rect 32450 34862 32452 34914
rect 32396 34850 32452 34862
rect 32620 35698 33236 35700
rect 32620 35646 33182 35698
rect 33234 35646 33236 35698
rect 32620 35644 33236 35646
rect 32620 34802 32676 35644
rect 33180 35634 33236 35644
rect 33628 35586 33684 36876
rect 33846 36876 34110 36886
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 33846 36810 34110 36820
rect 34188 36372 34244 37772
rect 34188 36306 34244 36316
rect 33740 36258 33796 36270
rect 33740 36206 33742 36258
rect 33794 36206 33796 36258
rect 33740 35924 33796 36206
rect 33740 35858 33796 35868
rect 33628 35534 33630 35586
rect 33682 35534 33684 35586
rect 33628 35522 33684 35534
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 34300 35140 34356 39200
rect 34972 36820 35028 39200
rect 35196 37268 35252 39676
rect 35616 39200 35728 40000
rect 36288 39200 36400 40000
rect 36960 39200 37072 40000
rect 37632 39200 37744 40000
rect 34636 36764 35028 36820
rect 35084 37212 35252 37268
rect 34412 36596 34468 36606
rect 34412 36502 34468 36540
rect 34524 35700 34580 35710
rect 34524 35606 34580 35644
rect 33964 35084 34356 35140
rect 32620 34750 32622 34802
rect 32674 34750 32676 34802
rect 32620 34738 32676 34750
rect 33516 34804 33572 34814
rect 33516 34710 33572 34748
rect 33964 34802 34020 35084
rect 34636 35028 34692 36764
rect 35084 36036 35140 37212
rect 35308 36372 35364 36382
rect 35308 36278 35364 36316
rect 35084 35980 35252 36036
rect 34748 35812 34804 35822
rect 34748 35718 34804 35756
rect 35084 35812 35140 35822
rect 35084 35718 35140 35756
rect 33964 34750 33966 34802
rect 34018 34750 34020 34802
rect 33964 34738 34020 34750
rect 34076 34972 34692 35028
rect 34748 35364 34804 35374
rect 34076 34580 34132 34972
rect 34300 34804 34356 34814
rect 34300 34802 34580 34804
rect 34300 34750 34302 34802
rect 34354 34750 34580 34802
rect 34300 34748 34580 34750
rect 34300 34738 34356 34748
rect 33628 34524 34132 34580
rect 33628 34354 33684 34524
rect 33628 34302 33630 34354
rect 33682 34302 33684 34354
rect 33628 34290 33684 34302
rect 34076 34244 34132 34254
rect 34076 34150 34132 34188
rect 34412 34130 34468 34142
rect 34412 34078 34414 34130
rect 34466 34078 34468 34130
rect 33846 33740 34110 33750
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 33846 33674 34110 33684
rect 31612 31154 31668 31164
rect 32620 33236 32676 33246
rect 5874 30604 6138 30614
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 5874 30538 6138 30548
rect 15198 30604 15462 30614
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15198 30538 15462 30548
rect 24522 30604 24786 30614
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24522 30538 24786 30548
rect 10444 30322 10500 30334
rect 10444 30270 10446 30322
rect 10498 30270 10500 30322
rect 9436 29988 9492 29998
rect 5874 29036 6138 29046
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 5874 28970 6138 28980
rect 8652 28756 8708 28766
rect 5516 27972 5572 27982
rect 2380 26402 2436 26414
rect 2380 26350 2382 26402
rect 2434 26350 2436 26402
rect 1596 26066 1652 26078
rect 1596 26014 1598 26066
rect 1650 26014 1652 26066
rect 1484 25396 1540 25406
rect 1484 21812 1540 25340
rect 1596 24836 1652 26014
rect 2156 25396 2212 25406
rect 2156 25302 2212 25340
rect 1596 24770 1652 24780
rect 2268 24836 2324 24846
rect 2268 24742 2324 24780
rect 2268 24052 2324 24062
rect 2380 24052 2436 26350
rect 4284 26292 4340 26302
rect 3500 25620 3556 25630
rect 3500 25526 3556 25564
rect 4060 24724 4116 24734
rect 2268 24050 2436 24052
rect 2268 23998 2270 24050
rect 2322 23998 2436 24050
rect 2268 23996 2436 23998
rect 3500 24610 3556 24622
rect 3500 24558 3502 24610
rect 3554 24558 3556 24610
rect 2268 23986 2324 23996
rect 1932 23828 1988 23838
rect 1932 22482 1988 23772
rect 2940 23826 2996 23838
rect 2940 23774 2942 23826
rect 2994 23774 2996 23826
rect 2940 23378 2996 23774
rect 3500 23492 3556 24558
rect 4060 24050 4116 24668
rect 4060 23998 4062 24050
rect 4114 23998 4116 24050
rect 4060 23986 4116 23998
rect 3500 23426 3556 23436
rect 3724 23716 3780 23726
rect 2940 23326 2942 23378
rect 2994 23326 2996 23378
rect 2940 23314 2996 23326
rect 3724 23378 3780 23660
rect 3724 23326 3726 23378
rect 3778 23326 3780 23378
rect 3724 23314 3780 23326
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 22418 1988 22430
rect 4060 22484 4116 22494
rect 4060 22390 4116 22428
rect 2268 22258 2324 22270
rect 2268 22206 2270 22258
rect 2322 22206 2324 22258
rect 1596 21812 1652 21822
rect 1484 21810 1652 21812
rect 1484 21758 1598 21810
rect 1650 21758 1652 21810
rect 1484 21756 1652 21758
rect 1596 21746 1652 21756
rect 2268 21810 2324 22206
rect 2268 21758 2270 21810
rect 2322 21758 2324 21810
rect 2268 21746 2324 21758
rect 3052 22258 3108 22270
rect 3052 22206 3054 22258
rect 3106 22206 3108 22258
rect 3052 21700 3108 22206
rect 3052 21634 3108 21644
rect 4172 21588 4228 21598
rect 3948 21476 4004 21486
rect 3052 20916 3108 20926
rect 3836 20916 3892 20926
rect 3052 20690 3108 20860
rect 3052 20638 3054 20690
rect 3106 20638 3108 20690
rect 3052 20626 3108 20638
rect 3724 20914 3892 20916
rect 3724 20862 3838 20914
rect 3890 20862 3892 20914
rect 3724 20860 3892 20862
rect 3612 20020 3668 20030
rect 3612 19926 3668 19964
rect 3052 19796 3108 19806
rect 3052 19122 3108 19740
rect 3052 19070 3054 19122
rect 3106 19070 3108 19122
rect 3052 19058 3108 19070
rect 2380 19012 2436 19022
rect 1820 17442 1876 17454
rect 1820 17390 1822 17442
rect 1874 17390 1876 17442
rect 1708 15988 1764 15998
rect 1820 15988 1876 17390
rect 2156 16884 2212 16894
rect 2156 16790 2212 16828
rect 1708 15986 1876 15988
rect 1708 15934 1710 15986
rect 1762 15934 1876 15986
rect 1708 15932 1876 15934
rect 1596 15090 1652 15102
rect 1596 15038 1598 15090
rect 1650 15038 1652 15090
rect 1596 11732 1652 15038
rect 1708 14868 1764 15932
rect 2044 15876 2100 15886
rect 2044 15874 2212 15876
rect 2044 15822 2046 15874
rect 2098 15822 2212 15874
rect 2044 15820 2212 15822
rect 2044 15810 2100 15820
rect 1708 14802 1764 14812
rect 1932 14418 1988 14430
rect 1932 14366 1934 14418
rect 1986 14366 1988 14418
rect 1596 11666 1652 11676
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 12178 1876 13694
rect 1932 13524 1988 14366
rect 1932 13074 1988 13468
rect 2044 14306 2100 14318
rect 2044 14254 2046 14306
rect 2098 14254 2100 14306
rect 2044 13300 2100 14254
rect 2044 13234 2100 13244
rect 1932 13022 1934 13074
rect 1986 13022 1988 13074
rect 1932 13010 1988 13022
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 8428 1876 12126
rect 2156 12178 2212 15820
rect 2380 15538 2436 18956
rect 3724 18676 3780 20860
rect 3836 20850 3892 20860
rect 3948 20188 4004 21420
rect 3836 20132 4004 20188
rect 4060 21364 4116 21374
rect 3836 20130 3892 20132
rect 3836 20078 3838 20130
rect 3890 20078 3892 20130
rect 3836 20066 3892 20078
rect 4060 19346 4116 21308
rect 4172 20018 4228 21532
rect 4284 21028 4340 26236
rect 4620 26290 4676 26302
rect 4620 26238 4622 26290
rect 4674 26238 4676 26290
rect 4620 25620 4676 26238
rect 5292 26292 5348 26302
rect 5292 26198 5348 26236
rect 5516 25730 5572 27916
rect 7980 27972 8036 27982
rect 7980 27878 8036 27916
rect 6972 27746 7028 27758
rect 6972 27694 6974 27746
rect 7026 27694 7028 27746
rect 5874 27468 6138 27478
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 5874 27402 6138 27412
rect 6076 26964 6132 26974
rect 5516 25678 5518 25730
rect 5570 25678 5572 25730
rect 5516 25666 5572 25678
rect 5628 26292 5684 26302
rect 4620 25554 4676 25564
rect 5180 25284 5236 25294
rect 4956 25228 5180 25284
rect 4956 24722 5012 25228
rect 5180 25218 5236 25228
rect 5628 25284 5684 26236
rect 6076 26290 6132 26908
rect 6972 26964 7028 27694
rect 8316 27748 8372 27758
rect 6972 26898 7028 26908
rect 7084 27186 7140 27198
rect 7084 27134 7086 27186
rect 7138 27134 7140 27186
rect 6076 26238 6078 26290
rect 6130 26238 6132 26290
rect 6076 26226 6132 26238
rect 5874 25900 6138 25910
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 5874 25834 6138 25844
rect 6300 25396 6356 25406
rect 6300 25302 6356 25340
rect 5628 25218 5684 25228
rect 4956 24670 4958 24722
rect 5010 24670 5012 24722
rect 4732 23380 4788 23390
rect 4732 21586 4788 23324
rect 4732 21534 4734 21586
rect 4786 21534 4788 21586
rect 4732 21522 4788 21534
rect 4956 23156 5012 24670
rect 5292 24724 5348 24734
rect 5292 24630 5348 24668
rect 5874 24332 6138 24342
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 5874 24266 6138 24276
rect 5740 23828 5796 23838
rect 5740 23734 5796 23772
rect 6300 23828 6356 23838
rect 6636 23828 6692 23838
rect 6356 23772 6580 23828
rect 6300 23762 6356 23772
rect 5852 23716 5908 23726
rect 5852 23622 5908 23660
rect 4956 21588 5012 23100
rect 5964 23492 6020 23502
rect 5964 23154 6020 23436
rect 6524 23380 6580 23772
rect 6636 23734 6692 23772
rect 7084 23492 7140 27134
rect 8092 26962 8148 26974
rect 8092 26910 8094 26962
rect 8146 26910 8148 26962
rect 8092 25508 8148 26910
rect 8316 26514 8372 27692
rect 8316 26462 8318 26514
rect 8370 26462 8372 26514
rect 8316 26450 8372 26462
rect 8428 26516 8484 26526
rect 8092 25442 8148 25452
rect 7868 24946 7924 24958
rect 7868 24894 7870 24946
rect 7922 24894 7924 24946
rect 7084 23426 7140 23436
rect 7644 24050 7700 24062
rect 7644 23998 7646 24050
rect 7698 23998 7700 24050
rect 6524 23324 6916 23380
rect 6860 23268 6916 23324
rect 7532 23268 7588 23278
rect 6860 23266 7588 23268
rect 6860 23214 6862 23266
rect 6914 23214 7534 23266
rect 7586 23214 7588 23266
rect 6860 23212 7588 23214
rect 6860 23202 6916 23212
rect 5964 23102 5966 23154
rect 6018 23102 6020 23154
rect 5964 23090 6020 23102
rect 6412 23156 6468 23166
rect 6412 23062 6468 23100
rect 5874 22764 6138 22774
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 5874 22698 6138 22708
rect 5516 22148 5572 22158
rect 5516 22146 5796 22148
rect 5516 22094 5518 22146
rect 5570 22094 5796 22146
rect 5516 22092 5796 22094
rect 5516 22082 5572 22092
rect 5068 21588 5124 21598
rect 5404 21588 5460 21598
rect 4956 21586 5404 21588
rect 4956 21534 5070 21586
rect 5122 21534 5404 21586
rect 4956 21532 5404 21534
rect 5068 21522 5124 21532
rect 5404 21494 5460 21532
rect 4284 20962 4340 20972
rect 5628 20690 5684 20702
rect 5628 20638 5630 20690
rect 5682 20638 5684 20690
rect 5628 20132 5684 20638
rect 5740 20188 5796 22092
rect 6076 22146 6132 22158
rect 6076 22094 6078 22146
rect 6130 22094 6132 22146
rect 5964 21586 6020 21598
rect 5964 21534 5966 21586
rect 6018 21534 6020 21586
rect 5964 21364 6020 21534
rect 6076 21476 6132 22094
rect 6076 21410 6132 21420
rect 5964 21298 6020 21308
rect 5874 21196 6138 21206
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 6972 21026 7028 23212
rect 7532 23202 7588 23212
rect 6972 20974 6974 21026
rect 7026 20974 7028 21026
rect 5964 20804 6020 20814
rect 5740 20132 5908 20188
rect 4956 20076 5684 20132
rect 4172 19966 4174 20018
rect 4226 19966 4228 20018
rect 4172 19954 4228 19966
rect 4732 20018 4788 20030
rect 4732 19966 4734 20018
rect 4786 19966 4788 20018
rect 4060 19294 4062 19346
rect 4114 19294 4116 19346
rect 4060 19282 4116 19294
rect 3724 18610 3780 18620
rect 3052 18562 3108 18574
rect 3052 18510 3054 18562
rect 3106 18510 3108 18562
rect 3052 18340 3108 18510
rect 3052 18274 3108 18284
rect 3948 18452 4004 18462
rect 3948 17778 4004 18396
rect 4060 18338 4116 18350
rect 4060 18286 4062 18338
rect 4114 18286 4116 18338
rect 4060 18228 4116 18286
rect 4060 18162 4116 18172
rect 3948 17726 3950 17778
rect 4002 17726 4004 17778
rect 3948 17714 4004 17726
rect 3052 17556 3108 17566
rect 3052 17462 3108 17500
rect 2604 16996 2660 17006
rect 2604 16882 2660 16940
rect 2604 16830 2606 16882
rect 2658 16830 2660 16882
rect 2604 16818 2660 16830
rect 3500 16996 3556 17006
rect 3052 16772 3108 16782
rect 2380 15486 2382 15538
rect 2434 15486 2436 15538
rect 2380 15474 2436 15486
rect 2940 16660 2996 16670
rect 2268 14644 2324 14654
rect 2268 13746 2324 14588
rect 2268 13694 2270 13746
rect 2322 13694 2324 13746
rect 2268 13682 2324 13694
rect 2156 12126 2158 12178
rect 2210 12126 2212 12178
rect 2156 12114 2212 12126
rect 2268 12850 2324 12862
rect 2268 12798 2270 12850
rect 2322 12798 2324 12850
rect 2268 11172 2324 12798
rect 2268 11106 2324 11116
rect 2380 11732 2436 11742
rect 2380 9714 2436 11676
rect 2940 11282 2996 16604
rect 3052 15986 3108 16716
rect 3052 15934 3054 15986
rect 3106 15934 3108 15986
rect 3052 15922 3108 15934
rect 2940 11230 2942 11282
rect 2994 11230 2996 11282
rect 2940 11218 2996 11230
rect 3388 11956 3444 11966
rect 2492 10724 2548 10734
rect 2492 10630 2548 10668
rect 3388 10498 3444 11900
rect 3388 10446 3390 10498
rect 3442 10446 3444 10498
rect 3388 10434 3444 10446
rect 3500 9938 3556 16940
rect 4060 16210 4116 16222
rect 4060 16158 4062 16210
rect 4114 16158 4116 16210
rect 4060 16100 4116 16158
rect 4732 16212 4788 19966
rect 4956 17106 5012 20076
rect 5852 19908 5908 20132
rect 5404 19852 5908 19908
rect 5964 20020 6020 20748
rect 6972 20804 7028 20974
rect 6972 20738 7028 20748
rect 7084 23042 7140 23054
rect 7084 22990 7086 23042
rect 7138 22990 7140 23042
rect 7084 20242 7140 22990
rect 7644 22596 7700 23998
rect 7868 23266 7924 24894
rect 8428 24946 8484 26460
rect 8652 25506 8708 28700
rect 8652 25454 8654 25506
rect 8706 25454 8708 25506
rect 8652 25442 8708 25454
rect 8988 27074 9044 27086
rect 8988 27022 8990 27074
rect 9042 27022 9044 27074
rect 8988 25508 9044 27022
rect 9436 27074 9492 29932
rect 10444 29988 10500 30270
rect 14476 30322 14532 30334
rect 14476 30270 14478 30322
rect 14530 30270 14532 30322
rect 10444 29922 10500 29932
rect 11452 30098 11508 30110
rect 11452 30046 11454 30098
rect 11506 30046 11508 30098
rect 10536 29820 10800 29830
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10536 29754 10800 29764
rect 9660 28756 9716 28766
rect 9660 28662 9716 28700
rect 10892 28530 10948 28542
rect 10892 28478 10894 28530
rect 10946 28478 10948 28530
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 10668 27748 10724 27758
rect 10668 27654 10724 27692
rect 9436 27022 9438 27074
rect 9490 27022 9492 27074
rect 9436 27010 9492 27022
rect 9996 27412 10052 27422
rect 9100 26852 9156 26862
rect 9100 26514 9156 26796
rect 9100 26462 9102 26514
rect 9154 26462 9156 26514
rect 9100 26450 9156 26462
rect 9772 26404 9828 26414
rect 9436 26402 9828 26404
rect 9436 26350 9774 26402
rect 9826 26350 9828 26402
rect 9436 26348 9828 26350
rect 9324 25508 9380 25518
rect 8988 25506 9380 25508
rect 8988 25454 8990 25506
rect 9042 25454 9326 25506
rect 9378 25454 9380 25506
rect 8988 25452 9380 25454
rect 8428 24894 8430 24946
rect 8482 24894 8484 24946
rect 8428 24882 8484 24894
rect 8988 25284 9044 25452
rect 9324 25442 9380 25452
rect 7868 23214 7870 23266
rect 7922 23214 7924 23266
rect 7868 23202 7924 23214
rect 7644 22530 7700 22540
rect 8428 22484 8484 22494
rect 7756 21588 7812 21598
rect 7756 20802 7812 21532
rect 7756 20750 7758 20802
rect 7810 20750 7812 20802
rect 7756 20738 7812 20750
rect 8092 20804 8148 20814
rect 7084 20190 7086 20242
rect 7138 20190 7140 20242
rect 7084 20178 7140 20190
rect 7532 20690 7588 20702
rect 7532 20638 7534 20690
rect 7586 20638 7588 20690
rect 7532 20244 7588 20638
rect 7532 20178 7588 20188
rect 4956 17054 4958 17106
rect 5010 17054 5012 17106
rect 4956 17042 5012 17054
rect 5292 18450 5348 18462
rect 5292 18398 5294 18450
rect 5346 18398 5348 18450
rect 5068 16884 5124 16894
rect 5292 16884 5348 18398
rect 5124 16828 5348 16884
rect 4732 16156 4900 16212
rect 4060 16034 4116 16044
rect 4732 15988 4788 15998
rect 4620 15316 4676 15326
rect 3836 15314 4676 15316
rect 3836 15262 4622 15314
rect 4674 15262 4676 15314
rect 3836 15260 4676 15262
rect 3612 14644 3668 14654
rect 3612 14550 3668 14588
rect 3836 13074 3892 15260
rect 4620 15250 4676 15260
rect 4732 13970 4788 15932
rect 4732 13918 4734 13970
rect 4786 13918 4788 13970
rect 4732 13906 4788 13918
rect 4844 13524 4900 16156
rect 5068 15876 5124 16828
rect 5404 16100 5460 19852
rect 5964 19796 6020 19964
rect 8092 20018 8148 20748
rect 8428 20802 8484 22428
rect 8652 22370 8708 22382
rect 8652 22318 8654 22370
rect 8706 22318 8708 22370
rect 8540 21812 8596 21822
rect 8540 21718 8596 21756
rect 8428 20750 8430 20802
rect 8482 20750 8484 20802
rect 8428 20738 8484 20750
rect 8092 19966 8094 20018
rect 8146 19966 8148 20018
rect 8092 19954 8148 19966
rect 8316 19906 8372 19918
rect 8316 19854 8318 19906
rect 8370 19854 8372 19906
rect 5740 19740 6020 19796
rect 7756 19796 7812 19806
rect 5740 19236 5796 19740
rect 7756 19702 7812 19740
rect 5874 19628 6138 19638
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 5874 19562 6138 19572
rect 5852 19236 5908 19246
rect 5740 19234 5908 19236
rect 5740 19182 5854 19234
rect 5906 19182 5908 19234
rect 5740 19180 5908 19182
rect 5852 19170 5908 19180
rect 5852 19012 5908 19022
rect 6972 19012 7028 19022
rect 5852 18918 5908 18956
rect 6860 19010 7028 19012
rect 6860 18958 6974 19010
rect 7026 18958 7028 19010
rect 6860 18956 7028 18958
rect 5852 18452 5908 18462
rect 5852 18358 5908 18396
rect 5874 18060 6138 18070
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 5874 17994 6138 18004
rect 5516 17556 5572 17566
rect 5516 17462 5572 17500
rect 6188 17442 6244 17454
rect 6188 17390 6190 17442
rect 6242 17390 6244 17442
rect 6188 16994 6244 17390
rect 6188 16942 6190 16994
rect 6242 16942 6244 16994
rect 6188 16930 6244 16942
rect 5964 16884 6020 16894
rect 5740 16828 5964 16884
rect 5628 16660 5684 16670
rect 5628 16566 5684 16604
rect 5068 15782 5124 15820
rect 5180 16044 5460 16100
rect 5740 16100 5796 16828
rect 5964 16790 6020 16828
rect 6860 16772 6916 18956
rect 6972 18946 7028 18956
rect 7756 19010 7812 19022
rect 7756 18958 7758 19010
rect 7810 18958 7812 19010
rect 7756 18452 7812 18958
rect 8316 18674 8372 19854
rect 8316 18622 8318 18674
rect 8370 18622 8372 18674
rect 8316 18610 8372 18622
rect 7756 18386 7812 18396
rect 8652 18228 8708 22318
rect 8988 22372 9044 25228
rect 9436 25060 9492 26348
rect 9772 26338 9828 26348
rect 9100 25004 9492 25060
rect 9548 25508 9604 25518
rect 9100 24162 9156 25004
rect 9100 24110 9102 24162
rect 9154 24110 9156 24162
rect 9100 24098 9156 24110
rect 9548 23828 9604 25452
rect 9996 25506 10052 27356
rect 10536 26684 10800 26694
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10536 26618 10800 26628
rect 10892 26516 10948 28478
rect 10892 26450 10948 26460
rect 11004 27746 11060 27758
rect 11004 27694 11006 27746
rect 11058 27694 11060 27746
rect 9996 25454 9998 25506
rect 10050 25454 10052 25506
rect 9996 25442 10052 25454
rect 10108 25396 10164 25406
rect 10108 24834 10164 25340
rect 10536 25116 10800 25126
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10536 25050 10800 25060
rect 11004 25060 11060 27694
rect 11452 26964 11508 30046
rect 12460 29540 12516 29550
rect 12348 29314 12404 29326
rect 12348 29262 12350 29314
rect 12402 29262 12404 29314
rect 12236 29092 12292 29102
rect 12124 28756 12180 28766
rect 11788 27860 11844 27870
rect 11788 27766 11844 27804
rect 11452 26898 11508 26908
rect 11676 26964 11732 26974
rect 11676 26870 11732 26908
rect 11116 26178 11172 26190
rect 11116 26126 11118 26178
rect 11170 26126 11172 26178
rect 11116 25172 11172 26126
rect 11116 25106 11172 25116
rect 11900 25172 11956 25182
rect 10108 24782 10110 24834
rect 10162 24782 10164 24834
rect 10108 24770 10164 24782
rect 10332 24724 10388 24734
rect 10332 24630 10388 24668
rect 11004 24724 11060 25004
rect 11004 24630 11060 24668
rect 11452 24724 11508 24734
rect 11452 24630 11508 24668
rect 11900 24722 11956 25116
rect 11900 24670 11902 24722
rect 11954 24670 11956 24722
rect 11900 24658 11956 24670
rect 9324 23772 9604 23828
rect 10892 24610 10948 24622
rect 10892 24558 10894 24610
rect 10946 24558 10948 24610
rect 9324 22594 9380 23772
rect 9324 22542 9326 22594
rect 9378 22542 9380 22594
rect 9324 22530 9380 22542
rect 9884 23714 9940 23726
rect 9884 23662 9886 23714
rect 9938 23662 9940 23714
rect 9212 22372 9268 22382
rect 8988 22316 9212 22372
rect 9212 22278 9268 22316
rect 9884 22148 9940 23662
rect 10536 23548 10800 23558
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10536 23482 10800 23492
rect 10332 23044 10388 23054
rect 10332 22372 10388 22988
rect 9884 22082 9940 22092
rect 10108 22146 10164 22158
rect 10108 22094 10110 22146
rect 10162 22094 10164 22146
rect 9660 21812 9716 21822
rect 9660 21718 9716 21756
rect 9100 21700 9156 21710
rect 9100 21606 9156 21644
rect 9548 21474 9604 21486
rect 9548 21422 9550 21474
rect 9602 21422 9604 21474
rect 9548 20804 9604 21422
rect 9548 20738 9604 20748
rect 9996 21476 10052 21486
rect 8652 18162 8708 18172
rect 8764 20244 8820 20254
rect 8764 19906 8820 20188
rect 8764 19854 8766 19906
rect 8818 19854 8820 19906
rect 7980 17668 8036 17678
rect 8652 17668 8708 17678
rect 6972 17444 7028 17454
rect 6972 16994 7028 17388
rect 6972 16942 6974 16994
rect 7026 16942 7028 16994
rect 6972 16930 7028 16942
rect 6860 16706 6916 16716
rect 7532 16772 7588 16782
rect 5874 16492 6138 16502
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 5874 16426 6138 16436
rect 7532 16210 7588 16716
rect 7980 16770 8036 17612
rect 7980 16718 7982 16770
rect 8034 16718 8036 16770
rect 7980 16706 8036 16718
rect 8428 17666 8708 17668
rect 8428 17614 8654 17666
rect 8706 17614 8708 17666
rect 8428 17612 8708 17614
rect 7532 16158 7534 16210
rect 7586 16158 7588 16210
rect 7532 16146 7588 16158
rect 8092 16212 8148 16222
rect 5852 16100 5908 16110
rect 5740 16098 5908 16100
rect 5740 16046 5854 16098
rect 5906 16046 5908 16098
rect 5740 16044 5908 16046
rect 4956 14756 5012 14766
rect 4956 14418 5012 14700
rect 4956 14366 4958 14418
rect 5010 14366 5012 14418
rect 4956 14354 5012 14366
rect 3836 13022 3838 13074
rect 3890 13022 3892 13074
rect 3836 13010 3892 13022
rect 4060 13468 4900 13524
rect 4060 11506 4116 13468
rect 4508 13300 4564 13310
rect 4508 12402 4564 13244
rect 4956 12852 5012 12862
rect 5180 12852 5236 16044
rect 5628 15988 5684 15998
rect 5628 15894 5684 15932
rect 5292 15876 5348 15886
rect 5292 15428 5348 15820
rect 5740 15652 5796 16044
rect 5852 16034 5908 16044
rect 7756 16098 7812 16110
rect 7756 16046 7758 16098
rect 7810 16046 7812 16098
rect 6412 15876 6468 15886
rect 6412 15782 6468 15820
rect 7420 15876 7476 15886
rect 7756 15876 7812 16046
rect 7420 15874 7700 15876
rect 7420 15822 7422 15874
rect 7474 15822 7700 15874
rect 7420 15820 7700 15822
rect 7420 15810 7476 15820
rect 5628 15596 5796 15652
rect 5292 15372 5572 15428
rect 5292 15314 5348 15372
rect 5292 15262 5294 15314
rect 5346 15262 5348 15314
rect 5292 15250 5348 15262
rect 5404 15090 5460 15102
rect 5404 15038 5406 15090
rect 5458 15038 5460 15090
rect 4956 12850 5236 12852
rect 4956 12798 4958 12850
rect 5010 12798 5236 12850
rect 4956 12796 5236 12798
rect 5292 13522 5348 13534
rect 5292 13470 5294 13522
rect 5346 13470 5348 13522
rect 4956 12786 5012 12796
rect 4508 12350 4510 12402
rect 4562 12350 4564 12402
rect 4508 12338 4564 12350
rect 5292 12180 5348 13470
rect 4060 11454 4062 11506
rect 4114 11454 4116 11506
rect 4060 11442 4116 11454
rect 5180 12124 5348 12180
rect 4732 10724 4788 10734
rect 4732 10630 4788 10668
rect 3500 9886 3502 9938
rect 3554 9886 3556 9938
rect 3500 9874 3556 9886
rect 4732 10052 4788 10062
rect 2380 9662 2382 9714
rect 2434 9662 2436 9714
rect 2380 9650 2436 9662
rect 3052 9042 3108 9054
rect 3052 8990 3054 9042
rect 3106 8990 3108 9042
rect 3052 8932 3108 8990
rect 2156 8876 3052 8932
rect 2156 8428 2212 8876
rect 3052 8838 3108 8876
rect 3724 9042 3780 9054
rect 3724 8990 3726 9042
rect 3778 8990 3780 9042
rect 1820 8372 2212 8428
rect 2268 8372 2324 8382
rect 1820 7474 1876 8372
rect 1820 7422 1822 7474
rect 1874 7422 1876 7474
rect 1820 7410 1876 7422
rect 2268 7474 2324 8316
rect 3612 8372 3668 8382
rect 3612 8278 3668 8316
rect 2268 7422 2270 7474
rect 2322 7422 2324 7474
rect 2268 7410 2324 7422
rect 3724 5796 3780 8990
rect 4732 7698 4788 9996
rect 4956 9940 5012 9950
rect 4956 8146 5012 9884
rect 4956 8094 4958 8146
rect 5010 8094 5012 8146
rect 4956 8082 5012 8094
rect 5180 8148 5236 12124
rect 5292 11954 5348 11966
rect 5292 11902 5294 11954
rect 5346 11902 5348 11954
rect 5292 10500 5348 11902
rect 5292 10434 5348 10444
rect 5404 9940 5460 15038
rect 5516 13748 5572 15372
rect 5628 14420 5684 15596
rect 5964 15540 6020 15550
rect 5740 15538 6020 15540
rect 5740 15486 5966 15538
rect 6018 15486 6020 15538
rect 5740 15484 6020 15486
rect 5740 14644 5796 15484
rect 5964 15474 6020 15484
rect 7084 15316 7140 15326
rect 5874 14924 6138 14934
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 5874 14858 6138 14868
rect 5852 14644 5908 14654
rect 5740 14642 5908 14644
rect 5740 14590 5854 14642
rect 5906 14590 5908 14642
rect 5740 14588 5908 14590
rect 5852 14578 5908 14588
rect 5628 14418 5796 14420
rect 5628 14366 5630 14418
rect 5682 14366 5796 14418
rect 5628 14364 5796 14366
rect 5628 14354 5684 14364
rect 5628 13748 5684 13758
rect 5516 13746 5684 13748
rect 5516 13694 5630 13746
rect 5682 13694 5684 13746
rect 5516 13692 5684 13694
rect 5628 12180 5684 13692
rect 5740 13524 5796 14364
rect 7084 14418 7140 15260
rect 7084 14366 7086 14418
rect 7138 14366 7140 14418
rect 7084 14354 7140 14366
rect 7644 13972 7700 15820
rect 7756 15810 7812 15820
rect 8092 14642 8148 16156
rect 8316 16100 8372 16110
rect 8316 16006 8372 16044
rect 8092 14590 8094 14642
rect 8146 14590 8148 14642
rect 8092 14578 8148 14590
rect 8316 13972 8372 13982
rect 7644 13970 8372 13972
rect 7644 13918 8318 13970
rect 8370 13918 8372 13970
rect 7644 13916 8372 13918
rect 8316 13906 8372 13916
rect 6076 13746 6132 13758
rect 6076 13694 6078 13746
rect 6130 13694 6132 13746
rect 6076 13524 6132 13694
rect 6076 13468 6692 13524
rect 5740 12964 5796 13468
rect 5874 13356 6138 13366
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 5874 13290 6138 13300
rect 5964 12964 6020 12974
rect 5740 12962 6020 12964
rect 5740 12910 5966 12962
rect 6018 12910 6020 12962
rect 5740 12908 6020 12910
rect 5964 12852 6020 12908
rect 5964 12786 6020 12796
rect 6188 12852 6244 12862
rect 6188 12850 6356 12852
rect 6188 12798 6190 12850
rect 6242 12798 6356 12850
rect 6188 12796 6356 12798
rect 6188 12786 6244 12796
rect 5516 11284 5572 11294
rect 5516 10834 5572 11228
rect 5628 11172 5684 12124
rect 5964 12178 6020 12190
rect 5964 12126 5966 12178
rect 6018 12126 6020 12178
rect 5964 11956 6020 12126
rect 5964 11890 6020 11900
rect 5874 11788 6138 11798
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 5874 11722 6138 11732
rect 5740 11172 5796 11182
rect 5628 11170 5796 11172
rect 5628 11118 5742 11170
rect 5794 11118 5796 11170
rect 5628 11116 5796 11118
rect 5516 10782 5518 10834
rect 5570 10782 5572 10834
rect 5516 10770 5572 10782
rect 5404 9874 5460 9884
rect 5180 8082 5236 8092
rect 5516 9602 5572 9614
rect 5516 9550 5518 9602
rect 5570 9550 5572 9602
rect 4732 7646 4734 7698
rect 4786 7646 4788 7698
rect 4732 7634 4788 7646
rect 5292 7250 5348 7262
rect 5292 7198 5294 7250
rect 5346 7198 5348 7250
rect 5292 6020 5348 7198
rect 5516 6020 5572 9550
rect 5628 8932 5684 8942
rect 5740 8932 5796 11116
rect 5874 10220 6138 10230
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 5874 10154 6138 10164
rect 6300 10052 6356 12796
rect 6524 12850 6580 12862
rect 6524 12798 6526 12850
rect 6578 12798 6580 12850
rect 6188 9996 6356 10052
rect 6412 11172 6468 11182
rect 6188 9266 6244 9996
rect 6300 9716 6356 9726
rect 6412 9716 6468 11116
rect 6524 10052 6580 12798
rect 6524 9986 6580 9996
rect 6300 9714 6468 9716
rect 6300 9662 6302 9714
rect 6354 9662 6468 9714
rect 6300 9660 6468 9662
rect 6300 9650 6356 9660
rect 6188 9214 6190 9266
rect 6242 9214 6244 9266
rect 6188 9202 6244 9214
rect 5684 8876 5796 8932
rect 5628 7698 5684 8876
rect 5874 8652 6138 8662
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 5874 8586 6138 8596
rect 6076 8148 6132 8158
rect 6076 8054 6132 8092
rect 5628 7646 5630 7698
rect 5682 7646 5684 7698
rect 5628 7634 5684 7646
rect 6636 7700 6692 13468
rect 7644 12962 7700 12974
rect 8204 12964 8260 12974
rect 7644 12910 7646 12962
rect 7698 12910 7700 12962
rect 6860 12852 6916 12862
rect 6860 11844 6916 12796
rect 7308 12740 7364 12750
rect 7644 12740 7700 12910
rect 7308 12738 7700 12740
rect 7308 12686 7310 12738
rect 7362 12686 7700 12738
rect 7308 12684 7700 12686
rect 7980 12962 8260 12964
rect 7980 12910 8206 12962
rect 8258 12910 8260 12962
rect 7980 12908 8260 12910
rect 7308 12180 7364 12684
rect 7308 12114 7364 12124
rect 6860 11778 6916 11788
rect 7868 11844 7924 11854
rect 7868 11506 7924 11788
rect 7868 11454 7870 11506
rect 7922 11454 7924 11506
rect 7868 11442 7924 11454
rect 7532 11284 7588 11294
rect 7532 11190 7588 11228
rect 7756 10612 7812 10622
rect 7644 10610 7812 10612
rect 7644 10558 7758 10610
rect 7810 10558 7812 10610
rect 7644 10556 7812 10558
rect 6748 10500 6804 10510
rect 6804 10444 6916 10500
rect 6748 10434 6804 10444
rect 6636 7634 6692 7644
rect 6748 8818 6804 8830
rect 6748 8766 6750 8818
rect 6802 8766 6804 8818
rect 6748 7364 6804 8766
rect 6860 7586 6916 10444
rect 7084 8932 7140 8942
rect 7084 8838 7140 8876
rect 7308 8372 7364 8382
rect 7308 8278 7364 8316
rect 6860 7534 6862 7586
rect 6914 7534 6916 7586
rect 6860 7522 6916 7534
rect 6636 7308 6804 7364
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 6636 6578 6692 7308
rect 7644 6802 7700 10556
rect 7756 10546 7812 10556
rect 7980 10164 8036 12908
rect 8204 12898 8260 12908
rect 8316 12292 8372 12302
rect 8316 12198 8372 12236
rect 8092 12180 8148 12190
rect 8092 11732 8148 12124
rect 8092 11396 8148 11676
rect 8092 11394 8260 11396
rect 8092 11342 8094 11394
rect 8146 11342 8260 11394
rect 8092 11340 8260 11342
rect 8092 11330 8148 11340
rect 8204 10836 8260 11340
rect 8204 10610 8260 10780
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 8204 10546 8260 10558
rect 8428 10612 8484 17612
rect 8652 17602 8708 17612
rect 8764 17108 8820 19854
rect 9996 19234 10052 21420
rect 10108 21140 10164 22094
rect 10108 21074 10164 21084
rect 10332 20188 10388 22316
rect 10536 21980 10800 21990
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10536 21914 10800 21924
rect 10892 20578 10948 24558
rect 12124 23938 12180 28700
rect 12236 27858 12292 29036
rect 12236 27806 12238 27858
rect 12290 27806 12292 27858
rect 12236 27794 12292 27806
rect 12348 27412 12404 29262
rect 12348 27346 12404 27356
rect 12460 27298 12516 29484
rect 13356 29540 13412 29550
rect 13356 29446 13412 29484
rect 14476 29092 14532 30270
rect 31052 30322 31108 30334
rect 31052 30270 31054 30322
rect 31106 30270 31108 30322
rect 15708 30100 15764 30110
rect 15708 30098 15876 30100
rect 15708 30046 15710 30098
rect 15762 30046 15876 30098
rect 15708 30044 15876 30046
rect 15708 30034 15764 30044
rect 15260 29314 15316 29326
rect 15260 29262 15262 29314
rect 15314 29262 15316 29314
rect 15260 29204 15316 29262
rect 14476 29026 14532 29036
rect 15036 29148 15316 29204
rect 13020 28532 13076 28542
rect 12460 27246 12462 27298
rect 12514 27246 12516 27298
rect 12460 27234 12516 27246
rect 12572 27860 12628 27870
rect 12572 27076 12628 27804
rect 12572 26290 12628 27020
rect 12572 26238 12574 26290
rect 12626 26238 12628 26290
rect 12460 25282 12516 25294
rect 12460 25230 12462 25282
rect 12514 25230 12516 25282
rect 12460 24052 12516 25230
rect 12572 24724 12628 26238
rect 13020 26290 13076 28476
rect 15036 28532 15092 29148
rect 15198 29036 15462 29046
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15198 28970 15462 28980
rect 15260 28756 15316 28766
rect 15260 28662 15316 28700
rect 15708 28756 15764 28766
rect 15036 28466 15092 28476
rect 14700 28082 14756 28094
rect 15372 28084 15428 28094
rect 14700 28030 14702 28082
rect 14754 28030 14756 28082
rect 13244 27748 13300 27758
rect 13020 26238 13022 26290
rect 13074 26238 13076 26290
rect 13020 26226 13076 26238
rect 13132 27692 13244 27748
rect 13020 25732 13076 25742
rect 13132 25732 13188 27692
rect 13244 27682 13300 27692
rect 13692 27074 13748 27086
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 13468 26964 13524 26974
rect 13468 26870 13524 26908
rect 13020 25730 13188 25732
rect 13020 25678 13022 25730
rect 13074 25678 13188 25730
rect 13020 25676 13188 25678
rect 13692 26180 13748 27022
rect 14588 27076 14644 27086
rect 14588 26982 14644 27020
rect 14700 26516 14756 28030
rect 15260 28028 15372 28084
rect 15260 27970 15316 28028
rect 15372 28018 15428 28028
rect 15260 27918 15262 27970
rect 15314 27918 15316 27970
rect 15260 27906 15316 27918
rect 15198 27468 15462 27478
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15198 27402 15462 27412
rect 15260 27076 15316 27086
rect 15708 27076 15764 28700
rect 15820 27748 15876 30044
rect 19860 29820 20124 29830
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 19860 29754 20124 29764
rect 29184 29820 29448 29830
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29184 29754 29448 29764
rect 16268 29538 16324 29550
rect 16268 29486 16270 29538
rect 16322 29486 16324 29538
rect 15820 27682 15876 27692
rect 16044 28532 16100 28542
rect 15260 27074 15764 27076
rect 15260 27022 15262 27074
rect 15314 27022 15764 27074
rect 15260 27020 15764 27022
rect 15260 27010 15316 27020
rect 14700 26450 14756 26460
rect 16044 26514 16100 28476
rect 16268 28084 16324 29486
rect 29820 29540 29876 29550
rect 29820 29538 30100 29540
rect 29820 29486 29822 29538
rect 29874 29486 30100 29538
rect 29820 29484 30100 29486
rect 29820 29474 29876 29484
rect 28476 29314 28532 29326
rect 28476 29262 28478 29314
rect 28530 29262 28532 29314
rect 24522 29036 24786 29046
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24522 28970 24786 28980
rect 18060 28756 18116 28766
rect 18060 28662 18116 28700
rect 27020 28754 27076 28766
rect 27020 28702 27022 28754
rect 27074 28702 27076 28754
rect 16268 28018 16324 28028
rect 16604 28530 16660 28542
rect 16604 28478 16606 28530
rect 16658 28478 16660 28530
rect 16044 26462 16046 26514
rect 16098 26462 16100 26514
rect 16044 26450 16100 26462
rect 16380 26516 16436 26526
rect 16380 26422 16436 26460
rect 16604 26516 16660 28478
rect 19068 28532 19124 28542
rect 19068 28438 19124 28476
rect 26012 28532 26068 28542
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 18284 27972 18340 27982
rect 18284 27298 18340 27916
rect 19628 27972 19684 27982
rect 19628 27878 19684 27916
rect 21084 27972 21140 27982
rect 18284 27246 18286 27298
rect 18338 27246 18340 27298
rect 18284 27234 18340 27246
rect 18620 27746 18676 27758
rect 18620 27694 18622 27746
rect 18674 27694 18676 27746
rect 16604 26450 16660 26460
rect 17500 26850 17556 26862
rect 17500 26798 17502 26850
rect 17554 26798 17556 26850
rect 13020 25666 13076 25676
rect 13692 25396 13748 26124
rect 14140 26404 14196 26414
rect 14140 25618 14196 26348
rect 15260 26404 15316 26414
rect 15260 26310 15316 26348
rect 16268 26180 16324 26190
rect 16268 26086 16324 26124
rect 15198 25900 15462 25910
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15198 25834 15462 25844
rect 16716 25844 16772 25854
rect 14140 25566 14142 25618
rect 14194 25566 14196 25618
rect 14140 25554 14196 25566
rect 15932 25620 15988 25630
rect 15932 25618 16212 25620
rect 15932 25566 15934 25618
rect 15986 25566 16212 25618
rect 15932 25564 16212 25566
rect 15932 25554 15988 25564
rect 13804 25396 13860 25406
rect 13692 25394 13860 25396
rect 13692 25342 13806 25394
rect 13858 25342 13860 25394
rect 13692 25340 13860 25342
rect 13692 25060 13748 25340
rect 13804 25330 13860 25340
rect 14924 25396 14980 25406
rect 14924 25394 15092 25396
rect 14924 25342 14926 25394
rect 14978 25342 15092 25394
rect 14924 25340 15092 25342
rect 14924 25330 14980 25340
rect 12628 24668 12740 24724
rect 12572 24658 12628 24668
rect 12460 23986 12516 23996
rect 12124 23886 12126 23938
rect 12178 23886 12180 23938
rect 12124 23874 12180 23886
rect 12572 23938 12628 23950
rect 12572 23886 12574 23938
rect 12626 23886 12628 23938
rect 11452 23828 11508 23838
rect 11452 21026 11508 23772
rect 12572 23044 12628 23886
rect 12572 22978 12628 22988
rect 12684 23492 12740 24668
rect 13468 24052 13524 24062
rect 13468 23958 13524 23996
rect 12348 22372 12404 22382
rect 12684 22372 12740 23436
rect 13692 23938 13748 25004
rect 15036 24946 15092 25340
rect 15036 24894 15038 24946
rect 15090 24894 15092 24946
rect 15036 24882 15092 24894
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 12796 22372 12852 22382
rect 12684 22370 13412 22372
rect 12684 22318 12798 22370
rect 12850 22318 13412 22370
rect 12684 22316 13412 22318
rect 12348 22278 12404 22316
rect 12796 22306 12852 22316
rect 12684 21812 12740 21822
rect 11564 21476 11620 21486
rect 11564 21382 11620 21420
rect 11452 20974 11454 21026
rect 11506 20974 11508 21026
rect 11452 20962 11508 20974
rect 12460 21140 12516 21150
rect 10892 20526 10894 20578
rect 10946 20526 10948 20578
rect 10892 20514 10948 20526
rect 11900 20802 11956 20814
rect 11900 20750 11902 20802
rect 11954 20750 11956 20802
rect 11900 20580 11956 20750
rect 10536 20412 10800 20422
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10536 20346 10800 20356
rect 11564 20244 11620 20254
rect 11900 20188 11956 20524
rect 10332 20132 10500 20188
rect 9996 19182 9998 19234
rect 10050 19182 10052 19234
rect 9996 19170 10052 19182
rect 10444 19234 10500 20132
rect 11004 20130 11060 20142
rect 11564 20132 11956 20188
rect 11004 20078 11006 20130
rect 11058 20078 11060 20130
rect 11004 19460 11060 20078
rect 11004 19394 11060 19404
rect 10444 19182 10446 19234
rect 10498 19182 10500 19234
rect 10444 19170 10500 19182
rect 11116 19122 11172 19134
rect 11116 19070 11118 19122
rect 11170 19070 11172 19122
rect 11116 19012 11172 19070
rect 11452 19124 11508 19134
rect 11452 19030 11508 19068
rect 11788 19122 11844 19134
rect 11788 19070 11790 19122
rect 11842 19070 11844 19122
rect 10536 18844 10800 18854
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10536 18778 10800 18788
rect 10332 18564 10388 18574
rect 8988 18340 9044 18350
rect 8988 18246 9044 18284
rect 9772 18338 9828 18350
rect 9772 18286 9774 18338
rect 9826 18286 9828 18338
rect 9100 17668 9156 17678
rect 9324 17668 9380 17678
rect 9772 17668 9828 18286
rect 10108 18340 10164 18350
rect 10108 18246 10164 18284
rect 10332 18338 10388 18508
rect 11004 18564 11060 18574
rect 11116 18564 11172 18956
rect 11788 19012 11844 19070
rect 11788 18946 11844 18956
rect 11060 18508 11172 18564
rect 11004 18470 11060 18508
rect 11900 18452 11956 20132
rect 12012 20804 12068 20814
rect 12012 19906 12068 20748
rect 12012 19854 12014 19906
rect 12066 19854 12068 19906
rect 12012 19842 12068 19854
rect 12460 19346 12516 21084
rect 12460 19294 12462 19346
rect 12514 19294 12516 19346
rect 12460 19282 12516 19294
rect 12684 21026 12740 21756
rect 12684 20974 12686 21026
rect 12738 20974 12740 21026
rect 12684 19234 12740 20974
rect 12908 21698 12964 21710
rect 12908 21646 12910 21698
rect 12962 21646 12964 21698
rect 12684 19182 12686 19234
rect 12738 19182 12740 19234
rect 12684 19170 12740 19182
rect 12796 20580 12852 20590
rect 11676 18396 11956 18452
rect 12124 19122 12180 19134
rect 12124 19070 12126 19122
rect 12178 19070 12180 19122
rect 10332 18286 10334 18338
rect 10386 18286 10388 18338
rect 9100 17666 9828 17668
rect 9100 17614 9102 17666
rect 9154 17614 9326 17666
rect 9378 17614 9828 17666
rect 9100 17612 9828 17614
rect 9884 17666 9940 17678
rect 9884 17614 9886 17666
rect 9938 17614 9940 17666
rect 8988 17108 9044 17118
rect 8764 17106 9044 17108
rect 8764 17054 8990 17106
rect 9042 17054 9044 17106
rect 8764 17052 9044 17054
rect 8988 17042 9044 17052
rect 8540 16770 8596 16782
rect 8540 16718 8542 16770
rect 8594 16718 8596 16770
rect 8540 15876 8596 16718
rect 8540 15810 8596 15820
rect 9100 15428 9156 17612
rect 9324 17602 9380 17612
rect 9884 16212 9940 17614
rect 9996 16884 10052 16894
rect 9996 16790 10052 16828
rect 10332 16772 10388 18286
rect 10780 18340 10836 18350
rect 11564 18340 11620 18350
rect 11676 18340 11732 18396
rect 10780 18338 10948 18340
rect 10780 18286 10782 18338
rect 10834 18286 10948 18338
rect 10780 18284 10948 18286
rect 10780 18274 10836 18284
rect 10536 17276 10800 17286
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10536 17210 10800 17220
rect 10780 16996 10836 17006
rect 10780 16902 10836 16940
rect 10332 16706 10388 16716
rect 9884 16146 9940 16156
rect 10892 15874 10948 18284
rect 11564 18338 11732 18340
rect 11564 18286 11566 18338
rect 11618 18286 11732 18338
rect 11564 18284 11732 18286
rect 11564 16996 11620 18284
rect 11788 18226 11844 18238
rect 11788 18174 11790 18226
rect 11842 18174 11844 18226
rect 11788 17444 11844 18174
rect 11788 17378 11844 17388
rect 12124 17108 12180 19070
rect 12348 19124 12404 19134
rect 12348 18674 12404 19068
rect 12348 18622 12350 18674
rect 12402 18622 12404 18674
rect 12348 18610 12404 18622
rect 12124 17042 12180 17052
rect 12460 17442 12516 17454
rect 12460 17390 12462 17442
rect 12514 17390 12516 17442
rect 11564 16930 11620 16940
rect 11340 16884 11396 16894
rect 11340 16790 11396 16828
rect 11788 16882 11844 16894
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 10892 15822 10894 15874
rect 10946 15822 10948 15874
rect 10892 15810 10948 15822
rect 11452 15874 11508 15886
rect 11452 15822 11454 15874
rect 11506 15822 11508 15874
rect 10536 15708 10800 15718
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10536 15642 10800 15652
rect 8428 10546 8484 10556
rect 8540 15314 8596 15326
rect 8540 15262 8542 15314
rect 8594 15262 8596 15314
rect 8540 10276 8596 15262
rect 9100 15314 9156 15372
rect 9100 15262 9102 15314
rect 9154 15262 9156 15314
rect 8652 14308 8708 14318
rect 9100 14308 9156 15262
rect 11452 15316 11508 15822
rect 11452 15250 11508 15260
rect 10108 15204 10164 15214
rect 10108 14418 10164 15148
rect 10108 14366 10110 14418
rect 10162 14366 10164 14418
rect 10108 14354 10164 14366
rect 8652 14306 9156 14308
rect 8652 14254 8654 14306
rect 8706 14254 9102 14306
rect 9154 14254 9156 14306
rect 8652 14252 9156 14254
rect 8652 14242 8708 14252
rect 9100 13748 9156 14252
rect 9324 14308 9380 14318
rect 9324 14306 9604 14308
rect 9324 14254 9326 14306
rect 9378 14254 9604 14306
rect 9324 14252 9604 14254
rect 9324 14242 9380 14252
rect 9436 13748 9492 13758
rect 9100 13746 9492 13748
rect 9100 13694 9438 13746
rect 9490 13694 9492 13746
rect 9100 13692 9492 13694
rect 9436 13682 9492 13692
rect 9100 13524 9156 13534
rect 9100 13522 9268 13524
rect 9100 13470 9102 13522
rect 9154 13470 9268 13522
rect 9100 13468 9268 13470
rect 9100 13458 9156 13468
rect 9100 11954 9156 11966
rect 9100 11902 9102 11954
rect 9154 11902 9156 11954
rect 7756 10108 8036 10164
rect 8428 10220 8596 10276
rect 8652 11394 8708 11406
rect 8652 11342 8654 11394
rect 8706 11342 8708 11394
rect 7756 7364 7812 10108
rect 8428 9940 8484 10220
rect 8316 9884 8484 9940
rect 8316 8372 8372 9884
rect 8540 9828 8596 9838
rect 7756 7298 7812 7308
rect 7868 8316 8372 8372
rect 8428 9826 8596 9828
rect 8428 9774 8542 9826
rect 8594 9774 8596 9826
rect 8428 9772 8596 9774
rect 7868 7362 7924 8316
rect 8428 7812 8484 9772
rect 8540 9762 8596 9772
rect 8652 8596 8708 11342
rect 8764 10836 8820 10846
rect 8820 10780 9044 10836
rect 8764 10742 8820 10780
rect 8764 10612 8820 10622
rect 8820 10556 8932 10612
rect 8764 10546 8820 10556
rect 8764 8596 8820 8606
rect 8652 8540 8764 8596
rect 8764 8530 8820 8540
rect 8876 8372 8932 10556
rect 8988 10164 9044 10780
rect 8988 9826 9044 10108
rect 8988 9774 8990 9826
rect 9042 9774 9044 9826
rect 8988 9762 9044 9774
rect 8876 8306 8932 8316
rect 9100 8372 9156 11902
rect 9212 10052 9268 13468
rect 9548 12516 9604 14252
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 10108 13746 10164 13758
rect 10108 13694 10110 13746
rect 10162 13694 10164 13746
rect 10108 12964 10164 13694
rect 10108 12908 10948 12964
rect 9548 12450 9604 12460
rect 9772 12740 9828 12750
rect 9660 11284 9716 11294
rect 9660 10722 9716 11228
rect 9772 10834 9828 12684
rect 10556 12740 10612 12778
rect 10556 12674 10612 12684
rect 10536 12572 10800 12582
rect 10332 12516 10388 12526
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10536 12506 10800 12516
rect 10108 12292 10164 12302
rect 9772 10782 9774 10834
rect 9826 10782 9828 10834
rect 9772 10770 9828 10782
rect 9884 12066 9940 12078
rect 9884 12014 9886 12066
rect 9938 12014 9940 12066
rect 9884 11844 9940 12014
rect 10108 12066 10164 12236
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 10108 12002 10164 12014
rect 9660 10670 9662 10722
rect 9714 10670 9716 10722
rect 9660 10658 9716 10670
rect 9212 9986 9268 9996
rect 9660 10164 9716 10174
rect 9660 9266 9716 10108
rect 9884 9826 9940 11788
rect 10108 11172 10164 11182
rect 9996 11116 10108 11172
rect 9996 9938 10052 11116
rect 10108 11106 10164 11116
rect 10332 10724 10388 12460
rect 10668 12066 10724 12078
rect 10668 12014 10670 12066
rect 10722 12014 10724 12066
rect 10668 11954 10724 12014
rect 10668 11902 10670 11954
rect 10722 11902 10724 11954
rect 10668 11732 10724 11902
rect 10668 11666 10724 11676
rect 10536 11004 10800 11014
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10536 10938 10800 10948
rect 10444 10724 10500 10734
rect 10332 10722 10500 10724
rect 10332 10670 10446 10722
rect 10498 10670 10500 10722
rect 10332 10668 10500 10670
rect 10444 10658 10500 10668
rect 9996 9886 9998 9938
rect 10050 9886 10052 9938
rect 9996 9874 10052 9886
rect 9884 9774 9886 9826
rect 9938 9774 9940 9826
rect 9884 9762 9940 9774
rect 10536 9436 10800 9446
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10536 9370 10800 9380
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 9660 9202 9716 9214
rect 9100 8306 9156 8316
rect 10332 8596 10388 8606
rect 7868 7310 7870 7362
rect 7922 7310 7924 7362
rect 7868 7298 7924 7310
rect 7980 7756 8484 7812
rect 7644 6750 7646 6802
rect 7698 6750 7700 6802
rect 7644 6738 7700 6750
rect 6636 6526 6638 6578
rect 6690 6526 6692 6578
rect 6636 6514 6692 6526
rect 5740 6020 5796 6030
rect 5516 6018 5796 6020
rect 5516 5966 5742 6018
rect 5794 5966 5796 6018
rect 5516 5964 5796 5966
rect 5292 5954 5348 5964
rect 5740 5954 5796 5964
rect 6860 6020 6916 6030
rect 6860 5926 6916 5964
rect 4732 5796 4788 5806
rect 3724 5794 4788 5796
rect 3724 5742 4734 5794
rect 4786 5742 4788 5794
rect 3724 5740 4788 5742
rect 4732 5730 4788 5740
rect 7980 5794 8036 7756
rect 7980 5742 7982 5794
rect 8034 5742 8036 5794
rect 7980 5730 8036 5742
rect 10332 5796 10388 8540
rect 10892 8372 10948 12908
rect 11340 12740 11396 12750
rect 11116 12738 11396 12740
rect 11116 12686 11342 12738
rect 11394 12686 11396 12738
rect 11116 12684 11396 12686
rect 11004 11172 11060 11182
rect 11004 11078 11060 11116
rect 11116 10164 11172 12684
rect 11340 12674 11396 12684
rect 11676 12738 11732 12750
rect 11676 12686 11678 12738
rect 11730 12686 11732 12738
rect 11228 12068 11284 12078
rect 11676 12068 11732 12686
rect 11228 12066 11732 12068
rect 11228 12014 11230 12066
rect 11282 12014 11732 12066
rect 11228 12012 11732 12014
rect 11228 11954 11284 12012
rect 11228 11902 11230 11954
rect 11282 11902 11284 11954
rect 11228 11890 11284 11902
rect 11564 11732 11620 11742
rect 11116 10098 11172 10108
rect 11452 11676 11564 11732
rect 11452 9938 11508 11676
rect 11564 11666 11620 11676
rect 11676 11396 11732 12012
rect 11788 12066 11844 16830
rect 11788 12014 11790 12066
rect 11842 12014 11844 12066
rect 11788 12002 11844 12014
rect 12124 16772 12180 16782
rect 12124 15986 12180 16716
rect 12124 15934 12126 15986
rect 12178 15934 12180 15986
rect 12124 15316 12180 15934
rect 12124 12850 12180 15260
rect 12348 14532 12404 14542
rect 12124 12798 12126 12850
rect 12178 12798 12180 12850
rect 11676 11340 12068 11396
rect 11788 11172 11844 11182
rect 11788 11170 11956 11172
rect 11788 11118 11790 11170
rect 11842 11118 11956 11170
rect 11788 11116 11956 11118
rect 11788 11106 11844 11116
rect 11788 10500 11844 10510
rect 11788 10406 11844 10444
rect 11900 10276 11956 11116
rect 12012 11060 12068 11340
rect 12124 11284 12180 12798
rect 12236 14530 12404 14532
rect 12236 14478 12350 14530
rect 12402 14478 12404 14530
rect 12236 14476 12404 14478
rect 12236 11732 12292 14476
rect 12348 14466 12404 14476
rect 12236 11666 12292 11676
rect 12348 13858 12404 13870
rect 12348 13806 12350 13858
rect 12402 13806 12404 13858
rect 12348 11506 12404 13806
rect 12460 13074 12516 17390
rect 12796 16098 12852 20524
rect 12908 16772 12964 21646
rect 13244 21362 13300 21374
rect 13244 21310 13246 21362
rect 13298 21310 13300 21362
rect 13244 20916 13300 21310
rect 13244 20850 13300 20860
rect 13356 20018 13412 22316
rect 13692 21812 13748 23886
rect 14252 24834 14308 24846
rect 14252 24782 14254 24834
rect 14306 24782 14308 24834
rect 14028 23044 14084 23054
rect 13748 21756 13972 21812
rect 13692 21746 13748 21756
rect 13916 20916 13972 21756
rect 14028 21810 14084 22988
rect 14028 21758 14030 21810
rect 14082 21758 14084 21810
rect 14028 21746 14084 21758
rect 13916 20822 13972 20860
rect 14252 20914 14308 24782
rect 15198 24332 15462 24342
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15198 24266 15462 24276
rect 16044 23938 16100 23950
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 16044 23492 16100 23886
rect 14700 23156 14756 23166
rect 14700 23062 14756 23100
rect 15372 23156 15428 23166
rect 15372 23042 15428 23100
rect 15372 22990 15374 23042
rect 15426 22990 15428 23042
rect 15372 22932 15428 22990
rect 15372 22876 15652 22932
rect 15198 22764 15462 22774
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15198 22698 15462 22708
rect 15484 22372 15540 22382
rect 15596 22372 15652 22876
rect 15484 22370 15652 22372
rect 15484 22318 15486 22370
rect 15538 22318 15652 22370
rect 15484 22316 15652 22318
rect 16044 22482 16100 23436
rect 16044 22430 16046 22482
rect 16098 22430 16100 22482
rect 14252 20862 14254 20914
rect 14306 20862 14308 20914
rect 14252 20850 14308 20862
rect 14588 22148 14644 22158
rect 14588 20914 14644 22092
rect 15484 22148 15540 22316
rect 15484 22082 15540 22092
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 15036 21028 15092 21038
rect 14588 20862 14590 20914
rect 14642 20862 14644 20914
rect 14588 20850 14644 20862
rect 14812 20916 14868 20926
rect 14812 20802 14868 20860
rect 14812 20750 14814 20802
rect 14866 20750 14868 20802
rect 14812 20738 14868 20750
rect 13580 20580 13636 20590
rect 13580 20486 13636 20524
rect 13356 19966 13358 20018
rect 13410 19966 13412 20018
rect 13356 19954 13412 19966
rect 13804 20018 13860 20030
rect 13804 19966 13806 20018
rect 13858 19966 13860 20018
rect 13356 19460 13412 19470
rect 13356 19366 13412 19404
rect 13804 18676 13860 19966
rect 15036 19908 15092 20972
rect 16044 20802 16100 22430
rect 16156 21588 16212 25564
rect 16716 23938 16772 25788
rect 16716 23886 16718 23938
rect 16770 23886 16772 23938
rect 16716 23874 16772 23886
rect 17164 25506 17220 25518
rect 17164 25454 17166 25506
rect 17218 25454 17220 25506
rect 16716 23492 16772 23502
rect 16268 21588 16324 21598
rect 16156 21586 16324 21588
rect 16156 21534 16270 21586
rect 16322 21534 16324 21586
rect 16156 21532 16324 21534
rect 16268 21522 16324 21532
rect 16716 21586 16772 23436
rect 17164 23492 17220 25454
rect 17500 24834 17556 26798
rect 18508 26516 18564 26526
rect 17836 26180 17892 26190
rect 17836 25506 17892 26124
rect 17836 25454 17838 25506
rect 17890 25454 17892 25506
rect 17836 25442 17892 25454
rect 18508 24946 18564 26460
rect 18620 25844 18676 27694
rect 18620 25778 18676 25788
rect 18844 26962 18900 26974
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 18844 25284 18900 26910
rect 18844 25218 18900 25228
rect 18956 26850 19012 26862
rect 18956 26798 18958 26850
rect 19010 26798 19012 26850
rect 18508 24894 18510 24946
rect 18562 24894 18564 24946
rect 18508 24882 18564 24894
rect 17500 24782 17502 24834
rect 17554 24782 17556 24834
rect 17500 24770 17556 24782
rect 17164 23426 17220 23436
rect 17724 24722 17780 24734
rect 17724 24670 17726 24722
rect 17778 24670 17780 24722
rect 17724 23268 17780 24670
rect 18956 23826 19012 26798
rect 19860 26684 20124 26694
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 19860 26618 20124 26628
rect 21084 26514 21140 27916
rect 22316 27972 22372 27982
rect 22316 27878 22372 27916
rect 23436 27748 23492 27758
rect 22988 27746 23492 27748
rect 22988 27694 23438 27746
rect 23490 27694 23492 27746
rect 22988 27692 23492 27694
rect 22316 27074 22372 27086
rect 22316 27022 22318 27074
rect 22370 27022 22372 27074
rect 22316 26908 22372 27022
rect 22988 27074 23044 27692
rect 23436 27682 23492 27692
rect 24220 27748 24276 27758
rect 22988 27022 22990 27074
rect 23042 27022 23044 27074
rect 22988 27010 23044 27022
rect 21084 26462 21086 26514
rect 21138 26462 21140 26514
rect 21084 26450 21140 26462
rect 22204 26852 22372 26908
rect 20412 26404 20468 26414
rect 19740 26402 20468 26404
rect 19740 26350 20414 26402
rect 20466 26350 20468 26402
rect 19740 26348 20468 26350
rect 19404 26180 19460 26190
rect 19404 26086 19460 26124
rect 19292 24836 19348 24846
rect 19292 24742 19348 24780
rect 19740 24162 19796 26348
rect 20412 26338 20468 26348
rect 21868 26402 21924 26414
rect 21868 26350 21870 26402
rect 21922 26350 21924 26402
rect 21644 25620 21700 25630
rect 20860 25396 20916 25406
rect 20860 25302 20916 25340
rect 20188 25282 20244 25294
rect 20188 25230 20190 25282
rect 20242 25230 20244 25282
rect 19860 25116 20124 25126
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 19860 25050 20124 25060
rect 19740 24110 19742 24162
rect 19794 24110 19796 24162
rect 19740 24098 19796 24110
rect 20188 24050 20244 25230
rect 20188 23998 20190 24050
rect 20242 23998 20244 24050
rect 20188 23986 20244 23998
rect 20300 25284 20356 25294
rect 20300 23940 20356 25228
rect 21532 25284 21588 25294
rect 21308 24836 21364 24846
rect 21308 24050 21364 24780
rect 21308 23998 21310 24050
rect 21362 23998 21364 24050
rect 21308 23986 21364 23998
rect 20300 23938 20692 23940
rect 20300 23886 20302 23938
rect 20354 23886 20692 23938
rect 20300 23884 20692 23886
rect 20300 23874 20356 23884
rect 18956 23774 18958 23826
rect 19010 23774 19012 23826
rect 18956 23762 19012 23774
rect 19860 23548 20124 23558
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 19860 23482 20124 23492
rect 19516 23268 19572 23278
rect 17724 23266 17892 23268
rect 17724 23214 17726 23266
rect 17778 23214 17892 23266
rect 17724 23212 17892 23214
rect 17724 23202 17780 23212
rect 17388 23044 17444 23054
rect 17388 22950 17444 22988
rect 16716 21534 16718 21586
rect 16770 21534 16772 21586
rect 16716 21522 16772 21534
rect 17836 21700 17892 23212
rect 19404 23042 19460 23054
rect 19404 22990 19406 23042
rect 19458 22990 19460 23042
rect 19292 22372 19348 22382
rect 17836 21586 17892 21644
rect 18508 21700 18564 21710
rect 18508 21606 18564 21644
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 17612 21474 17668 21486
rect 17612 21422 17614 21474
rect 17666 21422 17668 21474
rect 16044 20750 16046 20802
rect 16098 20750 16100 20802
rect 16044 20188 16100 20750
rect 16380 20804 16436 20814
rect 16380 20710 16436 20748
rect 16716 20580 16772 20590
rect 16380 20244 16436 20282
rect 15036 19842 15092 19852
rect 15596 20132 16212 20188
rect 16380 20178 16436 20188
rect 15198 19628 15462 19638
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15198 19562 15462 19572
rect 14140 19012 14196 19022
rect 14140 18918 14196 18956
rect 13804 18610 13860 18620
rect 14924 18450 14980 18462
rect 14924 18398 14926 18450
rect 14978 18398 14980 18450
rect 14812 17892 14868 17902
rect 14700 17836 14812 17892
rect 13580 17666 13636 17678
rect 13580 17614 13582 17666
rect 13634 17614 13636 17666
rect 12908 16706 12964 16716
rect 13020 17442 13076 17454
rect 13020 17390 13022 17442
rect 13074 17390 13076 17442
rect 12796 16046 12798 16098
rect 12850 16046 12852 16098
rect 12796 16034 12852 16046
rect 12796 15428 12852 15438
rect 12796 15334 12852 15372
rect 13020 15148 13076 17390
rect 13580 16884 13636 17614
rect 13916 17668 13972 17678
rect 13916 17574 13972 17612
rect 14028 17108 14084 17118
rect 14028 17014 14084 17052
rect 13580 16100 13636 16828
rect 13580 16034 13636 16044
rect 14140 16100 14196 16110
rect 14140 16006 14196 16044
rect 14700 15986 14756 17836
rect 14812 17826 14868 17836
rect 14700 15934 14702 15986
rect 14754 15934 14756 15986
rect 14700 15922 14756 15934
rect 14812 16658 14868 16670
rect 14812 16606 14814 16658
rect 14866 16606 14868 16658
rect 13580 15874 13636 15886
rect 13580 15822 13582 15874
rect 13634 15822 13636 15874
rect 13580 15428 13636 15822
rect 14812 15540 14868 16606
rect 13580 15362 13636 15372
rect 14364 15484 14868 15540
rect 14924 15540 14980 18398
rect 15484 18452 15540 18462
rect 15596 18452 15652 20132
rect 16156 20020 16212 20132
rect 16156 19954 16212 19964
rect 16380 19236 16436 19246
rect 15484 18450 15652 18452
rect 15484 18398 15486 18450
rect 15538 18398 15652 18450
rect 15484 18396 15652 18398
rect 15932 19234 16436 19236
rect 15932 19182 16382 19234
rect 16434 19182 16436 19234
rect 15932 19180 16436 19182
rect 15484 18386 15540 18396
rect 15708 18338 15764 18350
rect 15708 18286 15710 18338
rect 15762 18286 15764 18338
rect 15198 18060 15462 18070
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15198 17994 15462 18004
rect 15260 17108 15316 17118
rect 15484 17108 15540 17118
rect 15260 17106 15484 17108
rect 15260 17054 15262 17106
rect 15314 17054 15484 17106
rect 15260 17052 15484 17054
rect 15260 17042 15316 17052
rect 15484 17042 15540 17052
rect 15198 16492 15462 16502
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15198 16426 15462 16436
rect 14924 15484 15652 15540
rect 12460 13022 12462 13074
rect 12514 13022 12516 13074
rect 12460 13010 12516 13022
rect 12796 15092 13076 15148
rect 12348 11454 12350 11506
rect 12402 11454 12404 11506
rect 12348 11442 12404 11454
rect 12460 12404 12516 12414
rect 12124 11190 12180 11228
rect 12236 11172 12292 11182
rect 12236 11060 12292 11116
rect 12012 11004 12292 11060
rect 12236 10834 12292 11004
rect 12236 10782 12238 10834
rect 12290 10782 12292 10834
rect 12236 10770 12292 10782
rect 12460 10612 12516 12348
rect 12796 12290 12852 15092
rect 12908 14700 13412 14756
rect 12908 14530 12964 14700
rect 12908 14478 12910 14530
rect 12962 14478 12964 14530
rect 12908 14466 12964 14478
rect 13020 14532 13076 14542
rect 13020 13074 13076 14476
rect 13356 13746 13412 14700
rect 13804 14532 13860 14542
rect 13804 14438 13860 14476
rect 13356 13694 13358 13746
rect 13410 13694 13412 13746
rect 13020 13022 13022 13074
rect 13074 13022 13076 13074
rect 13020 13010 13076 13022
rect 13132 13522 13188 13534
rect 13132 13470 13134 13522
rect 13186 13470 13188 13522
rect 12796 12238 12798 12290
rect 12850 12238 12852 12290
rect 12796 12226 12852 12238
rect 12908 11172 12964 11182
rect 12908 11078 12964 11116
rect 12460 10546 12516 10556
rect 13020 10388 13076 10398
rect 11452 9886 11454 9938
rect 11506 9886 11508 9938
rect 11452 9874 11508 9886
rect 11788 10220 11956 10276
rect 12012 10386 13076 10388
rect 12012 10334 13022 10386
rect 13074 10334 13076 10386
rect 12012 10332 13076 10334
rect 11788 9380 11844 10220
rect 11788 9314 11844 9324
rect 11900 10052 11956 10062
rect 11228 9044 11284 9054
rect 11228 8950 11284 8988
rect 11676 9042 11732 9054
rect 11676 8990 11678 9042
rect 11730 8990 11732 9042
rect 11452 8372 11508 8382
rect 10892 8370 11508 8372
rect 10892 8318 11454 8370
rect 11506 8318 11508 8370
rect 10892 8316 11508 8318
rect 11452 8306 11508 8316
rect 10536 7868 10800 7878
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10536 7802 10800 7812
rect 10668 7700 10724 7710
rect 10556 7364 10612 7374
rect 10556 7270 10612 7308
rect 10668 6802 10724 7644
rect 11676 7364 11732 8990
rect 11676 7298 11732 7308
rect 11788 8372 11844 8382
rect 10668 6750 10670 6802
rect 10722 6750 10724 6802
rect 10668 6738 10724 6750
rect 10536 6300 10800 6310
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10536 6234 10800 6244
rect 11788 6018 11844 8316
rect 11900 7586 11956 9996
rect 11900 7534 11902 7586
rect 11954 7534 11956 7586
rect 11900 7522 11956 7534
rect 12012 6578 12068 10332
rect 13020 10322 13076 10332
rect 12460 10164 12516 10174
rect 13132 10164 13188 13470
rect 13356 12964 13412 13694
rect 13916 13748 13972 13758
rect 13916 13746 14084 13748
rect 13916 13694 13918 13746
rect 13970 13694 14084 13746
rect 13916 13692 14084 13694
rect 13916 13682 13972 13692
rect 13468 12964 13524 12974
rect 13356 12962 13524 12964
rect 13356 12910 13470 12962
rect 13522 12910 13524 12962
rect 13356 12908 13524 12910
rect 13468 12180 13524 12908
rect 13916 12962 13972 12974
rect 13916 12910 13918 12962
rect 13970 12910 13972 12962
rect 13916 12404 13972 12910
rect 13916 12338 13972 12348
rect 13468 12178 13636 12180
rect 13468 12126 13470 12178
rect 13522 12126 13636 12178
rect 13468 12124 13636 12126
rect 13468 12114 13524 12124
rect 13580 11170 13636 12124
rect 13580 11118 13582 11170
rect 13634 11118 13636 11170
rect 13580 10612 13636 11118
rect 13916 12178 13972 12190
rect 13916 12126 13918 12178
rect 13970 12126 13972 12178
rect 13804 10724 13860 10734
rect 13804 10630 13860 10668
rect 13580 10546 13636 10556
rect 13916 10388 13972 12126
rect 13916 10322 13972 10332
rect 12460 8146 12516 10108
rect 12796 10108 13188 10164
rect 12796 9714 12852 10108
rect 14028 9940 14084 13692
rect 14364 11282 14420 15484
rect 14812 15314 14868 15326
rect 14812 15262 14814 15314
rect 14866 15262 14868 15314
rect 14812 14532 14868 15262
rect 15372 15314 15428 15326
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 15148 15204 15204 15214
rect 15148 15110 15204 15148
rect 15372 15204 15428 15262
rect 15372 15138 15428 15148
rect 15198 14924 15462 14934
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15198 14858 15462 14868
rect 14812 14466 14868 14476
rect 15198 13356 15462 13366
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15198 13290 15462 13300
rect 15198 11788 15462 11798
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15198 11722 15462 11732
rect 15372 11508 15428 11518
rect 15596 11508 15652 15484
rect 15708 15316 15764 18286
rect 15932 16210 15988 19180
rect 16380 19170 16436 19180
rect 16044 18340 16100 18350
rect 16044 18338 16324 18340
rect 16044 18286 16046 18338
rect 16098 18286 16324 18338
rect 16044 18284 16324 18286
rect 16044 18274 16100 18284
rect 16268 17554 16324 18284
rect 16268 17502 16270 17554
rect 16322 17502 16324 17554
rect 16268 17490 16324 17502
rect 16716 17108 16772 20524
rect 17612 20244 17668 21422
rect 17612 20178 17668 20188
rect 17276 20020 17332 20030
rect 16940 19794 16996 19806
rect 16940 19742 16942 19794
rect 16994 19742 16996 19794
rect 16716 16882 16772 17052
rect 16716 16830 16718 16882
rect 16770 16830 16772 16882
rect 16716 16818 16772 16830
rect 16828 18340 16884 18350
rect 15932 16158 15934 16210
rect 15986 16158 15988 16210
rect 15932 16146 15988 16158
rect 16044 16770 16100 16782
rect 16044 16718 16046 16770
rect 16098 16718 16100 16770
rect 15708 15250 15764 15260
rect 16044 15316 16100 16718
rect 16828 16436 16884 18284
rect 16940 17892 16996 19742
rect 17052 19236 17108 19246
rect 17276 19236 17332 19964
rect 17724 19348 17780 19358
rect 17836 19348 17892 21534
rect 19292 21586 19348 22316
rect 19292 21534 19294 21586
rect 19346 21534 19348 21586
rect 19292 21522 19348 21534
rect 18732 21474 18788 21486
rect 18732 21422 18734 21474
rect 18786 21422 18788 21474
rect 17948 21252 18004 21262
rect 17948 20018 18004 21196
rect 18732 20690 18788 21422
rect 19404 21252 19460 22990
rect 19404 21186 19460 21196
rect 19516 21026 19572 23212
rect 20412 23268 20468 23278
rect 20412 23174 20468 23212
rect 20636 22370 20692 23884
rect 21532 23938 21588 25228
rect 21644 24722 21700 25564
rect 21868 24948 21924 26350
rect 21868 24882 21924 24892
rect 22204 24724 22260 26852
rect 24220 26290 24276 27692
rect 25788 27524 25844 27534
rect 24522 27468 24786 27478
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24522 27402 24786 27412
rect 25452 26852 25508 26862
rect 25452 26850 25732 26852
rect 25452 26798 25454 26850
rect 25506 26798 25732 26850
rect 25452 26796 25732 26798
rect 25452 26786 25508 26796
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 24220 26226 24276 26238
rect 24668 26292 24724 26302
rect 24668 26198 24724 26236
rect 25340 26292 25396 26302
rect 24522 25900 24786 25910
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24522 25834 24786 25844
rect 22428 25620 22484 25630
rect 22428 25526 22484 25564
rect 23996 25620 24052 25630
rect 23548 25396 23604 25406
rect 23548 25302 23604 25340
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 21644 24658 21700 24670
rect 21868 24668 22204 24724
rect 21532 23886 21534 23938
rect 21586 23886 21588 23938
rect 21532 23874 21588 23886
rect 21308 23156 21364 23166
rect 21756 23156 21812 23166
rect 21308 23062 21364 23100
rect 21532 23154 21812 23156
rect 21532 23102 21758 23154
rect 21810 23102 21812 23154
rect 21532 23100 21812 23102
rect 20636 22318 20638 22370
rect 20690 22318 20692 22370
rect 20412 22258 20468 22270
rect 20412 22206 20414 22258
rect 20466 22206 20468 22258
rect 19740 22148 19796 22158
rect 19740 22054 19796 22092
rect 19860 21980 20124 21990
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 19860 21914 20124 21924
rect 19516 20974 19518 21026
rect 19570 20974 19572 21026
rect 19516 20962 19572 20974
rect 19628 21586 19684 21598
rect 19628 21534 19630 21586
rect 19682 21534 19684 21586
rect 18732 20638 18734 20690
rect 18786 20638 18788 20690
rect 18732 20626 18788 20638
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19954 18004 19966
rect 17724 19346 17892 19348
rect 17724 19294 17726 19346
rect 17778 19294 17892 19346
rect 17724 19292 17892 19294
rect 19516 19348 19572 19358
rect 19628 19348 19684 21534
rect 19860 20412 20124 20422
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 19860 20346 20124 20356
rect 20412 20242 20468 22206
rect 20636 21588 20692 22318
rect 20636 21522 20692 21532
rect 21308 21588 21364 21598
rect 20412 20190 20414 20242
rect 20466 20190 20468 20242
rect 20412 20178 20468 20190
rect 21308 20130 21364 21532
rect 21532 20244 21588 23100
rect 21756 23090 21812 23100
rect 21868 23156 21924 24668
rect 22204 24630 22260 24668
rect 23436 24724 23492 24734
rect 23436 23938 23492 24668
rect 23436 23886 23438 23938
rect 23490 23886 23492 23938
rect 23436 23874 23492 23886
rect 23996 23938 24052 25564
rect 25228 24948 25284 24958
rect 25228 24834 25284 24892
rect 25228 24782 25230 24834
rect 25282 24782 25284 24834
rect 25228 24770 25284 24782
rect 25340 24724 25396 26236
rect 25676 25732 25732 26796
rect 25788 26290 25844 27468
rect 26012 27298 26068 28476
rect 26012 27246 26014 27298
rect 26066 27246 26068 27298
rect 26012 27234 26068 27246
rect 26684 27858 26740 27870
rect 26684 27806 26686 27858
rect 26738 27806 26740 27858
rect 25788 26238 25790 26290
rect 25842 26238 25844 26290
rect 25788 26226 25844 26238
rect 25676 25676 25956 25732
rect 25564 25620 25620 25630
rect 25564 25526 25620 25564
rect 25900 24834 25956 25676
rect 25900 24782 25902 24834
rect 25954 24782 25956 24834
rect 25900 24770 25956 24782
rect 26572 25394 26628 25406
rect 26572 25342 26574 25394
rect 26626 25342 26628 25394
rect 25340 24658 25396 24668
rect 25564 24610 25620 24622
rect 25564 24558 25566 24610
rect 25618 24558 25620 24610
rect 24522 24332 24786 24342
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24522 24266 24786 24276
rect 23996 23886 23998 23938
rect 24050 23886 24052 23938
rect 23996 23874 24052 23886
rect 24780 24164 24836 24174
rect 24220 23380 24276 23390
rect 24220 23286 24276 23324
rect 24780 23378 24836 24108
rect 25564 23940 25620 24558
rect 25564 23874 25620 23884
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 23940 26292 24558
rect 26572 24164 26628 25342
rect 26684 24724 26740 27806
rect 27020 27524 27076 28702
rect 27132 28756 27188 28766
rect 27132 27858 27188 28700
rect 28028 28532 28084 28542
rect 28028 28438 28084 28476
rect 27132 27806 27134 27858
rect 27186 27806 27188 27858
rect 27132 27794 27188 27806
rect 28476 27748 28532 29262
rect 29932 28868 29988 28878
rect 28476 27682 28532 27692
rect 28812 28532 28868 28542
rect 27020 27458 27076 27468
rect 27580 26964 27636 26974
rect 27468 25508 27524 25518
rect 27580 25508 27636 26908
rect 28812 26514 28868 28476
rect 29596 28308 29652 28318
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 29372 27970 29428 27982
rect 29372 27918 29374 27970
rect 29426 27918 29428 27970
rect 29372 27186 29428 27918
rect 29372 27134 29374 27186
rect 29426 27134 29428 27186
rect 29372 27122 29428 27134
rect 29148 26964 29204 26974
rect 29148 26870 29204 26908
rect 29184 26684 29448 26694
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29184 26618 29448 26628
rect 28812 26462 28814 26514
rect 28866 26462 28868 26514
rect 28812 26450 28868 26462
rect 28028 26404 28084 26414
rect 27692 26402 28084 26404
rect 27692 26350 28030 26402
rect 28082 26350 28084 26402
rect 27692 26348 28084 26350
rect 27692 25618 27748 26348
rect 28028 26338 28084 26348
rect 27692 25566 27694 25618
rect 27746 25566 27748 25618
rect 27692 25554 27748 25566
rect 29148 26290 29204 26302
rect 29148 26238 29150 26290
rect 29202 26238 29204 26290
rect 27468 25506 27636 25508
rect 27468 25454 27470 25506
rect 27522 25454 27636 25506
rect 27468 25452 27636 25454
rect 29148 25508 29204 26238
rect 29596 26290 29652 28252
rect 29932 27972 29988 28812
rect 30044 28196 30100 29484
rect 30156 28756 30212 28766
rect 30156 28662 30212 28700
rect 31052 28308 31108 30270
rect 32060 30098 32116 30110
rect 32060 30046 32062 30098
rect 32114 30046 32116 30098
rect 32060 28868 32116 30046
rect 32060 28802 32116 28812
rect 31164 28532 31220 28542
rect 31164 28438 31220 28476
rect 31052 28242 31108 28252
rect 30044 28140 30436 28196
rect 30156 27972 30212 27982
rect 29932 27970 30212 27972
rect 29932 27918 30158 27970
rect 30210 27918 30212 27970
rect 29932 27916 30212 27918
rect 30156 27906 30212 27916
rect 30380 27298 30436 28140
rect 32284 27860 32340 27870
rect 32172 27858 32340 27860
rect 32172 27806 32286 27858
rect 32338 27806 32340 27858
rect 32172 27804 32340 27806
rect 32060 27748 32116 27758
rect 30380 27246 30382 27298
rect 30434 27246 30436 27298
rect 30380 27234 30436 27246
rect 31836 27746 32116 27748
rect 31836 27694 32062 27746
rect 32114 27694 32116 27746
rect 31836 27692 32116 27694
rect 29596 26238 29598 26290
rect 29650 26238 29652 26290
rect 29596 26226 29652 26238
rect 29708 27076 29764 27086
rect 29260 25508 29316 25518
rect 29148 25452 29260 25508
rect 27468 25442 27524 25452
rect 26684 24164 26740 24668
rect 27132 24722 27188 24734
rect 27132 24670 27134 24722
rect 27186 24670 27188 24722
rect 26684 24108 26964 24164
rect 26572 24098 26628 24108
rect 26236 23874 26292 23884
rect 26460 23828 26516 23838
rect 26460 23714 26516 23772
rect 26460 23662 26462 23714
rect 26514 23662 26516 23714
rect 26460 23650 26516 23662
rect 24780 23326 24782 23378
rect 24834 23326 24836 23378
rect 24780 23314 24836 23326
rect 21756 22372 21812 22382
rect 21868 22372 21924 23100
rect 26908 23042 26964 24108
rect 27132 24052 27188 24670
rect 27132 23986 27188 23996
rect 27580 23940 27636 25452
rect 29260 25414 29316 25452
rect 29708 25506 29764 27020
rect 31164 26852 31220 26862
rect 31164 26758 31220 26796
rect 29708 25454 29710 25506
rect 29762 25454 29764 25506
rect 29708 25442 29764 25454
rect 30156 26740 30212 26750
rect 29184 25116 29448 25126
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29184 25050 29448 25060
rect 29596 24948 29652 24958
rect 29596 24854 29652 24892
rect 30156 24946 30212 26684
rect 31836 26514 31892 27692
rect 32060 27682 32116 27692
rect 31836 26462 31838 26514
rect 31890 26462 31892 26514
rect 31836 26450 31892 26462
rect 32172 25508 32228 27804
rect 32284 27794 32340 27804
rect 32620 26514 32676 33180
rect 34076 33236 34132 33246
rect 34076 33142 34132 33180
rect 33846 32172 34110 32182
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 33846 32106 34110 32116
rect 34300 31890 34356 31902
rect 34300 31838 34302 31890
rect 34354 31838 34356 31890
rect 33846 30604 34110 30614
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 33846 30538 34110 30548
rect 33516 29428 33572 29438
rect 32956 28754 33012 28766
rect 32956 28702 32958 28754
rect 33010 28702 33012 28754
rect 32620 26462 32622 26514
rect 32674 26462 32676 26514
rect 32620 26450 32676 26462
rect 32732 28420 32788 28430
rect 32732 25730 32788 28364
rect 32956 27076 33012 28702
rect 33180 28532 33236 28542
rect 32956 27010 33012 27020
rect 33068 28476 33180 28532
rect 32956 26516 33012 26526
rect 33068 26516 33124 28476
rect 33180 28466 33236 28476
rect 33404 28196 33460 28206
rect 32956 26514 33124 26516
rect 32956 26462 32958 26514
rect 33010 26462 33124 26514
rect 32956 26460 33124 26462
rect 33180 26852 33236 26862
rect 32956 26450 33012 26460
rect 32732 25678 32734 25730
rect 32786 25678 32788 25730
rect 32732 25666 32788 25678
rect 33068 26292 33124 26302
rect 31948 25452 32228 25508
rect 33068 25508 33124 26236
rect 30156 24894 30158 24946
rect 30210 24894 30212 24946
rect 30156 24882 30212 24894
rect 30492 24948 30548 24958
rect 30492 24854 30548 24892
rect 31836 24724 31892 24734
rect 31948 24724 32004 25452
rect 33068 25414 33124 25452
rect 32060 25282 32116 25294
rect 32060 25230 32062 25282
rect 32114 25230 32116 25282
rect 32060 24834 32116 25230
rect 32060 24782 32062 24834
rect 32114 24782 32116 24834
rect 32060 24770 32116 24782
rect 33180 24834 33236 26796
rect 33404 25506 33460 28140
rect 33516 27074 33572 29372
rect 34300 29428 34356 31838
rect 34412 31108 34468 34078
rect 34524 33572 34580 34748
rect 34524 33506 34580 33516
rect 34636 34690 34692 34702
rect 34636 34638 34638 34690
rect 34690 34638 34692 34690
rect 34412 31042 34468 31052
rect 34300 29362 34356 29372
rect 34412 30882 34468 30894
rect 34412 30830 34414 30882
rect 34466 30830 34468 30882
rect 34076 29316 34132 29326
rect 34076 29314 34244 29316
rect 34076 29262 34078 29314
rect 34130 29262 34244 29314
rect 34076 29260 34244 29262
rect 34076 29250 34132 29260
rect 33846 29036 34110 29046
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 33846 28970 34110 28980
rect 34188 28756 34244 29260
rect 34188 28700 34356 28756
rect 34188 28530 34244 28542
rect 34188 28478 34190 28530
rect 34242 28478 34244 28530
rect 33846 27468 34110 27478
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 33846 27402 34110 27412
rect 33516 27022 33518 27074
rect 33570 27022 33572 27074
rect 33516 27010 33572 27022
rect 34076 27074 34132 27086
rect 34076 27022 34078 27074
rect 34130 27022 34132 27074
rect 33404 25454 33406 25506
rect 33458 25454 33460 25506
rect 33404 25442 33460 25454
rect 33628 26514 33684 26526
rect 33628 26462 33630 26514
rect 33682 26462 33684 26514
rect 33628 25508 33684 26462
rect 34076 26292 34132 27022
rect 34188 26740 34244 28478
rect 34300 27972 34356 28700
rect 34412 28196 34468 30830
rect 34412 28130 34468 28140
rect 34300 27916 34580 27972
rect 34300 27748 34356 27758
rect 34300 27746 34468 27748
rect 34300 27694 34302 27746
rect 34354 27694 34468 27746
rect 34300 27692 34468 27694
rect 34300 27682 34356 27692
rect 34188 26674 34244 26684
rect 34076 26226 34132 26236
rect 33846 25900 34110 25910
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 33846 25834 34110 25844
rect 33628 25452 34020 25508
rect 33852 25284 33908 25294
rect 33180 24782 33182 24834
rect 33234 24782 33236 24834
rect 33180 24770 33236 24782
rect 33628 25228 33852 25284
rect 31836 24722 31948 24724
rect 31836 24670 31838 24722
rect 31890 24670 31948 24722
rect 31836 24668 31948 24670
rect 31836 24658 31892 24668
rect 31948 24630 32004 24668
rect 33404 24724 33460 24734
rect 30380 24610 30436 24622
rect 30380 24558 30382 24610
rect 30434 24558 30436 24610
rect 30156 24050 30212 24062
rect 30156 23998 30158 24050
rect 30210 23998 30212 24050
rect 27244 23828 27300 23838
rect 27244 23734 27300 23772
rect 27580 23826 27636 23884
rect 28252 23940 28308 23978
rect 28252 23874 28308 23884
rect 27580 23774 27582 23826
rect 27634 23774 27636 23826
rect 27020 23716 27076 23726
rect 27020 23622 27076 23660
rect 26908 22990 26910 23042
rect 26962 22990 26964 23042
rect 25788 22820 25844 22830
rect 24522 22764 24786 22774
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24522 22698 24786 22708
rect 21812 22316 21924 22372
rect 22204 22484 22260 22494
rect 22204 22370 22260 22428
rect 22204 22318 22206 22370
rect 22258 22318 22260 22370
rect 21756 22278 21812 22316
rect 22204 22306 22260 22318
rect 22764 22260 22820 22270
rect 22764 21810 22820 22204
rect 22764 21758 22766 21810
rect 22818 21758 22820 21810
rect 22764 21746 22820 21758
rect 23772 22148 23828 22158
rect 21980 21700 22036 21710
rect 21532 20178 21588 20188
rect 21644 21698 22036 21700
rect 21644 21646 21982 21698
rect 22034 21646 22036 21698
rect 21644 21644 22036 21646
rect 21308 20078 21310 20130
rect 21362 20078 21364 20130
rect 21308 20066 21364 20078
rect 21644 20130 21700 21644
rect 21980 21634 22036 21644
rect 21756 21476 21812 21486
rect 21756 20914 21812 21420
rect 21756 20862 21758 20914
rect 21810 20862 21812 20914
rect 21756 20850 21812 20862
rect 22316 20802 22372 20814
rect 23772 20804 23828 22092
rect 24556 22146 24612 22158
rect 24556 22094 24558 22146
rect 24610 22094 24612 22146
rect 24556 21810 24612 22094
rect 24556 21758 24558 21810
rect 24610 21758 24612 21810
rect 24556 21746 24612 21758
rect 25228 22146 25284 22158
rect 25228 22094 25230 22146
rect 25282 22094 25284 22146
rect 24668 21476 24724 21486
rect 24668 21382 24724 21420
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20580 22372 20750
rect 23100 20748 23828 20804
rect 22316 20514 22372 20524
rect 22988 20580 23044 20590
rect 21644 20078 21646 20130
rect 21698 20078 21700 20130
rect 21644 20066 21700 20078
rect 22092 19908 22148 19918
rect 20972 19796 21028 19806
rect 19516 19346 19684 19348
rect 19516 19294 19518 19346
rect 19570 19294 19684 19346
rect 19516 19292 19684 19294
rect 20636 19794 21028 19796
rect 20636 19742 20974 19794
rect 21026 19742 21028 19794
rect 20636 19740 21028 19742
rect 17724 19282 17780 19292
rect 19516 19282 19572 19292
rect 17052 19234 17332 19236
rect 17052 19182 17054 19234
rect 17106 19182 17332 19234
rect 17052 19180 17332 19182
rect 17052 18452 17108 19180
rect 17388 19122 17444 19134
rect 17388 19070 17390 19122
rect 17442 19070 17444 19122
rect 17388 19012 17444 19070
rect 20636 19122 20692 19740
rect 20972 19730 21028 19740
rect 22092 19234 22148 19852
rect 22092 19182 22094 19234
rect 22146 19182 22148 19234
rect 22092 19170 22148 19182
rect 22988 19236 23044 20524
rect 23100 20188 23156 20748
rect 23436 20578 23492 20590
rect 23436 20526 23438 20578
rect 23490 20526 23492 20578
rect 23436 20188 23492 20526
rect 23100 20132 23380 20188
rect 23324 20020 23380 20132
rect 23436 20122 23492 20132
rect 23324 19964 23716 20020
rect 23212 19908 23268 19918
rect 23212 19814 23268 19852
rect 22988 19170 23044 19180
rect 20636 19070 20638 19122
rect 20690 19070 20692 19122
rect 20636 19058 20692 19070
rect 17388 18946 17444 18956
rect 19860 18844 20124 18854
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 19860 18778 20124 18788
rect 21868 18564 21924 18574
rect 21756 18562 21924 18564
rect 21756 18510 21870 18562
rect 21922 18510 21924 18562
rect 21756 18508 21924 18510
rect 17052 18386 17108 18396
rect 18956 18452 19012 18462
rect 19516 18452 19572 18462
rect 18956 18358 19012 18396
rect 19180 18450 19572 18452
rect 19180 18398 19518 18450
rect 19570 18398 19572 18450
rect 19180 18396 19572 18398
rect 17612 18340 17668 18350
rect 17612 18246 17668 18284
rect 18060 18340 18116 18350
rect 18060 18246 18116 18284
rect 16940 17826 16996 17836
rect 17948 17892 18004 17902
rect 17948 17554 18004 17836
rect 17948 17502 17950 17554
rect 18002 17502 18004 17554
rect 17948 17490 18004 17502
rect 16380 16380 16884 16436
rect 17052 17442 17108 17454
rect 17052 17390 17054 17442
rect 17106 17390 17108 17442
rect 17052 16436 17108 17390
rect 17164 17444 17220 17454
rect 17164 17442 17892 17444
rect 17164 17390 17166 17442
rect 17218 17390 17892 17442
rect 17164 17388 17892 17390
rect 17164 17378 17220 17388
rect 17836 16994 17892 17388
rect 17836 16942 17838 16994
rect 17890 16942 17892 16994
rect 17836 16930 17892 16942
rect 19180 16770 19236 18396
rect 19516 18386 19572 18396
rect 20636 18340 20692 18350
rect 19180 16718 19182 16770
rect 19234 16718 19236 16770
rect 19180 16706 19236 16718
rect 19404 17668 19460 17678
rect 17052 16380 17220 16436
rect 16380 16100 16436 16380
rect 16380 16006 16436 16044
rect 16604 15540 16660 16380
rect 16716 16268 17108 16324
rect 16716 16098 16772 16268
rect 16716 16046 16718 16098
rect 16770 16046 16772 16098
rect 16716 16034 16772 16046
rect 16716 15540 16772 15550
rect 16604 15538 16884 15540
rect 16604 15486 16718 15538
rect 16770 15486 16884 15538
rect 16604 15484 16884 15486
rect 16716 15474 16772 15484
rect 16044 15222 16100 15260
rect 16268 15202 16324 15214
rect 16268 15150 16270 15202
rect 16322 15150 16324 15202
rect 16268 12850 16324 15150
rect 16380 15204 16436 15214
rect 16380 13970 16436 15148
rect 16380 13918 16382 13970
rect 16434 13918 16436 13970
rect 16380 13906 16436 13918
rect 16828 14644 16884 15484
rect 16268 12798 16270 12850
rect 16322 12798 16324 12850
rect 16268 12786 16324 12798
rect 16380 12402 16436 12414
rect 16380 12350 16382 12402
rect 16434 12350 16436 12402
rect 16380 12292 16436 12350
rect 16380 12226 16436 12236
rect 15372 11506 15652 11508
rect 15372 11454 15374 11506
rect 15426 11454 15652 11506
rect 15372 11452 15652 11454
rect 15708 11620 15764 11630
rect 15372 11442 15428 11452
rect 14364 11230 14366 11282
rect 14418 11230 14420 11282
rect 14364 11218 14420 11230
rect 14028 9874 14084 9884
rect 14924 10612 14980 10622
rect 14812 9716 14868 9726
rect 12796 9662 12798 9714
rect 12850 9662 12852 9714
rect 12796 9650 12852 9662
rect 14140 9714 14868 9716
rect 14140 9662 14814 9714
rect 14866 9662 14868 9714
rect 14140 9660 14868 9662
rect 14140 9266 14196 9660
rect 14812 9650 14868 9660
rect 14140 9214 14142 9266
rect 14194 9214 14196 9266
rect 14140 9202 14196 9214
rect 14364 9380 14420 9390
rect 12460 8094 12462 8146
rect 12514 8094 12516 8146
rect 12460 8082 12516 8094
rect 14364 7586 14420 9324
rect 14924 9044 14980 10556
rect 15596 10500 15652 10510
rect 15198 10220 15462 10230
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15198 10154 15462 10164
rect 15148 9940 15204 9950
rect 15596 9940 15652 10444
rect 15148 9938 15652 9940
rect 15148 9886 15150 9938
rect 15202 9886 15652 9938
rect 15148 9884 15652 9886
rect 15148 9874 15204 9884
rect 15708 9714 15764 11564
rect 15932 11508 15988 11518
rect 16380 11508 16436 11518
rect 16828 11508 16884 14588
rect 16940 13522 16996 13534
rect 16940 13470 16942 13522
rect 16994 13470 16996 13522
rect 16940 12180 16996 13470
rect 17052 12964 17108 16268
rect 17164 14868 17220 16380
rect 18956 16212 19012 16222
rect 18956 15538 19012 16156
rect 19292 15988 19348 15998
rect 19292 15874 19348 15932
rect 19292 15822 19294 15874
rect 19346 15822 19348 15874
rect 19292 15810 19348 15822
rect 18956 15486 18958 15538
rect 19010 15486 19012 15538
rect 18956 15474 19012 15486
rect 17836 15316 17892 15326
rect 17500 15204 17556 15214
rect 17500 15110 17556 15148
rect 17836 15202 17892 15260
rect 17836 15150 17838 15202
rect 17890 15150 17892 15202
rect 17164 14802 17220 14812
rect 17276 14644 17332 14654
rect 17276 13746 17332 14588
rect 17276 13694 17278 13746
rect 17330 13694 17332 13746
rect 17276 13682 17332 13694
rect 17052 12898 17108 12908
rect 16940 12114 16996 12124
rect 17052 12738 17108 12750
rect 17052 12686 17054 12738
rect 17106 12686 17108 12738
rect 16940 11954 16996 11966
rect 16940 11902 16942 11954
rect 16994 11902 16996 11954
rect 16940 11620 16996 11902
rect 17052 11620 17108 12686
rect 17164 12740 17220 12750
rect 17164 12738 17444 12740
rect 17164 12686 17166 12738
rect 17218 12686 17444 12738
rect 17164 12684 17444 12686
rect 17164 12674 17220 12684
rect 17052 11564 17332 11620
rect 16940 11554 16996 11564
rect 15932 11506 16884 11508
rect 15932 11454 15934 11506
rect 15986 11454 16382 11506
rect 16434 11454 16884 11506
rect 15932 11452 16884 11454
rect 15932 11442 15988 11452
rect 16380 11442 16436 11452
rect 16156 10610 16212 10622
rect 16156 10558 16158 10610
rect 16210 10558 16212 10610
rect 15708 9662 15710 9714
rect 15762 9662 15764 9714
rect 15708 9650 15764 9662
rect 15932 10388 15988 10398
rect 15036 9044 15092 9054
rect 14924 8988 15036 9044
rect 15036 8950 15092 8988
rect 14364 7534 14366 7586
rect 14418 7534 14420 7586
rect 14364 7522 14420 7534
rect 14700 8818 14756 8830
rect 14700 8766 14702 8818
rect 14754 8766 14756 8818
rect 14700 7476 14756 8766
rect 15198 8652 15462 8662
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15198 8586 15462 8596
rect 15932 8370 15988 10332
rect 16156 8428 16212 10558
rect 16492 10612 16548 11452
rect 16828 11394 16884 11452
rect 17164 11396 17220 11406
rect 16828 11342 16830 11394
rect 16882 11342 16884 11394
rect 16828 11330 16884 11342
rect 16940 11394 17220 11396
rect 16940 11342 17166 11394
rect 17218 11342 17220 11394
rect 16940 11340 17220 11342
rect 16492 10518 16548 10556
rect 16940 9938 16996 11340
rect 17164 11330 17220 11340
rect 16940 9886 16942 9938
rect 16994 9886 16996 9938
rect 16940 9874 16996 9886
rect 17276 8428 17332 11564
rect 17388 10948 17444 12684
rect 17724 12292 17780 12302
rect 17724 12198 17780 12236
rect 17836 12068 17892 15150
rect 18172 15090 18228 15102
rect 18172 15038 18174 15090
rect 18226 15038 18228 15090
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13076 18004 13694
rect 17948 13010 18004 13020
rect 17948 12852 18004 12862
rect 17948 12758 18004 12796
rect 17948 12178 18004 12190
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17948 12068 18004 12126
rect 17388 10882 17444 10892
rect 17612 12012 17948 12068
rect 17388 10724 17444 10734
rect 17388 10630 17444 10668
rect 17612 10610 17668 12012
rect 17948 11974 18004 12012
rect 18172 11396 18228 15038
rect 19292 14644 19348 14654
rect 18620 13076 18676 13086
rect 18284 12964 18340 12974
rect 18284 11732 18340 12908
rect 18284 11676 18452 11732
rect 18172 11340 18340 11396
rect 18172 11172 18228 11182
rect 18172 10836 18228 11116
rect 17612 10558 17614 10610
rect 17666 10558 17668 10610
rect 17612 10500 17668 10558
rect 17612 10434 17668 10444
rect 17836 10834 18228 10836
rect 17836 10782 18174 10834
rect 18226 10782 18228 10834
rect 17836 10780 18228 10782
rect 17388 9940 17444 9950
rect 17836 9940 17892 10780
rect 18172 10770 18228 10780
rect 18284 10724 18340 11340
rect 18284 10658 18340 10668
rect 17388 9938 17892 9940
rect 17388 9886 17390 9938
rect 17442 9886 17838 9938
rect 17890 9886 17892 9938
rect 17388 9884 17892 9886
rect 17388 9874 17444 9884
rect 17836 9874 17892 9884
rect 18396 8930 18452 11676
rect 18396 8878 18398 8930
rect 18450 8878 18452 8930
rect 18396 8866 18452 8878
rect 16156 8372 16884 8428
rect 15932 8318 15934 8370
rect 15986 8318 15988 8370
rect 15932 8306 15988 8318
rect 14700 7410 14756 7420
rect 15708 7476 15764 7486
rect 13356 7364 13412 7374
rect 13356 7270 13412 7308
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 12012 6526 12014 6578
rect 12066 6526 12068 6578
rect 12012 6514 12068 6526
rect 15708 6578 15764 7420
rect 16828 6802 16884 8372
rect 17164 8372 17332 8428
rect 18620 8428 18676 13020
rect 18844 12180 18900 12190
rect 18900 12124 19012 12180
rect 18844 12114 18900 12124
rect 18732 12068 18788 12078
rect 18732 11974 18788 12012
rect 18956 10276 19012 12124
rect 19292 12178 19348 14588
rect 19292 12126 19294 12178
rect 19346 12126 19348 12178
rect 19068 12066 19124 12078
rect 19068 12014 19070 12066
rect 19122 12014 19124 12066
rect 19068 11620 19124 12014
rect 19068 11554 19124 11564
rect 19292 11284 19348 12126
rect 19292 11218 19348 11228
rect 19404 10498 19460 17612
rect 20188 17668 20244 17678
rect 20188 17574 20244 17612
rect 20636 17666 20692 18284
rect 21756 17778 21812 18508
rect 21868 18498 21924 18508
rect 22876 18338 22932 18350
rect 22876 18286 22878 18338
rect 22930 18286 22932 18338
rect 21756 17726 21758 17778
rect 21810 17726 21812 17778
rect 21756 17714 21812 17726
rect 22652 18226 22708 18238
rect 22652 18174 22654 18226
rect 22706 18174 22708 18226
rect 20636 17614 20638 17666
rect 20690 17614 20692 17666
rect 20636 17602 20692 17614
rect 22204 17666 22260 17678
rect 22204 17614 22206 17666
rect 22258 17614 22260 17666
rect 21980 17554 22036 17566
rect 21980 17502 21982 17554
rect 22034 17502 22036 17554
rect 19860 17276 20124 17286
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 19860 17210 20124 17220
rect 21980 17220 22036 17502
rect 20636 16884 20692 16894
rect 20636 16790 20692 16828
rect 21084 16882 21140 16894
rect 21084 16830 21086 16882
rect 21138 16830 21140 16882
rect 21084 16100 21140 16830
rect 21084 16034 21140 16044
rect 21532 16884 21588 16894
rect 20076 15988 20132 15998
rect 20076 15894 20132 15932
rect 20412 15986 20468 15998
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 19852 15876 19908 15886
rect 19628 15874 19908 15876
rect 19628 15822 19854 15874
rect 19906 15822 19908 15874
rect 19628 15820 19908 15822
rect 19516 15204 19572 15214
rect 19516 14642 19572 15148
rect 19516 14590 19518 14642
rect 19570 14590 19572 14642
rect 19516 14532 19572 14590
rect 19516 14466 19572 14476
rect 19516 11620 19572 11630
rect 19516 11282 19572 11564
rect 19516 11230 19518 11282
rect 19570 11230 19572 11282
rect 19516 11218 19572 11230
rect 19628 11284 19684 15820
rect 19852 15810 19908 15820
rect 19860 15708 20124 15718
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 19860 15642 20124 15652
rect 20412 15316 20468 15934
rect 20412 15250 20468 15260
rect 21308 15314 21364 15326
rect 21308 15262 21310 15314
rect 21362 15262 21364 15314
rect 19964 14644 20020 14654
rect 19964 14550 20020 14588
rect 20748 14308 20804 14318
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 20412 13970 20468 13982
rect 20412 13918 20414 13970
rect 20466 13918 20468 13970
rect 20412 13300 20468 13918
rect 20412 13234 20468 13244
rect 20188 12962 20244 12974
rect 20188 12910 20190 12962
rect 20242 12910 20244 12962
rect 19860 12572 20124 12582
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 19860 12506 20124 12516
rect 19964 12180 20020 12190
rect 19628 11218 19684 11228
rect 19740 12178 20020 12180
rect 19740 12126 19966 12178
rect 20018 12126 20020 12178
rect 19740 12124 20020 12126
rect 19404 10446 19406 10498
rect 19458 10446 19460 10498
rect 19404 10434 19460 10446
rect 19628 10948 19684 10958
rect 18956 10220 19460 10276
rect 19292 9940 19348 9950
rect 19292 9846 19348 9884
rect 19404 9154 19460 10220
rect 19404 9102 19406 9154
rect 19458 9102 19460 9154
rect 19404 9090 19460 9102
rect 19628 8428 19684 10892
rect 19740 10500 19796 12124
rect 19964 12114 20020 12124
rect 20188 11508 20244 12910
rect 20188 11442 20244 11452
rect 20300 11170 20356 11182
rect 20300 11118 20302 11170
rect 20354 11118 20356 11170
rect 19860 11004 20124 11014
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 19860 10938 20124 10948
rect 20188 10724 20244 10734
rect 20188 10630 20244 10668
rect 19740 10434 19796 10444
rect 20300 10052 20356 11118
rect 20636 11172 20692 11182
rect 20636 11078 20692 11116
rect 20300 9986 20356 9996
rect 20636 9716 20692 9726
rect 20748 9716 20804 14252
rect 21308 13972 21364 15262
rect 21308 13906 21364 13916
rect 21532 15316 21588 16828
rect 21644 16212 21700 16222
rect 21644 16118 21700 16156
rect 21980 16210 22036 17164
rect 22204 16884 22260 17614
rect 22204 16818 22260 16828
rect 21980 16158 21982 16210
rect 22034 16158 22036 16210
rect 21980 16146 22036 16158
rect 22652 15428 22708 18174
rect 22876 17892 22932 18286
rect 23212 18340 23268 18350
rect 23212 18246 23268 18284
rect 23548 18338 23604 18350
rect 23548 18286 23550 18338
rect 23602 18286 23604 18338
rect 22876 17826 22932 17836
rect 22876 17666 22932 17678
rect 22876 17614 22878 17666
rect 22930 17614 22932 17666
rect 22876 17108 22932 17614
rect 22876 17042 22932 17052
rect 23548 17106 23604 18286
rect 23548 17054 23550 17106
rect 23602 17054 23604 17106
rect 23548 17042 23604 17054
rect 23436 16772 23492 16782
rect 23436 16322 23492 16716
rect 23436 16270 23438 16322
rect 23490 16270 23492 16322
rect 23436 16258 23492 16270
rect 23100 16100 23156 16110
rect 22764 15540 22820 15550
rect 22764 15446 22820 15484
rect 22652 15362 22708 15372
rect 21644 15316 21700 15326
rect 21532 15314 21700 15316
rect 21532 15262 21646 15314
rect 21698 15262 21700 15314
rect 21532 15260 21700 15262
rect 21084 13748 21140 13758
rect 21532 13748 21588 15260
rect 21644 15250 21700 15260
rect 23100 15202 23156 16044
rect 23660 15540 23716 19964
rect 23660 15474 23716 15484
rect 23772 19122 23828 20748
rect 24220 20580 24276 20590
rect 24220 20486 24276 20524
rect 25228 20188 25284 22094
rect 25564 22148 25620 22158
rect 25564 22054 25620 22092
rect 25340 21588 25396 21598
rect 25340 21494 25396 21532
rect 25788 21586 25844 22764
rect 26460 22484 26516 22494
rect 26460 22390 26516 22428
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25788 21522 25844 21534
rect 26908 21588 26964 22990
rect 27468 22260 27524 22270
rect 27468 22166 27524 22204
rect 26572 20802 26628 20814
rect 26572 20750 26574 20802
rect 26626 20750 26628 20802
rect 24220 20132 24276 20142
rect 25228 20132 26292 20188
rect 24220 20038 24276 20076
rect 26012 19796 26068 19806
rect 26012 19702 26068 19740
rect 24522 19628 24786 19638
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24522 19562 24786 19572
rect 23772 19070 23774 19122
rect 23826 19070 23828 19122
rect 23100 15150 23102 15202
rect 23154 15150 23156 15202
rect 23100 15138 23156 15150
rect 23772 15204 23828 19070
rect 23884 18340 23940 18350
rect 23884 17220 23940 18284
rect 24522 18060 24786 18070
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24522 17994 24786 18004
rect 26236 17554 26292 20132
rect 26572 19012 26628 20750
rect 26908 20802 26964 21532
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26908 20738 26964 20750
rect 27580 21476 27636 23774
rect 28252 23714 28308 23726
rect 28252 23662 28254 23714
rect 28306 23662 28308 23714
rect 28252 21810 28308 23662
rect 29184 23548 29448 23558
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29184 23482 29448 23492
rect 28364 23380 28420 23390
rect 28364 22482 28420 23324
rect 29372 23154 29428 23166
rect 29372 23102 29374 23154
rect 29426 23102 29428 23154
rect 28364 22430 28366 22482
rect 28418 22430 28420 22482
rect 28364 22418 28420 22430
rect 28812 22932 28868 22942
rect 28588 22372 28644 22382
rect 28588 22260 28644 22316
rect 28252 21758 28254 21810
rect 28306 21758 28308 21810
rect 28252 21746 28308 21758
rect 28476 22258 28644 22260
rect 28476 22206 28590 22258
rect 28642 22206 28644 22258
rect 28476 22204 28644 22206
rect 27580 20802 27636 21420
rect 28476 21476 28532 22204
rect 28588 22194 28644 22204
rect 28812 21810 28868 22876
rect 29260 22370 29316 22382
rect 29260 22318 29262 22370
rect 29314 22318 29316 22370
rect 29260 22260 29316 22318
rect 29260 22194 29316 22204
rect 29372 22148 29428 23102
rect 30156 22820 30212 23998
rect 30380 23940 30436 24558
rect 32956 24052 33012 24062
rect 32956 23958 33012 23996
rect 30380 23874 30436 23884
rect 31164 23826 31220 23838
rect 31164 23774 31166 23826
rect 31218 23774 31220 23826
rect 31164 23716 31220 23774
rect 31164 23650 31220 23660
rect 33180 23156 33236 23166
rect 30156 22754 30212 22764
rect 31388 23042 31444 23054
rect 31388 22990 31390 23042
rect 31442 22990 31444 23042
rect 29708 22482 29764 22494
rect 29708 22430 29710 22482
rect 29762 22430 29764 22482
rect 29484 22372 29540 22382
rect 29708 22372 29764 22430
rect 29540 22316 29764 22372
rect 31164 22372 31220 22382
rect 31388 22372 31444 22990
rect 31164 22370 31444 22372
rect 31164 22318 31166 22370
rect 31218 22318 31444 22370
rect 31164 22316 31444 22318
rect 33180 22482 33236 23100
rect 33180 22430 33182 22482
rect 33234 22430 33236 22482
rect 29484 22306 29540 22316
rect 29372 22082 29428 22092
rect 29820 22260 29876 22270
rect 29184 21980 29448 21990
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29184 21914 29448 21924
rect 28812 21758 28814 21810
rect 28866 21758 28868 21810
rect 28812 21746 28868 21758
rect 28476 21410 28532 21420
rect 28924 21586 28980 21598
rect 28924 21534 28926 21586
rect 28978 21534 28980 21586
rect 27580 20750 27582 20802
rect 27634 20750 27636 20802
rect 27580 20738 27636 20750
rect 28924 20804 28980 21534
rect 29596 21588 29652 21598
rect 29596 21494 29652 21532
rect 26796 20692 26852 20702
rect 26796 20130 26852 20636
rect 27356 20690 27412 20702
rect 27356 20638 27358 20690
rect 27410 20638 27412 20690
rect 27356 20580 27412 20638
rect 28252 20692 28308 20702
rect 28252 20598 28308 20636
rect 28588 20692 28644 20702
rect 27356 20514 27412 20524
rect 28588 20188 28644 20636
rect 26796 20078 26798 20130
rect 26850 20078 26852 20130
rect 26796 20066 26852 20078
rect 28364 20132 28644 20188
rect 28924 20188 28980 20748
rect 29820 20802 29876 22204
rect 30828 22260 30884 22270
rect 30828 22166 30884 22204
rect 31164 22148 31220 22316
rect 31164 22082 31220 22092
rect 32060 21810 32116 21822
rect 32060 21758 32062 21810
rect 32114 21758 32116 21810
rect 32060 21700 32116 21758
rect 32060 21634 32116 21644
rect 33068 21700 33124 21710
rect 33068 21606 33124 21644
rect 31724 21476 31780 21486
rect 29820 20750 29822 20802
rect 29874 20750 29876 20802
rect 29184 20412 29448 20422
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29184 20346 29448 20356
rect 28924 20132 29540 20188
rect 26572 18946 26628 18956
rect 26908 19908 26964 19918
rect 26460 18900 26516 18910
rect 26236 17502 26238 17554
rect 26290 17502 26292 17554
rect 26236 17490 26292 17502
rect 26348 18450 26404 18462
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 25228 17442 25284 17454
rect 25228 17390 25230 17442
rect 25282 17390 25284 17442
rect 23884 17154 23940 17164
rect 24668 17220 24724 17230
rect 24108 16996 24164 17006
rect 24108 16902 24164 16940
rect 24668 16994 24724 17164
rect 24668 16942 24670 16994
rect 24722 16942 24724 16994
rect 24668 16930 24724 16942
rect 25228 16994 25284 17390
rect 25900 17444 25956 17454
rect 25900 17442 26180 17444
rect 25900 17390 25902 17442
rect 25954 17390 26180 17442
rect 25900 17388 26180 17390
rect 25900 17378 25956 17388
rect 25228 16942 25230 16994
rect 25282 16942 25284 16994
rect 25228 16930 25284 16942
rect 25564 17220 25620 17230
rect 25564 16994 25620 17164
rect 25564 16942 25566 16994
rect 25618 16942 25620 16994
rect 25564 16930 25620 16942
rect 26012 16884 26068 16894
rect 25788 16828 26012 16884
rect 24332 16770 24388 16782
rect 24332 16718 24334 16770
rect 24386 16718 24388 16770
rect 24220 15876 24276 15886
rect 24220 15782 24276 15820
rect 24108 15428 24164 15438
rect 24108 15334 24164 15372
rect 23772 15138 23828 15148
rect 23660 14308 23716 14318
rect 23660 14214 23716 14252
rect 24332 14306 24388 16718
rect 24522 16492 24786 16502
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24522 16426 24786 16436
rect 25788 15202 25844 16828
rect 26012 16790 26068 16828
rect 25788 15150 25790 15202
rect 25842 15150 25844 15202
rect 24522 14924 24786 14934
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24522 14858 24786 14868
rect 24332 14254 24334 14306
rect 24386 14254 24388 14306
rect 24332 14242 24388 14254
rect 22316 13972 22372 13982
rect 21084 13746 21588 13748
rect 21084 13694 21086 13746
rect 21138 13694 21588 13746
rect 21084 13692 21588 13694
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 20972 13522 21028 13534
rect 20972 13470 20974 13522
rect 21026 13470 21028 13522
rect 20972 13188 21028 13470
rect 20972 13122 21028 13132
rect 20860 12964 20916 12974
rect 21084 12964 21140 13692
rect 20860 12962 21084 12964
rect 20860 12910 20862 12962
rect 20914 12910 21084 12962
rect 20860 12908 21084 12910
rect 20860 12898 20916 12908
rect 21084 12870 21140 12908
rect 21532 12852 21588 12862
rect 21532 12292 21588 12796
rect 21756 12628 21812 13694
rect 22204 13076 22260 13086
rect 22204 12982 22260 13020
rect 21868 12852 21924 12862
rect 21868 12850 22260 12852
rect 21868 12798 21870 12850
rect 21922 12798 22260 12850
rect 21868 12796 22260 12798
rect 21868 12786 21924 12796
rect 21756 12562 21812 12572
rect 22204 12402 22260 12796
rect 22204 12350 22206 12402
rect 22258 12350 22260 12402
rect 22204 12338 22260 12350
rect 21532 12226 21588 12236
rect 22316 11506 22372 13916
rect 24220 13970 24276 13982
rect 24220 13918 24222 13970
rect 24274 13918 24276 13970
rect 23212 13524 23268 13534
rect 22876 13188 22932 13198
rect 22428 12962 22484 12974
rect 22428 12910 22430 12962
rect 22482 12910 22484 12962
rect 22428 12852 22484 12910
rect 22428 12786 22484 12796
rect 22316 11454 22318 11506
rect 22370 11454 22372 11506
rect 22316 11442 22372 11454
rect 22428 11508 22484 11518
rect 21980 10500 22036 10510
rect 21980 10406 22036 10444
rect 22428 9938 22484 11452
rect 22876 10724 22932 13132
rect 23212 12964 23268 13468
rect 23324 13300 23380 13310
rect 23380 13244 23492 13300
rect 23324 13234 23380 13244
rect 23212 12870 23268 12908
rect 23324 12852 23380 12862
rect 23324 12178 23380 12796
rect 23324 12126 23326 12178
rect 23378 12126 23380 12178
rect 23324 12114 23380 12126
rect 23436 12066 23492 13244
rect 23436 12014 23438 12066
rect 23490 12014 23492 12066
rect 23436 12002 23492 12014
rect 23884 12962 23940 12974
rect 23884 12910 23886 12962
rect 23938 12910 23940 12962
rect 22988 11954 23044 11966
rect 22988 11902 22990 11954
rect 23042 11902 23044 11954
rect 22988 11620 23044 11902
rect 22988 11554 23044 11564
rect 23548 11284 23604 11294
rect 23548 11190 23604 11228
rect 22988 10724 23044 10734
rect 22876 10722 23044 10724
rect 22876 10670 22990 10722
rect 23042 10670 23044 10722
rect 22876 10668 23044 10670
rect 22988 10658 23044 10668
rect 23884 10500 23940 12910
rect 24220 12290 24276 13918
rect 25228 13746 25284 13758
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 24780 13524 24836 13534
rect 25228 13524 25284 13694
rect 24780 13522 24948 13524
rect 24780 13470 24782 13522
rect 24834 13470 24948 13522
rect 24780 13468 24948 13470
rect 24780 13458 24836 13468
rect 24522 13356 24786 13366
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24522 13290 24786 13300
rect 24220 12238 24222 12290
rect 24274 12238 24276 12290
rect 24220 12226 24276 12238
rect 24556 12292 24612 12302
rect 24556 12198 24612 12236
rect 24892 12068 24948 13468
rect 25228 13458 25284 13468
rect 25676 13746 25732 13758
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 24892 12002 24948 12012
rect 25116 12628 25172 12638
rect 24522 11788 24786 11798
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24522 11722 24786 11732
rect 25116 11506 25172 12572
rect 25564 12292 25620 12302
rect 25676 12292 25732 13694
rect 25788 13524 25844 15150
rect 25788 13458 25844 13468
rect 26124 13412 26180 17388
rect 26348 16884 26404 18398
rect 26348 16818 26404 16828
rect 26460 13748 26516 18844
rect 26908 18450 26964 19852
rect 27916 19236 27972 19246
rect 27916 19142 27972 19180
rect 26908 18398 26910 18450
rect 26962 18398 26964 18450
rect 26908 18386 26964 18398
rect 27356 19012 27412 19022
rect 27356 17778 27412 18956
rect 27356 17726 27358 17778
rect 27410 17726 27412 17778
rect 27356 17714 27412 17726
rect 27580 19010 27636 19022
rect 27580 18958 27582 19010
rect 27634 18958 27636 19010
rect 27580 17220 27636 18958
rect 26572 16882 26628 16894
rect 26572 16830 26574 16882
rect 26626 16830 26628 16882
rect 26572 16324 26628 16830
rect 26684 16884 26740 16894
rect 26740 16828 26852 16884
rect 26684 16818 26740 16828
rect 26796 16772 26852 16828
rect 26796 16716 26964 16772
rect 26572 16268 26740 16324
rect 26572 16098 26628 16110
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 14084 26628 16046
rect 26572 14018 26628 14028
rect 26124 13346 26180 13356
rect 26348 13692 26516 13748
rect 26124 12740 26180 12750
rect 26012 12738 26180 12740
rect 26012 12686 26126 12738
rect 26178 12686 26180 12738
rect 26012 12684 26180 12686
rect 25676 12236 25844 12292
rect 25564 12068 25620 12236
rect 25788 12180 25844 12236
rect 26012 12290 26068 12684
rect 26124 12674 26180 12684
rect 26012 12238 26014 12290
rect 26066 12238 26068 12290
rect 26012 12226 26068 12238
rect 25788 12114 25844 12124
rect 25676 12068 25732 12078
rect 25564 12066 25732 12068
rect 25564 12014 25678 12066
rect 25730 12014 25732 12066
rect 25564 12012 25732 12014
rect 25676 12002 25732 12012
rect 25116 11454 25118 11506
rect 25170 11454 25172 11506
rect 25116 11442 25172 11454
rect 26124 11620 26180 11630
rect 26124 11282 26180 11564
rect 26124 11230 26126 11282
rect 26178 11230 26180 11282
rect 26124 11218 26180 11230
rect 23884 10434 23940 10444
rect 26236 10500 26292 10510
rect 26236 10406 26292 10444
rect 24522 10220 24786 10230
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24522 10154 24786 10164
rect 22428 9886 22430 9938
rect 22482 9886 22484 9938
rect 22428 9874 22484 9886
rect 23548 10052 23604 10062
rect 20636 9714 20804 9716
rect 20636 9662 20638 9714
rect 20690 9662 20804 9714
rect 20636 9660 20804 9662
rect 23548 9714 23604 9996
rect 23548 9662 23550 9714
rect 23602 9662 23604 9714
rect 20636 9650 20692 9660
rect 23548 9650 23604 9662
rect 19860 9436 20124 9446
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 19860 9370 20124 9380
rect 24522 8652 24786 8662
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24522 8586 24786 8596
rect 18620 8372 18788 8428
rect 19628 8372 19796 8428
rect 17164 8146 17220 8372
rect 18732 8370 18788 8372
rect 18732 8318 18734 8370
rect 18786 8318 18788 8370
rect 18732 8306 18788 8318
rect 17164 8094 17166 8146
rect 17218 8094 17220 8146
rect 17164 8082 17220 8094
rect 19740 8146 19796 8372
rect 21980 8260 22036 8270
rect 21980 8258 22148 8260
rect 21980 8206 21982 8258
rect 22034 8206 22148 8258
rect 21980 8204 22148 8206
rect 21980 8194 22036 8204
rect 19740 8094 19742 8146
rect 19794 8094 19796 8146
rect 19740 8082 19796 8094
rect 19860 7868 20124 7878
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 19860 7802 20124 7812
rect 16828 6750 16830 6802
rect 16882 6750 16884 6802
rect 16828 6738 16884 6750
rect 15708 6526 15710 6578
rect 15762 6526 15764 6578
rect 15708 6514 15764 6526
rect 19860 6300 20124 6310
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 19860 6234 20124 6244
rect 11788 5966 11790 6018
rect 11842 5966 11844 6018
rect 11788 5954 11844 5966
rect 10556 5796 10612 5806
rect 10332 5794 10612 5796
rect 10332 5742 10558 5794
rect 10610 5742 10612 5794
rect 10332 5740 10612 5742
rect 10556 5730 10612 5740
rect 5874 5516 6138 5526
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 5874 5450 6138 5460
rect 15198 5516 15462 5526
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15198 5450 15462 5460
rect 10536 4732 10800 4742
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10536 4666 10800 4676
rect 19860 4732 20124 4742
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 19860 4666 20124 4676
rect 5874 3948 6138 3958
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 5874 3882 6138 3892
rect 15198 3948 15462 3958
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15198 3882 15462 3892
rect 21532 3444 21588 3454
rect 21756 3444 21812 3454
rect 21532 3442 21812 3444
rect 21532 3390 21534 3442
rect 21586 3390 21758 3442
rect 21810 3390 21812 3442
rect 21532 3388 21812 3390
rect 10536 3164 10800 3174
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10536 3098 10800 3108
rect 19860 3164 20124 3174
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 19860 3098 20124 3108
rect 21532 800 21588 3388
rect 21756 3378 21812 3388
rect 22092 3442 22148 8204
rect 22204 8036 22260 8046
rect 22204 8034 22484 8036
rect 22204 7982 22206 8034
rect 22258 7982 22484 8034
rect 22204 7980 22484 7982
rect 22204 7970 22260 7980
rect 22428 3554 22484 7980
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 26348 6580 26404 13692
rect 26684 13524 26740 16268
rect 26908 16100 26964 16716
rect 27580 16210 27636 17164
rect 27580 16158 27582 16210
rect 27634 16158 27636 16210
rect 26908 16098 27188 16100
rect 26908 16046 26910 16098
rect 26962 16046 27188 16098
rect 26908 16044 27188 16046
rect 26908 16034 26964 16044
rect 26684 13458 26740 13468
rect 26796 14530 26852 14542
rect 26796 14478 26798 14530
rect 26850 14478 26852 14530
rect 26348 6514 26404 6524
rect 26460 11620 26516 11630
rect 26460 6020 26516 11564
rect 26572 11172 26628 11182
rect 26572 9714 26628 11116
rect 26572 9662 26574 9714
rect 26626 9662 26628 9714
rect 26572 9650 26628 9662
rect 26796 8932 26852 14478
rect 27132 14530 27188 16044
rect 27132 14478 27134 14530
rect 27186 14478 27188 14530
rect 27132 14466 27188 14478
rect 27580 14418 27636 16158
rect 28252 18228 28308 18238
rect 27692 15876 27748 15886
rect 27692 15782 27748 15820
rect 27580 14366 27582 14418
rect 27634 14366 27636 14418
rect 27356 14084 27412 14094
rect 26908 12738 26964 12750
rect 26908 12686 26910 12738
rect 26962 12686 26964 12738
rect 26908 11732 26964 12686
rect 26908 11666 26964 11676
rect 27244 12068 27300 12078
rect 27244 10722 27300 12012
rect 27356 12066 27412 14028
rect 27580 12292 27636 14366
rect 27916 14420 27972 14430
rect 27916 14418 28084 14420
rect 27916 14366 27918 14418
rect 27970 14366 28084 14418
rect 27916 14364 28084 14366
rect 27916 14354 27972 14364
rect 28028 13970 28084 14364
rect 28028 13918 28030 13970
rect 28082 13918 28084 13970
rect 28028 13906 28084 13918
rect 27580 12226 27636 12236
rect 27356 12014 27358 12066
rect 27410 12014 27412 12066
rect 27356 12002 27412 12014
rect 27244 10670 27246 10722
rect 27298 10670 27300 10722
rect 27244 10658 27300 10670
rect 27580 11620 27636 11630
rect 27244 10500 27300 10510
rect 27132 10444 27244 10500
rect 26796 8866 26852 8876
rect 27020 10388 27076 10398
rect 27020 8428 27076 10332
rect 26572 8372 27076 8428
rect 26572 8146 26628 8372
rect 26572 8094 26574 8146
rect 26626 8094 26628 8146
rect 26572 8082 26628 8094
rect 27132 6916 27188 10444
rect 27244 10434 27300 10444
rect 27580 9938 27636 11564
rect 27580 9886 27582 9938
rect 27634 9886 27636 9938
rect 27580 9874 27636 9886
rect 28252 9716 28308 18172
rect 28364 16098 28420 20132
rect 29148 20020 29204 20030
rect 29148 19926 29204 19964
rect 29484 20018 29540 20132
rect 29484 19966 29486 20018
rect 29538 19966 29540 20018
rect 29484 19954 29540 19966
rect 29820 20132 29876 20750
rect 31052 20804 31108 20814
rect 31052 20710 31108 20748
rect 31612 20802 31668 20814
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 30380 20692 30436 20702
rect 30380 20598 30436 20636
rect 29820 19348 29876 20076
rect 30604 20132 30660 20142
rect 30604 20038 30660 20076
rect 30940 19908 30996 19918
rect 30940 19814 30996 19852
rect 29820 19282 29876 19292
rect 30380 19348 30436 19358
rect 28588 19236 28644 19246
rect 28588 19142 28644 19180
rect 29260 19236 29316 19246
rect 29260 19142 29316 19180
rect 29708 19234 29764 19246
rect 29708 19182 29710 19234
rect 29762 19182 29764 19234
rect 29184 18844 29448 18854
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29184 18778 29448 18788
rect 29148 18564 29204 18574
rect 28588 18562 29204 18564
rect 28588 18510 29150 18562
rect 29202 18510 29204 18562
rect 28588 18508 29204 18510
rect 28588 17220 28644 18508
rect 29148 18498 29204 18508
rect 28476 17164 28644 17220
rect 29036 17442 29092 17454
rect 29036 17390 29038 17442
rect 29090 17390 29092 17442
rect 28476 16210 28532 17164
rect 28924 16996 28980 17006
rect 28476 16158 28478 16210
rect 28530 16158 28532 16210
rect 28476 16146 28532 16158
rect 28588 16994 28980 16996
rect 28588 16942 28926 16994
rect 28978 16942 28980 16994
rect 28588 16940 28980 16942
rect 28364 16046 28366 16098
rect 28418 16046 28420 16098
rect 28364 14530 28420 16046
rect 28588 15652 28644 16940
rect 28924 16930 28980 16940
rect 28476 15596 28644 15652
rect 28476 14642 28532 15596
rect 29036 15316 29092 17390
rect 29184 17276 29448 17286
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29184 17210 29448 17220
rect 29708 16884 29764 19182
rect 30380 18676 30436 19292
rect 30156 18674 30772 18676
rect 30156 18622 30382 18674
rect 30434 18622 30772 18674
rect 30156 18620 30772 18622
rect 29932 18228 29988 18238
rect 29932 18134 29988 18172
rect 29820 17444 29876 17454
rect 29820 17350 29876 17388
rect 29708 16818 29764 16828
rect 29708 16660 29764 16670
rect 29708 16566 29764 16604
rect 30156 16210 30212 18620
rect 30380 18610 30436 18620
rect 30716 18562 30772 18620
rect 30716 18510 30718 18562
rect 30770 18510 30772 18562
rect 30716 18498 30772 18510
rect 30940 17108 30996 17118
rect 30156 16158 30158 16210
rect 30210 16158 30212 16210
rect 30156 16146 30212 16158
rect 30492 16884 30548 16894
rect 29184 15708 29448 15718
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29184 15642 29448 15652
rect 29036 15250 29092 15260
rect 29372 15314 29428 15326
rect 29372 15262 29374 15314
rect 29426 15262 29428 15314
rect 29372 15204 29428 15262
rect 29372 15138 29428 15148
rect 28476 14590 28478 14642
rect 28530 14590 28532 14642
rect 28476 14578 28532 14590
rect 28364 14478 28366 14530
rect 28418 14478 28420 14530
rect 28364 14466 28420 14478
rect 29036 14532 29092 14542
rect 29036 13746 29092 14476
rect 29708 14532 29764 14542
rect 29708 14530 30100 14532
rect 29708 14478 29710 14530
rect 29762 14478 30100 14530
rect 29708 14476 30100 14478
rect 29708 14466 29764 14476
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 29036 13694 29038 13746
rect 29090 13694 29092 13746
rect 29036 13682 29092 13694
rect 29596 13748 29652 13758
rect 29596 13746 29764 13748
rect 29596 13694 29598 13746
rect 29650 13694 29764 13746
rect 29596 13692 29764 13694
rect 29596 13682 29652 13692
rect 28812 13524 28868 13534
rect 28812 13522 28980 13524
rect 28812 13470 28814 13522
rect 28866 13470 28980 13522
rect 28812 13468 28980 13470
rect 28812 13458 28868 13468
rect 28588 13412 28644 13422
rect 28588 12290 28644 13356
rect 28588 12238 28590 12290
rect 28642 12238 28644 12290
rect 28588 12226 28644 12238
rect 28924 10276 28980 13468
rect 29596 12738 29652 12750
rect 29596 12686 29598 12738
rect 29650 12686 29652 12738
rect 29184 12572 29448 12582
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29184 12506 29448 12516
rect 29036 12180 29092 12190
rect 29036 10498 29092 12124
rect 29596 11172 29652 12686
rect 29708 11620 29764 13692
rect 30044 12180 30100 14476
rect 30380 12740 30436 12750
rect 30380 12646 30436 12684
rect 30156 12180 30212 12190
rect 30044 12124 30156 12180
rect 30156 12114 30212 12124
rect 30492 12066 30548 16828
rect 30604 16770 30660 16782
rect 30604 16718 30606 16770
rect 30658 16718 30660 16770
rect 30604 16100 30660 16718
rect 30940 16770 30996 17052
rect 30940 16718 30942 16770
rect 30994 16718 30996 16770
rect 30940 16706 30996 16718
rect 30604 15204 30660 16044
rect 30828 16324 30884 16334
rect 30828 16098 30884 16268
rect 31500 16324 31556 16334
rect 30828 16046 30830 16098
rect 30882 16046 30884 16098
rect 30828 16034 30884 16046
rect 31276 16100 31332 16110
rect 31276 16006 31332 16044
rect 31500 15314 31556 16268
rect 31500 15262 31502 15314
rect 31554 15262 31556 15314
rect 31500 15250 31556 15262
rect 30604 15138 30660 15148
rect 31500 14084 31556 14094
rect 31388 13524 31444 13534
rect 30716 13188 30772 13198
rect 30492 12014 30494 12066
rect 30546 12014 30548 12066
rect 30492 12002 30548 12014
rect 30604 13132 30716 13188
rect 30268 11732 30324 11742
rect 30324 11676 30436 11732
rect 30268 11666 30324 11676
rect 29708 11554 29764 11564
rect 29596 11106 29652 11116
rect 30268 11170 30324 11182
rect 30268 11118 30270 11170
rect 30322 11118 30324 11170
rect 29184 11004 29448 11014
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29184 10938 29448 10948
rect 29036 10446 29038 10498
rect 29090 10446 29092 10498
rect 29036 10434 29092 10446
rect 28924 10220 29988 10276
rect 28252 9650 28308 9660
rect 29596 9828 29652 9838
rect 29184 9436 29448 9446
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29184 9370 29448 9380
rect 27580 9044 27636 9054
rect 27580 8370 27636 8988
rect 28924 8932 28980 8942
rect 28924 8838 28980 8876
rect 27916 8596 27972 8606
rect 27580 8318 27582 8370
rect 27634 8318 27636 8370
rect 27580 8306 27636 8318
rect 27692 8484 27748 8494
rect 27692 7586 27748 8428
rect 27692 7534 27694 7586
rect 27746 7534 27748 7586
rect 27692 7522 27748 7534
rect 27356 7476 27412 7486
rect 27020 6860 27188 6916
rect 27244 6916 27300 6926
rect 27020 6804 27076 6860
rect 26796 6748 27076 6804
rect 26684 6692 26740 6702
rect 26348 5964 26516 6020
rect 26572 6020 26628 6030
rect 24522 5516 24786 5526
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24522 5450 24786 5460
rect 26348 4900 26404 5964
rect 26460 5794 26516 5806
rect 26460 5742 26462 5794
rect 26514 5742 26516 5794
rect 26460 5684 26516 5742
rect 26460 5618 26516 5628
rect 26348 4834 26404 4844
rect 23100 4450 23156 4462
rect 23100 4398 23102 4450
rect 23154 4398 23156 4450
rect 22428 3502 22430 3554
rect 22482 3502 22484 3554
rect 22428 3490 22484 3502
rect 22876 3666 22932 3678
rect 22876 3614 22878 3666
rect 22930 3614 22932 3666
rect 22092 3390 22094 3442
rect 22146 3390 22148 3442
rect 22092 3378 22148 3390
rect 22876 2324 22932 3614
rect 22204 2268 22932 2324
rect 22204 800 22260 2268
rect 23100 2212 23156 4398
rect 26124 4452 26180 4462
rect 26124 4358 26180 4396
rect 26460 4340 26516 4350
rect 26572 4340 26628 5964
rect 26684 6018 26740 6636
rect 26684 5966 26686 6018
rect 26738 5966 26740 6018
rect 26684 5954 26740 5966
rect 26796 5122 26852 6748
rect 27244 6690 27300 6860
rect 27244 6638 27246 6690
rect 27298 6638 27300 6690
rect 27244 6626 27300 6638
rect 27356 6244 27412 7420
rect 27692 6692 27748 6702
rect 27692 6598 27748 6636
rect 27916 6578 27972 8540
rect 29184 7868 29448 7878
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29184 7802 29448 7812
rect 29596 7700 29652 9772
rect 29932 9154 29988 10220
rect 29932 9102 29934 9154
rect 29986 9102 29988 9154
rect 29932 9090 29988 9102
rect 29820 8260 29876 8270
rect 29820 8166 29876 8204
rect 30044 8036 30100 8046
rect 30044 7942 30100 7980
rect 29484 7644 29652 7700
rect 28700 7364 28756 7374
rect 28700 7270 28756 7308
rect 29260 7362 29316 7374
rect 29260 7310 29262 7362
rect 29314 7310 29316 7362
rect 29148 7250 29204 7262
rect 29148 7198 29150 7250
rect 29202 7198 29204 7250
rect 28588 7028 28644 7038
rect 27916 6526 27918 6578
rect 27970 6526 27972 6578
rect 27916 6514 27972 6526
rect 28252 6578 28308 6590
rect 28252 6526 28254 6578
rect 28306 6526 28308 6578
rect 26908 6188 27412 6244
rect 26908 5796 26964 6188
rect 27692 6132 27748 6142
rect 27692 6038 27748 6076
rect 27020 6020 27076 6030
rect 28028 6020 28084 6030
rect 27020 6018 27300 6020
rect 27020 5966 27022 6018
rect 27074 5966 27300 6018
rect 27020 5964 27300 5966
rect 27020 5954 27076 5964
rect 26908 5740 27076 5796
rect 26796 5070 26798 5122
rect 26850 5070 26852 5122
rect 26796 5058 26852 5070
rect 26908 5348 26964 5358
rect 26684 4564 26740 4574
rect 26684 4470 26740 4508
rect 26460 4338 26628 4340
rect 26460 4286 26462 4338
rect 26514 4286 26628 4338
rect 26460 4284 26628 4286
rect 26460 4274 26516 4284
rect 24522 3948 24786 3958
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24522 3882 24786 3892
rect 26908 3554 26964 5292
rect 27020 5010 27076 5740
rect 27020 4958 27022 5010
rect 27074 4958 27076 5010
rect 27020 4946 27076 4958
rect 27132 5460 27188 5470
rect 27132 4452 27188 5404
rect 27244 4676 27300 5964
rect 28028 5926 28084 5964
rect 27468 5906 27524 5918
rect 27468 5854 27470 5906
rect 27522 5854 27524 5906
rect 27468 5684 27524 5854
rect 27468 5618 27524 5628
rect 27692 5796 27748 5806
rect 27244 4610 27300 4620
rect 27356 5010 27412 5022
rect 27356 4958 27358 5010
rect 27410 4958 27412 5010
rect 27356 4562 27412 4958
rect 27692 5010 27748 5740
rect 28028 5012 28084 5022
rect 27692 4958 27694 5010
rect 27746 4958 27748 5010
rect 27692 4946 27748 4958
rect 27804 5010 28084 5012
rect 27804 4958 28030 5010
rect 28082 4958 28084 5010
rect 27804 4956 28084 4958
rect 27356 4510 27358 4562
rect 27410 4510 27412 4562
rect 27356 4498 27412 4510
rect 27132 4338 27188 4396
rect 27132 4286 27134 4338
rect 27186 4286 27188 4338
rect 27132 4274 27188 4286
rect 27692 4338 27748 4350
rect 27692 4286 27694 4338
rect 27746 4286 27748 4338
rect 26908 3502 26910 3554
rect 26962 3502 26964 3554
rect 26908 3490 26964 3502
rect 27132 4116 27188 4126
rect 26124 3444 26180 3454
rect 26124 3350 26180 3388
rect 27132 3442 27188 4060
rect 27692 3780 27748 4286
rect 27692 3714 27748 3724
rect 27132 3390 27134 3442
rect 27186 3390 27188 3442
rect 27132 3378 27188 3390
rect 27580 3554 27636 3566
rect 27580 3502 27582 3554
rect 27634 3502 27636 3554
rect 27580 3444 27636 3502
rect 24556 3332 24612 3342
rect 22876 2156 23156 2212
rect 24220 3330 24612 3332
rect 24220 3278 24558 3330
rect 24610 3278 24612 3330
rect 24220 3276 24612 3278
rect 22876 800 22932 2156
rect 24220 800 24276 3276
rect 24556 3266 24612 3276
rect 26460 3332 26516 3342
rect 26460 3330 26740 3332
rect 26460 3278 26462 3330
rect 26514 3278 26740 3330
rect 26460 3276 26740 3278
rect 26460 3266 26516 3276
rect 26684 1764 26740 3276
rect 26684 1708 26964 1764
rect 26908 800 26964 1708
rect 27580 800 27636 3388
rect 27804 3442 27860 4956
rect 28028 4946 28084 4956
rect 28252 4564 28308 6526
rect 28588 6578 28644 6972
rect 28588 6526 28590 6578
rect 28642 6526 28644 6578
rect 28588 6514 28644 6526
rect 28812 6804 28868 6814
rect 28364 6020 28420 6030
rect 28364 5926 28420 5964
rect 28812 5906 28868 6748
rect 29148 6578 29204 7198
rect 29260 6692 29316 7310
rect 29260 6626 29316 6636
rect 29148 6526 29150 6578
rect 29202 6526 29204 6578
rect 29148 6468 29204 6526
rect 29484 6578 29540 7644
rect 29820 7362 29876 7374
rect 29820 7310 29822 7362
rect 29874 7310 29876 7362
rect 29820 7250 29876 7310
rect 29820 7198 29822 7250
rect 29874 7198 29876 7250
rect 29820 7186 29876 7198
rect 29484 6526 29486 6578
rect 29538 6526 29540 6578
rect 29484 6514 29540 6526
rect 30156 6578 30212 6590
rect 30156 6526 30158 6578
rect 30210 6526 30212 6578
rect 28812 5854 28814 5906
rect 28866 5854 28868 5906
rect 28812 5842 28868 5854
rect 28924 6412 29204 6468
rect 29820 6466 29876 6478
rect 29820 6414 29822 6466
rect 29874 6414 29876 6466
rect 28364 4900 28420 4910
rect 28700 4900 28756 4910
rect 28364 4898 28644 4900
rect 28364 4846 28366 4898
rect 28418 4846 28644 4898
rect 28364 4844 28644 4846
rect 28364 4834 28420 4844
rect 28252 4498 28308 4508
rect 28364 4676 28420 4686
rect 28028 4450 28084 4462
rect 28028 4398 28030 4450
rect 28082 4398 28084 4450
rect 28028 3556 28084 4398
rect 28364 4450 28420 4620
rect 28364 4398 28366 4450
rect 28418 4398 28420 4450
rect 28364 4386 28420 4398
rect 28028 3490 28084 3500
rect 28588 3554 28644 4844
rect 28700 4562 28756 4844
rect 28700 4510 28702 4562
rect 28754 4510 28756 4562
rect 28700 4498 28756 4510
rect 28924 4228 28980 6412
rect 29184 6300 29448 6310
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29184 6234 29448 6244
rect 29036 6020 29092 6030
rect 29036 6018 29316 6020
rect 29036 5966 29038 6018
rect 29090 5966 29316 6018
rect 29036 5964 29316 5966
rect 29036 5954 29092 5964
rect 29260 5124 29316 5964
rect 29372 6018 29428 6030
rect 29372 5966 29374 6018
rect 29426 5966 29428 6018
rect 29372 5348 29428 5966
rect 29372 5282 29428 5292
rect 29596 6020 29652 6030
rect 29596 5236 29652 5964
rect 29708 5908 29764 5918
rect 29708 5814 29764 5852
rect 29708 5236 29764 5246
rect 29596 5234 29764 5236
rect 29596 5182 29710 5234
rect 29762 5182 29764 5234
rect 29596 5180 29764 5182
rect 29708 5170 29764 5180
rect 29260 5068 29652 5124
rect 29260 4900 29316 4938
rect 29260 4834 29316 4844
rect 29184 4732 29448 4742
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29184 4666 29448 4676
rect 29036 4564 29092 4574
rect 29036 4470 29092 4508
rect 29372 4340 29428 4350
rect 29036 4228 29092 4238
rect 28924 4172 29036 4228
rect 29036 4162 29092 4172
rect 28924 3668 28980 3678
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 28700 3666 28980 3668
rect 28700 3614 28926 3666
rect 28978 3614 28980 3666
rect 28700 3612 28980 3614
rect 27804 3390 27806 3442
rect 27858 3390 27860 3442
rect 27804 3378 27860 3390
rect 28700 3388 28756 3612
rect 28924 3602 28980 3612
rect 29372 3388 29428 4284
rect 29596 4116 29652 5068
rect 29820 4338 29876 6414
rect 30156 5012 30212 6526
rect 30268 6018 30324 11118
rect 30380 10722 30436 11676
rect 30380 10670 30382 10722
rect 30434 10670 30436 10722
rect 30380 10658 30436 10670
rect 30492 7588 30548 7598
rect 30604 7588 30660 13132
rect 30716 13122 30772 13132
rect 30940 12180 30996 12190
rect 30940 9938 30996 12124
rect 31052 11172 31108 11182
rect 31052 11078 31108 11116
rect 30940 9886 30942 9938
rect 30994 9886 30996 9938
rect 30940 9874 30996 9886
rect 31276 10612 31332 10622
rect 31164 9156 31220 9166
rect 31164 9062 31220 9100
rect 30940 9042 30996 9054
rect 30940 8990 30942 9042
rect 30994 8990 30996 9042
rect 30940 8820 30996 8990
rect 30996 8764 31220 8820
rect 30940 8754 30996 8764
rect 31164 8370 31220 8764
rect 31164 8318 31166 8370
rect 31218 8318 31220 8370
rect 31164 8306 31220 8318
rect 31276 8148 31332 10556
rect 31388 8370 31444 13468
rect 31500 10388 31556 14028
rect 31612 13076 31668 20750
rect 31724 18338 31780 21420
rect 32620 21362 32676 21374
rect 32620 21310 32622 21362
rect 32674 21310 32676 21362
rect 32620 20188 32676 21310
rect 33180 20804 33236 22430
rect 33404 21700 33460 24668
rect 33628 23154 33684 25228
rect 33852 25218 33908 25228
rect 33964 24834 34020 25452
rect 33964 24782 33966 24834
rect 34018 24782 34020 24834
rect 33964 24770 34020 24782
rect 34188 24724 34244 24734
rect 33846 24332 34110 24342
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 33846 24266 34110 24276
rect 34188 24052 34244 24668
rect 34188 23986 34244 23996
rect 33628 23102 33630 23154
rect 33682 23102 33684 23154
rect 33628 23090 33684 23102
rect 33964 23826 34020 23838
rect 33964 23774 33966 23826
rect 34018 23774 34020 23826
rect 33964 22932 34020 23774
rect 33964 22866 34020 22876
rect 33846 22764 34110 22774
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 33846 22698 34110 22708
rect 33852 21700 33908 21710
rect 33404 21698 33908 21700
rect 33404 21646 33406 21698
rect 33458 21646 33854 21698
rect 33906 21646 33908 21698
rect 33404 21644 33908 21646
rect 33404 21476 33460 21644
rect 33852 21634 33908 21644
rect 33404 21410 33460 21420
rect 34188 21474 34244 21486
rect 34188 21422 34190 21474
rect 34242 21422 34244 21474
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 33236 20748 33796 20804
rect 33180 20738 33236 20748
rect 31948 20130 32004 20142
rect 31948 20078 31950 20130
rect 32002 20078 32004 20130
rect 31948 19796 32004 20078
rect 31948 19730 32004 19740
rect 32060 20132 32676 20188
rect 33068 20692 33124 20702
rect 33068 20188 33124 20636
rect 33292 20244 33348 20254
rect 33068 20132 33348 20188
rect 31724 18286 31726 18338
rect 31778 18286 31780 18338
rect 31724 18274 31780 18286
rect 31948 16996 32004 17006
rect 31948 16902 32004 16940
rect 32060 16772 32116 20132
rect 33292 20018 33348 20132
rect 33292 19966 33294 20018
rect 33346 19966 33348 20018
rect 33068 19908 33124 19918
rect 32172 19906 33124 19908
rect 32172 19854 33070 19906
rect 33122 19854 33124 19906
rect 32172 19852 33124 19854
rect 32172 19010 32228 19852
rect 33068 19842 33124 19852
rect 32956 19236 33012 19246
rect 32172 18958 32174 19010
rect 32226 18958 32228 19010
rect 32172 18946 32228 18958
rect 32732 19012 32788 19022
rect 32732 18918 32788 18956
rect 32956 18450 33012 19180
rect 32956 18398 32958 18450
rect 33010 18398 33012 18450
rect 32172 17666 32228 17678
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 32172 16996 32228 17614
rect 32172 16930 32228 16940
rect 32732 17668 32788 17678
rect 32844 17668 32900 17678
rect 32956 17668 33012 18398
rect 32732 17666 33012 17668
rect 32732 17614 32734 17666
rect 32786 17614 32846 17666
rect 32898 17614 33012 17666
rect 32732 17612 33012 17614
rect 32732 16884 32788 17612
rect 32844 17602 32900 17612
rect 33068 17444 33124 17454
rect 33068 16994 33124 17388
rect 33068 16942 33070 16994
rect 33122 16942 33124 16994
rect 33068 16930 33124 16942
rect 32732 16818 32788 16828
rect 33292 16882 33348 19966
rect 33740 20018 33796 20748
rect 34188 20578 34244 21422
rect 34188 20526 34190 20578
rect 34242 20526 34244 20578
rect 34188 20514 34244 20526
rect 33740 19966 33742 20018
rect 33794 19966 33796 20018
rect 33740 19954 33796 19966
rect 34300 20018 34356 20030
rect 34300 19966 34302 20018
rect 34354 19966 34356 20018
rect 33846 19628 34110 19638
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 33846 19562 34110 19572
rect 33516 19236 33572 19246
rect 33516 19142 33572 19180
rect 34300 18564 34356 19966
rect 34412 20020 34468 27692
rect 34524 26516 34580 27916
rect 34636 27076 34692 34638
rect 34748 34354 34804 35308
rect 35196 35140 35252 35980
rect 35644 35812 35700 39200
rect 36316 36596 36372 39200
rect 35644 35746 35700 35756
rect 36092 36540 36372 36596
rect 35420 35700 35476 35710
rect 35196 35074 35252 35084
rect 35308 35698 35476 35700
rect 35308 35646 35422 35698
rect 35474 35646 35476 35698
rect 35308 35644 35476 35646
rect 34972 34804 35028 34814
rect 34748 34302 34750 34354
rect 34802 34302 34804 34354
rect 34748 34290 34804 34302
rect 34860 34802 35028 34804
rect 34860 34750 34974 34802
rect 35026 34750 35028 34802
rect 34860 34748 35028 34750
rect 34860 31948 34916 34748
rect 34972 34738 35028 34748
rect 35308 34802 35364 35644
rect 35420 35634 35476 35644
rect 35644 35140 35700 35150
rect 35644 35046 35700 35084
rect 35308 34750 35310 34802
rect 35362 34750 35364 34802
rect 35308 34738 35364 34750
rect 35196 34356 35252 34366
rect 35084 34130 35140 34142
rect 35084 34078 35086 34130
rect 35138 34078 35140 34130
rect 34972 33684 35028 33694
rect 34972 32786 35028 33628
rect 34972 32734 34974 32786
rect 35026 32734 35028 32786
rect 34972 32722 35028 32734
rect 34748 31892 34916 31948
rect 34748 28084 34804 31892
rect 34748 28018 34804 28028
rect 34860 31108 34916 31118
rect 34636 27010 34692 27020
rect 34860 26516 34916 31052
rect 34524 26460 34692 26516
rect 34524 26292 34580 26302
rect 34524 24722 34580 26236
rect 34524 24670 34526 24722
rect 34578 24670 34580 24722
rect 34524 23156 34580 24670
rect 34524 21586 34580 23100
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 34524 21522 34580 21534
rect 34636 21588 34692 26460
rect 34860 26450 34916 26460
rect 34972 30322 35028 30334
rect 34972 30270 34974 30322
rect 35026 30270 35028 30322
rect 34972 25284 35028 30270
rect 35084 30212 35140 34078
rect 35196 32676 35252 34300
rect 35420 34242 35476 34254
rect 35420 34190 35422 34242
rect 35474 34190 35476 34242
rect 35308 33458 35364 33470
rect 35308 33406 35310 33458
rect 35362 33406 35364 33458
rect 35308 32900 35364 33406
rect 35420 33348 35476 34190
rect 36092 34244 36148 36540
rect 36988 36484 37044 39200
rect 37548 39060 37604 39070
rect 36988 36428 37492 36484
rect 36092 34178 36148 34188
rect 36204 36370 36260 36382
rect 36204 36318 36206 36370
rect 36258 36318 36260 36370
rect 35980 34020 36036 34030
rect 35980 34018 36148 34020
rect 35980 33966 35982 34018
rect 36034 33966 36148 34018
rect 35980 33964 36148 33966
rect 35980 33954 36036 33964
rect 35420 33282 35476 33292
rect 35308 32844 35924 32900
rect 35420 32676 35476 32686
rect 35196 32674 35476 32676
rect 35196 32622 35422 32674
rect 35474 32622 35476 32674
rect 35196 32620 35476 32622
rect 35420 32610 35476 32620
rect 35756 32450 35812 32462
rect 35756 32398 35758 32450
rect 35810 32398 35812 32450
rect 35420 32340 35476 32350
rect 35084 30146 35140 30156
rect 35308 31666 35364 31678
rect 35308 31614 35310 31666
rect 35362 31614 35364 31666
rect 35196 29538 35252 29550
rect 35196 29486 35198 29538
rect 35250 29486 35252 29538
rect 35196 28196 35252 29486
rect 35308 28420 35364 31614
rect 35420 31444 35476 32284
rect 35420 31378 35476 31388
rect 35420 31106 35476 31118
rect 35420 31054 35422 31106
rect 35474 31054 35476 31106
rect 35420 28532 35476 31054
rect 35420 28466 35476 28476
rect 35308 28354 35364 28364
rect 35196 28140 35476 28196
rect 34972 25218 35028 25228
rect 35308 27970 35364 27982
rect 35308 27918 35310 27970
rect 35362 27918 35364 27970
rect 35196 24724 35252 24734
rect 35196 24630 35252 24668
rect 35308 23492 35364 27918
rect 35420 24612 35476 28140
rect 35420 24546 35476 24556
rect 34636 21522 34692 21532
rect 34748 23436 35364 23492
rect 34748 21026 34804 23436
rect 35196 21588 35252 21598
rect 35756 21588 35812 32398
rect 35868 26292 35924 32844
rect 35980 26292 36036 26302
rect 35868 26290 36036 26292
rect 35868 26238 35982 26290
rect 36034 26238 36036 26290
rect 35868 26236 36036 26238
rect 35980 26226 36036 26236
rect 35980 25396 36036 25406
rect 35980 25282 36036 25340
rect 35980 25230 35982 25282
rect 36034 25230 36036 25282
rect 35980 25218 36036 25230
rect 36092 24724 36148 33964
rect 36204 31948 36260 36318
rect 36428 36372 36484 36382
rect 36428 35586 36484 36316
rect 36540 36260 36596 36270
rect 36540 36258 36932 36260
rect 36540 36206 36542 36258
rect 36594 36206 36932 36258
rect 36540 36204 36932 36206
rect 36540 36194 36596 36204
rect 36428 35534 36430 35586
rect 36482 35534 36484 35586
rect 36428 35522 36484 35534
rect 36652 35924 36708 35934
rect 36428 34692 36484 34702
rect 36316 34690 36484 34692
rect 36316 34638 36430 34690
rect 36482 34638 36484 34690
rect 36316 34636 36484 34638
rect 36316 33236 36372 34636
rect 36428 34626 36484 34636
rect 36652 33460 36708 35868
rect 36876 35476 36932 36204
rect 36988 36258 37044 36270
rect 36988 36206 36990 36258
rect 37042 36206 37044 36258
rect 36988 35924 37044 36206
rect 36988 35858 37044 35868
rect 37100 35698 37156 35710
rect 37100 35646 37102 35698
rect 37154 35646 37156 35698
rect 36876 35420 37044 35476
rect 36988 34914 37044 35420
rect 37100 35364 37156 35646
rect 37100 35298 37156 35308
rect 36988 34862 36990 34914
rect 37042 34862 37044 34914
rect 36988 34850 37044 34862
rect 36316 33170 36372 33180
rect 36428 33404 36708 33460
rect 36988 34242 37044 34254
rect 36988 34190 36990 34242
rect 37042 34190 37044 34242
rect 36204 31892 36372 31948
rect 36204 31778 36260 31790
rect 36204 31726 36206 31778
rect 36258 31726 36260 31778
rect 36204 31332 36260 31726
rect 36204 31266 36260 31276
rect 36204 30098 36260 30110
rect 36204 30046 36206 30098
rect 36258 30046 36260 30098
rect 36204 24948 36260 30046
rect 36316 29876 36372 31892
rect 36428 31666 36484 33404
rect 36988 33348 37044 34190
rect 37324 33460 37380 33470
rect 36428 31614 36430 31666
rect 36482 31614 36484 31666
rect 36428 31602 36484 31614
rect 36540 33292 37044 33348
rect 37100 33348 37156 33358
rect 36428 31444 36484 31454
rect 36428 31218 36484 31388
rect 36428 31166 36430 31218
rect 36482 31166 36484 31218
rect 36428 31154 36484 31166
rect 36316 29810 36372 29820
rect 36428 26292 36484 26302
rect 36428 26198 36484 26236
rect 36540 25730 36596 33292
rect 37100 33254 37156 33292
rect 36876 32788 36932 32798
rect 36876 31218 36932 32732
rect 36876 31166 36878 31218
rect 36930 31166 36932 31218
rect 36876 31154 36932 31166
rect 36988 32674 37044 32686
rect 36988 32622 36990 32674
rect 37042 32622 37044 32674
rect 36764 29652 36820 29662
rect 36764 29558 36820 29596
rect 36876 27076 36932 27086
rect 36988 27076 37044 32622
rect 37324 31778 37380 33404
rect 37324 31726 37326 31778
rect 37378 31726 37380 31778
rect 37324 31714 37380 31726
rect 37436 33236 37492 36428
rect 37548 33458 37604 39004
rect 37660 38612 37716 39200
rect 37660 38556 37940 38612
rect 37772 38388 37828 38398
rect 37660 37044 37716 37054
rect 37660 35026 37716 36988
rect 37772 36706 37828 38332
rect 37772 36654 37774 36706
rect 37826 36654 37828 36706
rect 37772 36642 37828 36654
rect 37660 34974 37662 35026
rect 37714 34974 37716 35026
rect 37660 34962 37716 34974
rect 37772 35474 37828 35486
rect 37772 35422 37774 35474
rect 37826 35422 37828 35474
rect 37772 35028 37828 35422
rect 37772 34962 37828 34972
rect 37884 34804 37940 38556
rect 37884 34738 37940 34748
rect 38220 37716 38276 37726
rect 37548 33406 37550 33458
rect 37602 33406 37604 33458
rect 37548 33394 37604 33406
rect 37772 33572 37828 33582
rect 37436 33180 37716 33236
rect 37100 31668 37156 31678
rect 37100 30098 37156 31612
rect 37212 31220 37268 31230
rect 37212 31126 37268 31164
rect 37436 30994 37492 33180
rect 37660 32786 37716 33180
rect 37660 32734 37662 32786
rect 37714 32734 37716 32786
rect 37660 32722 37716 32734
rect 37548 31556 37604 31566
rect 37548 31462 37604 31500
rect 37436 30942 37438 30994
rect 37490 30942 37492 30994
rect 37436 30930 37492 30942
rect 37660 30996 37716 31006
rect 37100 30046 37102 30098
rect 37154 30046 37156 30098
rect 37100 30034 37156 30046
rect 37548 30324 37604 30334
rect 37548 30098 37604 30268
rect 37548 30046 37550 30098
rect 37602 30046 37604 30098
rect 37548 30034 37604 30046
rect 37548 29652 37604 29662
rect 37660 29652 37716 30940
rect 37772 30884 37828 33516
rect 38220 33460 38276 37660
rect 38508 36092 38772 36102
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38508 36026 38772 36036
rect 38220 33366 38276 33404
rect 38332 35700 38388 35710
rect 37884 33236 37940 33246
rect 37884 31666 37940 33180
rect 38220 32788 38276 32798
rect 38332 32788 38388 35644
rect 38508 34524 38772 34534
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38508 34458 38772 34468
rect 38508 32956 38772 32966
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38508 32890 38772 32900
rect 38220 32786 38388 32788
rect 38220 32734 38222 32786
rect 38274 32734 38388 32786
rect 38220 32732 38388 32734
rect 38220 31948 38276 32732
rect 37884 31614 37886 31666
rect 37938 31614 37940 31666
rect 37884 31602 37940 31614
rect 38108 31892 38276 31948
rect 37884 31332 37940 31342
rect 37884 31218 37940 31276
rect 37884 31166 37886 31218
rect 37938 31166 37940 31218
rect 37884 31154 37940 31166
rect 38108 31108 38164 31892
rect 38220 31666 38276 31678
rect 38220 31614 38222 31666
rect 38274 31614 38276 31666
rect 38220 31556 38276 31614
rect 38220 31490 38276 31500
rect 38508 31388 38772 31398
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38508 31322 38772 31332
rect 38220 31108 38276 31118
rect 38108 31106 38276 31108
rect 38108 31054 38222 31106
rect 38274 31054 38276 31106
rect 38108 31052 38276 31054
rect 38220 31042 38276 31052
rect 37772 30828 37940 30884
rect 37548 29650 37716 29652
rect 37548 29598 37550 29650
rect 37602 29598 37716 29650
rect 37548 29596 37716 29598
rect 37772 30212 37828 30222
rect 37548 29586 37604 29596
rect 37772 29428 37828 30156
rect 37884 30098 37940 30828
rect 37884 30046 37886 30098
rect 37938 30046 37940 30098
rect 37884 30034 37940 30046
rect 38220 30098 38276 30110
rect 38220 30046 38222 30098
rect 38274 30046 38276 30098
rect 37884 29876 37940 29886
rect 37884 29650 37940 29820
rect 37884 29598 37886 29650
rect 37938 29598 37940 29650
rect 37884 29586 37940 29598
rect 38220 29652 38276 30046
rect 38508 29820 38772 29830
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38508 29754 38772 29764
rect 38220 29586 38276 29596
rect 37772 29372 37940 29428
rect 37212 29314 37268 29326
rect 37212 29262 37214 29314
rect 37266 29262 37268 29314
rect 37212 28980 37268 29262
rect 37212 28914 37268 28924
rect 37660 28644 37716 28654
rect 37660 28550 37716 28588
rect 37884 28530 37940 29372
rect 38220 29426 38276 29438
rect 38220 29374 38222 29426
rect 38274 29374 38276 29426
rect 38220 28980 38276 29374
rect 38220 28914 38276 28924
rect 38108 28644 38164 28654
rect 38108 28550 38164 28588
rect 37884 28478 37886 28530
rect 37938 28478 37940 28530
rect 37884 28466 37940 28478
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 37884 28084 37940 28094
rect 37884 27990 37940 28028
rect 38220 27858 38276 27870
rect 38220 27806 38222 27858
rect 38274 27806 38276 27858
rect 37660 27746 37716 27758
rect 37660 27694 37662 27746
rect 37714 27694 37716 27746
rect 37660 27636 37716 27694
rect 37660 27570 37716 27580
rect 38220 27636 38276 27806
rect 38220 27570 38276 27580
rect 36988 27020 37156 27076
rect 36876 26964 36932 27020
rect 36876 26908 37044 26964
rect 36988 26850 37044 26908
rect 36988 26798 36990 26850
rect 37042 26798 37044 26850
rect 36988 26786 37044 26798
rect 36540 25678 36542 25730
rect 36594 25678 36596 25730
rect 36540 25666 36596 25678
rect 36988 25396 37044 25406
rect 36988 25302 37044 25340
rect 36204 24882 36260 24892
rect 36092 24658 36148 24668
rect 36988 24052 37044 24062
rect 36988 23958 37044 23996
rect 37100 23604 37156 27020
rect 37772 26962 37828 26974
rect 37772 26910 37774 26962
rect 37826 26910 37828 26962
rect 37548 26402 37604 26414
rect 37548 26350 37550 26402
rect 37602 26350 37604 26402
rect 37548 25620 37604 26350
rect 37772 26292 37828 26910
rect 38220 26852 38276 26862
rect 37884 26516 37940 26526
rect 37884 26422 37940 26460
rect 37772 26226 37828 26236
rect 38220 26402 38276 26796
rect 38508 26684 38772 26694
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38508 26618 38772 26628
rect 38220 26350 38222 26402
rect 38274 26350 38276 26402
rect 38220 25620 38276 26350
rect 38332 25620 38388 25630
rect 38220 25618 38388 25620
rect 38220 25566 38334 25618
rect 38386 25566 38388 25618
rect 38220 25564 38388 25566
rect 37548 25554 37604 25564
rect 38332 25554 38388 25564
rect 36876 23548 37156 23604
rect 37212 25506 37268 25518
rect 37212 25454 37214 25506
rect 37266 25454 37268 25506
rect 37212 24052 37268 25454
rect 38508 25116 38772 25126
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38508 25050 38772 25060
rect 38220 24948 38276 24958
rect 38220 24854 38276 24892
rect 37436 24834 37492 24846
rect 37436 24782 37438 24834
rect 37490 24782 37492 24834
rect 36092 23380 36148 23390
rect 36092 23286 36148 23324
rect 36652 23380 36708 23390
rect 36876 23380 36932 23548
rect 36652 23378 36932 23380
rect 36652 23326 36654 23378
rect 36706 23326 36932 23378
rect 36652 23324 36932 23326
rect 36988 23380 37044 23390
rect 36652 23314 36708 23324
rect 36988 22482 37044 23324
rect 36988 22430 36990 22482
rect 37042 22430 37044 22482
rect 36988 22418 37044 22430
rect 37212 22484 37268 23996
rect 37324 24052 37380 24062
rect 37436 24052 37492 24782
rect 37324 24050 37492 24052
rect 37324 23998 37326 24050
rect 37378 23998 37492 24050
rect 37324 23996 37492 23998
rect 38220 24612 38276 24622
rect 37324 23986 37380 23996
rect 37660 22484 37716 22494
rect 37212 22482 37716 22484
rect 37212 22430 37662 22482
rect 37714 22430 37716 22482
rect 37212 22428 37716 22430
rect 37212 22370 37268 22428
rect 37660 22418 37716 22428
rect 37212 22318 37214 22370
rect 37266 22318 37268 22370
rect 37212 22306 37268 22318
rect 37772 22146 37828 22158
rect 37772 22094 37774 22146
rect 37826 22094 37828 22146
rect 37660 21812 37716 21822
rect 37772 21812 37828 22094
rect 37660 21810 37828 21812
rect 37660 21758 37662 21810
rect 37714 21758 37828 21810
rect 37660 21756 37828 21758
rect 38220 21810 38276 24556
rect 38508 23548 38772 23558
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38508 23482 38772 23492
rect 38508 21980 38772 21990
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38508 21914 38772 21924
rect 38220 21758 38222 21810
rect 38274 21758 38276 21810
rect 37660 21746 37716 21756
rect 38220 21746 38276 21758
rect 35196 21586 35812 21588
rect 35196 21534 35198 21586
rect 35250 21534 35812 21586
rect 35196 21532 35812 21534
rect 35196 21522 35252 21532
rect 34748 20974 34750 21026
rect 34802 20974 34804 21026
rect 34748 20962 34804 20974
rect 34972 20690 35028 20702
rect 34972 20638 34974 20690
rect 35026 20638 35028 20690
rect 34972 20244 35028 20638
rect 34860 20132 35028 20188
rect 35084 20578 35140 20590
rect 35084 20526 35086 20578
rect 35138 20526 35140 20578
rect 35084 20188 35140 20526
rect 38332 20578 38388 20590
rect 38332 20526 38334 20578
rect 38386 20526 38388 20578
rect 36764 20242 36820 20254
rect 36764 20190 36766 20242
rect 36818 20190 36820 20242
rect 36764 20188 36820 20190
rect 38332 20188 38388 20526
rect 38508 20412 38772 20422
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38508 20346 38772 20356
rect 35084 20132 35812 20188
rect 36764 20132 37044 20188
rect 34860 20066 34916 20076
rect 34412 19954 34468 19964
rect 34300 18498 34356 18508
rect 35084 19236 35140 19246
rect 33628 18452 33684 18462
rect 33628 18450 34244 18452
rect 33628 18398 33630 18450
rect 33682 18398 34244 18450
rect 33628 18396 34244 18398
rect 33628 18386 33684 18396
rect 33846 18060 34110 18070
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 33846 17994 34110 18004
rect 33516 17666 33572 17678
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33516 17108 33572 17614
rect 33516 17042 33572 17052
rect 33292 16830 33294 16882
rect 33346 16830 33348 16882
rect 33292 16818 33348 16830
rect 31948 16716 32116 16772
rect 31612 13010 31668 13020
rect 31724 15316 31780 15326
rect 31724 12290 31780 15260
rect 31836 13860 31892 13870
rect 31836 13766 31892 13804
rect 31948 12852 32004 16716
rect 33846 16492 34110 16502
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 33846 16426 34110 16436
rect 33740 15988 33796 15998
rect 33740 15538 33796 15932
rect 33740 15486 33742 15538
rect 33794 15486 33796 15538
rect 33740 15474 33796 15486
rect 32956 15204 33012 15214
rect 32956 15110 33012 15148
rect 34188 15148 34244 18396
rect 34972 17108 35028 17118
rect 34636 16996 34692 17006
rect 34300 16884 34356 16894
rect 34300 15988 34356 16828
rect 34636 16660 34692 16940
rect 34748 16884 34804 16894
rect 34748 16790 34804 16828
rect 34636 16604 34804 16660
rect 34636 15988 34692 15998
rect 34300 15986 34692 15988
rect 34300 15934 34638 15986
rect 34690 15934 34692 15986
rect 34300 15932 34692 15934
rect 34636 15316 34692 15932
rect 32284 15092 32340 15102
rect 32284 14998 32340 15036
rect 33292 15092 33348 15102
rect 34188 15092 34356 15148
rect 32844 14532 32900 14542
rect 32900 14476 33012 14532
rect 32844 14438 32900 14476
rect 32172 14308 32228 14318
rect 32172 14214 32228 14252
rect 32732 14308 32788 14318
rect 32732 14306 32900 14308
rect 32732 14254 32734 14306
rect 32786 14254 32900 14306
rect 32732 14252 32900 14254
rect 32732 14242 32788 14252
rect 32732 13972 32788 13982
rect 32620 13522 32676 13534
rect 32620 13470 32622 13522
rect 32674 13470 32676 13522
rect 32620 13188 32676 13470
rect 32620 13122 32676 13132
rect 31948 12786 32004 12796
rect 32620 12962 32676 12974
rect 32620 12910 32622 12962
rect 32674 12910 32676 12962
rect 31724 12238 31726 12290
rect 31778 12238 31780 12290
rect 31724 12226 31780 12238
rect 32396 11620 32452 11630
rect 32284 11564 32396 11620
rect 31500 10332 31780 10388
rect 31612 10164 31668 10174
rect 31500 9268 31556 9278
rect 31500 9154 31556 9212
rect 31500 9102 31502 9154
rect 31554 9102 31556 9154
rect 31500 9090 31556 9102
rect 31388 8318 31390 8370
rect 31442 8318 31444 8370
rect 31388 8306 31444 8318
rect 31276 8092 31444 8148
rect 30492 7586 30660 7588
rect 30492 7534 30494 7586
rect 30546 7534 30660 7586
rect 30492 7532 30660 7534
rect 30492 7522 30548 7532
rect 30604 7028 30660 7038
rect 30492 6804 30548 6814
rect 30492 6578 30548 6748
rect 30492 6526 30494 6578
rect 30546 6526 30548 6578
rect 30492 6514 30548 6526
rect 30268 5966 30270 6018
rect 30322 5966 30324 6018
rect 30268 5954 30324 5966
rect 30380 5348 30436 5358
rect 30380 5234 30436 5292
rect 30380 5182 30382 5234
rect 30434 5182 30436 5234
rect 30380 5170 30436 5182
rect 30156 4946 30212 4956
rect 30492 4900 30548 4910
rect 30492 4562 30548 4844
rect 30604 4676 30660 6972
rect 30604 4610 30660 4620
rect 30716 6690 30772 6702
rect 30716 6638 30718 6690
rect 30770 6638 30772 6690
rect 30716 6580 30772 6638
rect 31276 6580 31332 6590
rect 30716 6578 31332 6580
rect 30716 6526 31278 6578
rect 31330 6526 31332 6578
rect 30716 6524 31332 6526
rect 30492 4510 30494 4562
rect 30546 4510 30548 4562
rect 30492 4498 30548 4510
rect 29820 4286 29822 4338
rect 29874 4286 29876 4338
rect 29820 4274 29876 4286
rect 29596 4060 30100 4116
rect 29708 3780 29764 3790
rect 28252 3332 28756 3388
rect 28924 3332 29428 3388
rect 29596 3668 29652 3678
rect 28252 800 28308 3332
rect 28924 800 28980 3332
rect 29184 3164 29448 3174
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29184 3098 29448 3108
rect 29596 800 29652 3612
rect 29708 3666 29764 3724
rect 29708 3614 29710 3666
rect 29762 3614 29764 3666
rect 29708 3602 29764 3614
rect 30044 3554 30100 4060
rect 30492 3668 30548 3678
rect 30492 3574 30548 3612
rect 30044 3502 30046 3554
rect 30098 3502 30100 3554
rect 30044 3490 30100 3502
rect 30716 3388 30772 6524
rect 31276 6514 31332 6524
rect 31388 5794 31444 8092
rect 31500 7364 31556 7374
rect 31612 7364 31668 10108
rect 31500 7362 31668 7364
rect 31500 7310 31502 7362
rect 31554 7310 31668 7362
rect 31500 7308 31668 7310
rect 31500 7298 31556 7308
rect 31388 5742 31390 5794
rect 31442 5742 31444 5794
rect 31388 5730 31444 5742
rect 31500 7028 31556 7038
rect 30828 5124 30884 5134
rect 31500 5124 31556 6972
rect 30828 5122 31556 5124
rect 30828 5070 30830 5122
rect 30882 5070 31556 5122
rect 30828 5068 31556 5070
rect 30828 5058 30884 5068
rect 31612 5012 31668 5022
rect 31724 5012 31780 10332
rect 31948 9716 32004 9726
rect 31948 9622 32004 9660
rect 31836 9154 31892 9166
rect 31836 9102 31838 9154
rect 31890 9102 31892 9154
rect 31836 7252 31892 9102
rect 31836 7186 31892 7196
rect 32172 9154 32228 9166
rect 32172 9102 32174 9154
rect 32226 9102 32228 9154
rect 32172 7028 32228 9102
rect 32172 6962 32228 6972
rect 31948 5908 32004 5918
rect 31948 5794 32004 5852
rect 31948 5742 31950 5794
rect 32002 5742 32004 5794
rect 31948 5236 32004 5742
rect 32284 5236 32340 11564
rect 32396 11554 32452 11564
rect 32508 10724 32564 10734
rect 32396 9042 32452 9054
rect 32396 8990 32398 9042
rect 32450 8990 32452 9042
rect 32396 8596 32452 8990
rect 32396 8530 32452 8540
rect 32508 8146 32564 10668
rect 32508 8094 32510 8146
rect 32562 8094 32564 8146
rect 32508 8082 32564 8094
rect 32396 6804 32452 6814
rect 32620 6804 32676 12910
rect 32732 9156 32788 13916
rect 32844 10388 32900 14252
rect 32956 13748 33012 14476
rect 33068 14308 33124 14318
rect 33068 13858 33124 14252
rect 33068 13806 33070 13858
rect 33122 13806 33124 13858
rect 33068 13794 33124 13806
rect 32956 12964 33012 13692
rect 33292 13746 33348 15036
rect 33846 14924 34110 14934
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 33846 14858 34110 14868
rect 33404 14530 33460 14542
rect 33404 14478 33406 14530
rect 33458 14478 33460 14530
rect 33404 13972 33460 14478
rect 33404 13906 33460 13916
rect 33740 13860 33796 13870
rect 33740 13766 33796 13804
rect 33292 13694 33294 13746
rect 33346 13694 33348 13746
rect 33292 13636 33348 13694
rect 33964 13746 34020 13758
rect 33964 13694 33966 13746
rect 34018 13694 34020 13746
rect 33292 13570 33348 13580
rect 33628 13636 33684 13646
rect 33068 12964 33124 12974
rect 32956 12962 33460 12964
rect 32956 12910 33070 12962
rect 33122 12910 33460 12962
rect 32956 12908 33460 12910
rect 33068 12898 33124 12908
rect 33292 12740 33348 12750
rect 33292 12290 33348 12684
rect 33292 12238 33294 12290
rect 33346 12238 33348 12290
rect 33292 12226 33348 12238
rect 33404 12068 33460 12908
rect 33628 12404 33684 13580
rect 33964 13636 34020 13694
rect 33964 13570 34020 13580
rect 33846 13356 34110 13366
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 33846 13290 34110 13300
rect 33628 12348 34244 12404
rect 33628 12290 33684 12348
rect 33628 12238 33630 12290
rect 33682 12238 33684 12290
rect 33628 12226 33684 12238
rect 33852 12178 33908 12190
rect 33852 12126 33854 12178
rect 33906 12126 33908 12178
rect 33852 12068 33908 12126
rect 33180 12012 33908 12068
rect 33180 10610 33236 12012
rect 33180 10558 33182 10610
rect 33234 10558 33236 10610
rect 33180 10546 33236 10558
rect 33292 11394 33348 11406
rect 33292 11342 33294 11394
rect 33346 11342 33348 11394
rect 32844 10332 33236 10388
rect 32956 9602 33012 9614
rect 32956 9550 32958 9602
rect 33010 9550 33012 9602
rect 32956 9268 33012 9550
rect 32732 9100 32900 9156
rect 32396 6802 32676 6804
rect 32396 6750 32398 6802
rect 32450 6750 32676 6802
rect 32396 6748 32676 6750
rect 32732 8932 32788 8942
rect 32396 6738 32452 6748
rect 32396 5236 32452 5246
rect 32284 5234 32452 5236
rect 32284 5182 32398 5234
rect 32450 5182 32452 5234
rect 32284 5180 32452 5182
rect 31948 5170 32004 5180
rect 32396 5170 32452 5180
rect 31612 5010 31780 5012
rect 31612 4958 31614 5010
rect 31666 4958 31780 5010
rect 31612 4956 31780 4958
rect 32060 5124 32116 5134
rect 31612 4946 31668 4956
rect 30940 4340 30996 4350
rect 30940 4246 30996 4284
rect 31612 4228 31668 4238
rect 30268 3332 30772 3388
rect 30940 3780 30996 3790
rect 30268 800 30324 3332
rect 30940 800 30996 3724
rect 31612 800 31668 4172
rect 32060 4226 32116 5068
rect 32060 4174 32062 4226
rect 32114 4174 32116 4226
rect 32060 4162 32116 4174
rect 32284 4788 32340 4798
rect 32172 3556 32228 3566
rect 32172 3462 32228 3500
rect 32284 800 32340 4732
rect 32508 4564 32564 4574
rect 32732 4564 32788 8876
rect 32844 7364 32900 9100
rect 32956 8596 33012 9212
rect 32956 8530 33012 8540
rect 33068 7476 33124 7486
rect 32844 7298 32900 7308
rect 32956 7474 33124 7476
rect 32956 7422 33070 7474
rect 33122 7422 33124 7474
rect 32956 7420 33124 7422
rect 32956 6132 33012 7420
rect 33068 7410 33124 7420
rect 32956 6066 33012 6076
rect 33068 7252 33124 7262
rect 33068 6018 33124 7196
rect 33180 6578 33236 10332
rect 33292 10164 33348 11342
rect 33628 11396 33684 12012
rect 33846 11788 34110 11798
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 33846 11722 34110 11732
rect 33740 11396 33796 11406
rect 33628 11394 34132 11396
rect 33628 11342 33742 11394
rect 33794 11342 34132 11394
rect 33628 11340 34132 11342
rect 33740 11330 33796 11340
rect 34076 11060 34132 11340
rect 34188 11284 34244 12348
rect 34300 11732 34356 15092
rect 34636 13748 34692 15260
rect 34636 13682 34692 13692
rect 34636 13524 34692 13534
rect 34524 13076 34580 13086
rect 34524 12982 34580 13020
rect 34524 12178 34580 12190
rect 34524 12126 34526 12178
rect 34578 12126 34580 12178
rect 34300 11676 34468 11732
rect 34188 11218 34244 11228
rect 34300 11506 34356 11518
rect 34300 11454 34302 11506
rect 34354 11454 34356 11506
rect 34300 11172 34356 11454
rect 34300 11106 34356 11116
rect 34076 11004 34244 11060
rect 33628 10612 33684 10622
rect 33628 10518 33684 10556
rect 33846 10220 34110 10230
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 33846 10154 34110 10164
rect 33292 10098 33348 10108
rect 34076 10052 34132 10062
rect 33964 9996 34076 10052
rect 33852 9940 33908 9950
rect 33852 9846 33908 9884
rect 33404 9604 33460 9614
rect 33292 9154 33348 9166
rect 33292 9102 33294 9154
rect 33346 9102 33348 9154
rect 33292 6916 33348 9102
rect 33404 7698 33460 9548
rect 33964 9266 34020 9996
rect 34076 9986 34132 9996
rect 33964 9214 33966 9266
rect 34018 9214 34020 9266
rect 33964 9202 34020 9214
rect 33628 9156 33684 9166
rect 33628 9062 33684 9100
rect 34188 9042 34244 11004
rect 34188 8990 34190 9042
rect 34242 8990 34244 9042
rect 34188 8978 34244 8990
rect 34412 8820 34468 11676
rect 34524 11620 34580 12126
rect 34524 11554 34580 11564
rect 34524 11284 34580 11294
rect 34524 11190 34580 11228
rect 34188 8764 34468 8820
rect 33846 8652 34110 8662
rect 33404 7646 33406 7698
rect 33458 7646 33460 7698
rect 33404 7634 33460 7646
rect 33628 8596 33684 8606
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 33846 8586 34110 8596
rect 33292 6850 33348 6860
rect 33180 6526 33182 6578
rect 33234 6526 33236 6578
rect 33180 6514 33236 6526
rect 33404 6468 33460 6478
rect 33404 6130 33460 6412
rect 33404 6078 33406 6130
rect 33458 6078 33460 6130
rect 33404 6066 33460 6078
rect 33068 5966 33070 6018
rect 33122 5966 33124 6018
rect 33068 5954 33124 5966
rect 32508 4562 32788 4564
rect 32508 4510 32510 4562
rect 32562 4510 32788 4562
rect 32508 4508 32788 4510
rect 33180 5460 33236 5470
rect 32508 4498 32564 4508
rect 33068 4340 33124 4350
rect 32620 4338 33124 4340
rect 32620 4286 33070 4338
rect 33122 4286 33124 4338
rect 32620 4284 33124 4286
rect 32508 3444 32564 3454
rect 32620 3444 32676 4284
rect 33068 4274 33124 4284
rect 32508 3442 32676 3444
rect 32508 3390 32510 3442
rect 32562 3390 32676 3442
rect 32508 3388 32676 3390
rect 33068 3444 33124 3482
rect 32508 3378 32564 3388
rect 33068 3378 33124 3388
rect 33180 1764 33236 5404
rect 33628 5348 33684 8540
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 34076 6916 34132 6926
rect 34076 6580 34132 6860
rect 34188 6802 34244 8764
rect 34636 8708 34692 13468
rect 34748 9940 34804 16604
rect 34748 9874 34804 9884
rect 34748 9716 34804 9726
rect 34748 9622 34804 9660
rect 34972 9492 35028 17052
rect 34972 9426 35028 9436
rect 34748 9044 34804 9054
rect 34748 8950 34804 8988
rect 34188 6750 34190 6802
rect 34242 6750 34244 6802
rect 34188 6738 34244 6750
rect 34300 8652 34692 8708
rect 34076 6524 34244 6580
rect 33852 5906 33908 5918
rect 33852 5854 33854 5906
rect 33906 5854 33908 5906
rect 33852 5796 33908 5854
rect 33852 5730 33908 5740
rect 33846 5516 34110 5526
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 33846 5450 34110 5460
rect 33628 5292 33796 5348
rect 33516 4228 33572 4238
rect 33516 4134 33572 4172
rect 33740 4116 33796 5292
rect 34188 4228 34244 6524
rect 34188 4162 34244 4172
rect 33628 4060 33796 4116
rect 33628 3388 33684 4060
rect 33846 3948 34110 3958
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 33846 3882 34110 3892
rect 34300 3666 34356 8652
rect 34636 8372 34692 8382
rect 35084 8372 35140 19180
rect 35756 19122 35812 20132
rect 36988 19346 37044 20132
rect 37436 20132 37492 20142
rect 37324 19796 37380 19806
rect 36988 19294 36990 19346
rect 37042 19294 37044 19346
rect 36988 19282 37044 19294
rect 37100 19794 37380 19796
rect 37100 19742 37326 19794
rect 37378 19742 37380 19794
rect 37100 19740 37380 19742
rect 35756 19070 35758 19122
rect 35810 19070 35812 19122
rect 35756 19058 35812 19070
rect 36540 19010 36596 19022
rect 36540 18958 36542 19010
rect 36594 18958 36596 19010
rect 36092 18674 36148 18686
rect 36092 18622 36094 18674
rect 36146 18622 36148 18674
rect 36092 18452 36148 18622
rect 36092 18386 36148 18396
rect 35980 18340 36036 18350
rect 35868 18228 35924 18238
rect 35644 18172 35868 18228
rect 35196 13746 35252 13758
rect 35196 13694 35198 13746
rect 35250 13694 35252 13746
rect 35196 13524 35252 13694
rect 35196 13458 35252 13468
rect 35532 12852 35588 12862
rect 35532 12758 35588 12796
rect 35196 11172 35252 11182
rect 35196 11078 35252 11116
rect 35420 11170 35476 11182
rect 35420 11118 35422 11170
rect 35474 11118 35476 11170
rect 35420 10500 35476 11118
rect 35420 10434 35476 10444
rect 35532 9602 35588 9614
rect 35532 9550 35534 9602
rect 35586 9550 35588 9602
rect 35532 8932 35588 9550
rect 35532 8866 35588 8876
rect 34636 8370 35140 8372
rect 34636 8318 34638 8370
rect 34690 8318 35140 8370
rect 34636 8316 35140 8318
rect 34636 8306 34692 8316
rect 35644 8146 35700 18172
rect 35868 18162 35924 18172
rect 35980 17442 36036 18284
rect 36540 17668 36596 18958
rect 36764 18564 36820 18574
rect 36652 18228 36708 18238
rect 36652 18134 36708 18172
rect 36540 17612 36708 17668
rect 36540 17444 36596 17454
rect 35980 17390 35982 17442
rect 36034 17390 36036 17442
rect 35980 17378 36036 17390
rect 36092 17442 36596 17444
rect 36092 17390 36542 17442
rect 36594 17390 36596 17442
rect 36092 17388 36596 17390
rect 35980 15314 36036 15326
rect 35980 15262 35982 15314
rect 36034 15262 36036 15314
rect 35980 15204 36036 15262
rect 35980 15138 36036 15148
rect 35980 14306 36036 14318
rect 35980 14254 35982 14306
rect 36034 14254 36036 14306
rect 35980 13188 36036 14254
rect 35980 13122 36036 13132
rect 35980 12740 36036 12750
rect 35868 12684 35980 12740
rect 35756 11282 35812 11294
rect 35756 11230 35758 11282
rect 35810 11230 35812 11282
rect 35756 11172 35812 11230
rect 35756 11106 35812 11116
rect 35868 10834 35924 12684
rect 35980 12674 36036 12684
rect 36092 11396 36148 17388
rect 36540 17378 36596 17388
rect 35868 10782 35870 10834
rect 35922 10782 35924 10834
rect 35868 10770 35924 10782
rect 35980 11340 36148 11396
rect 36204 16884 36260 16894
rect 35980 10612 36036 11340
rect 35868 10556 36036 10612
rect 36092 11170 36148 11182
rect 36092 11118 36094 11170
rect 36146 11118 36148 11170
rect 35756 9828 35812 9838
rect 35756 9734 35812 9772
rect 35868 8484 35924 10556
rect 35980 10276 36036 10286
rect 35980 8932 36036 10220
rect 36092 9044 36148 11118
rect 36204 9940 36260 16828
rect 36428 15316 36484 15326
rect 36428 15222 36484 15260
rect 36540 14306 36596 14318
rect 36540 14254 36542 14306
rect 36594 14254 36596 14306
rect 36540 14084 36596 14254
rect 36540 14018 36596 14028
rect 36428 11282 36484 11294
rect 36428 11230 36430 11282
rect 36482 11230 36484 11282
rect 36428 10836 36484 11230
rect 36428 10770 36484 10780
rect 36652 10612 36708 17612
rect 36764 15148 36820 18508
rect 36876 18452 36932 18462
rect 36876 18358 36932 18396
rect 36988 15988 37044 15998
rect 36988 15894 37044 15932
rect 36764 15092 36932 15148
rect 36540 10556 36708 10612
rect 36540 10276 36596 10556
rect 36652 10388 36708 10398
rect 36652 10294 36708 10332
rect 36540 10210 36596 10220
rect 36204 9884 36820 9940
rect 36316 9604 36372 9614
rect 36316 9602 36484 9604
rect 36316 9550 36318 9602
rect 36370 9550 36484 9602
rect 36316 9548 36484 9550
rect 36316 9538 36372 9548
rect 36092 8988 36372 9044
rect 35980 8876 36260 8932
rect 35868 8428 36036 8484
rect 35644 8094 35646 8146
rect 35698 8094 35700 8146
rect 35644 8082 35700 8094
rect 35196 7924 35252 7934
rect 35084 7588 35140 7598
rect 34972 7364 35028 7374
rect 34972 7270 35028 7308
rect 34748 6916 34804 6926
rect 34300 3614 34302 3666
rect 34354 3614 34356 3666
rect 34300 3602 34356 3614
rect 34412 5794 34468 5806
rect 34412 5742 34414 5794
rect 34466 5742 34468 5794
rect 33628 3332 34020 3388
rect 32956 1708 33236 1764
rect 32956 800 33012 1708
rect 33964 1092 34020 3332
rect 34412 1876 34468 5742
rect 33964 1026 34020 1036
rect 34076 1820 34468 1876
rect 34524 5236 34580 5246
rect 33628 924 33908 980
rect 33628 800 33684 924
rect 33852 868 33908 924
rect 33852 812 34020 868
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 33964 756 34020 812
rect 34076 756 34132 1820
rect 34524 1764 34580 5180
rect 34636 4338 34692 4350
rect 34636 4286 34638 4338
rect 34690 4286 34692 4338
rect 34636 4116 34692 4286
rect 34636 4050 34692 4060
rect 34748 3444 34804 6860
rect 34972 6580 35028 6590
rect 34972 6486 35028 6524
rect 34748 3378 34804 3388
rect 34972 3668 35028 3678
rect 34300 1708 34580 1764
rect 34300 800 34356 1708
rect 34972 800 35028 3612
rect 35084 2772 35140 7532
rect 35196 5234 35252 7868
rect 35196 5182 35198 5234
rect 35250 5182 35252 5234
rect 35196 5170 35252 5182
rect 35868 6020 35924 6030
rect 35644 5124 35700 5134
rect 35196 4226 35252 4238
rect 35196 4174 35198 4226
rect 35250 4174 35252 4226
rect 35196 3780 35252 4174
rect 35196 3714 35252 3724
rect 35084 2706 35140 2716
rect 35644 800 35700 5068
rect 35868 3388 35924 5964
rect 35980 5012 36036 8428
rect 36092 8372 36148 8382
rect 36092 7586 36148 8316
rect 36092 7534 36094 7586
rect 36146 7534 36148 7586
rect 36092 7522 36148 7534
rect 36092 5012 36148 5022
rect 35980 5010 36148 5012
rect 35980 4958 36094 5010
rect 36146 4958 36148 5010
rect 35980 4956 36148 4958
rect 36092 4946 36148 4956
rect 35980 4676 36036 4686
rect 35980 3554 36036 4620
rect 36204 4676 36260 8876
rect 36316 8260 36372 8988
rect 36316 8194 36372 8204
rect 36316 8034 36372 8046
rect 36316 7982 36318 8034
rect 36370 7982 36372 8034
rect 36316 5684 36372 7982
rect 36428 6916 36484 9548
rect 36652 7588 36708 7598
rect 36652 7494 36708 7532
rect 36764 7364 36820 9884
rect 36428 6850 36484 6860
rect 36652 7308 36820 7364
rect 36316 5618 36372 5628
rect 36652 5572 36708 7308
rect 36764 5796 36820 5806
rect 36876 5796 36932 15092
rect 36988 14418 37044 14430
rect 36988 14366 36990 14418
rect 37042 14366 37044 14418
rect 36988 12402 37044 14366
rect 36988 12350 36990 12402
rect 37042 12350 37044 12402
rect 36988 12338 37044 12350
rect 36988 11396 37044 11406
rect 36988 11302 37044 11340
rect 36988 10610 37044 10622
rect 36988 10558 36990 10610
rect 37042 10558 37044 10610
rect 36988 10164 37044 10558
rect 36988 10098 37044 10108
rect 36988 9604 37044 9614
rect 36988 9510 37044 9548
rect 37100 8372 37156 19740
rect 37324 19730 37380 19740
rect 37324 19348 37380 19358
rect 37436 19348 37492 20076
rect 37884 20132 37940 20142
rect 38220 20132 38948 20188
rect 37884 20130 38164 20132
rect 37884 20078 37886 20130
rect 37938 20078 38164 20130
rect 37884 20076 38164 20078
rect 37884 20066 37940 20076
rect 37660 19348 37716 19358
rect 37212 19346 37716 19348
rect 37212 19294 37326 19346
rect 37378 19294 37662 19346
rect 37714 19294 37716 19346
rect 37212 19292 37716 19294
rect 37212 18562 37268 19292
rect 37324 19282 37380 19292
rect 37212 18510 37214 18562
rect 37266 18510 37268 18562
rect 37212 18498 37268 18510
rect 37548 18562 37604 19292
rect 37660 19282 37716 19292
rect 37548 18510 37550 18562
rect 37602 18510 37604 18562
rect 37548 18498 37604 18510
rect 37772 19010 37828 19022
rect 37772 18958 37774 19010
rect 37826 18958 37828 19010
rect 37772 18004 37828 18958
rect 37884 18340 37940 18350
rect 37884 18246 37940 18284
rect 37212 17948 37828 18004
rect 37212 17106 37268 17948
rect 37212 17054 37214 17106
rect 37266 17054 37268 17106
rect 37212 17042 37268 17054
rect 37548 17778 37604 17790
rect 37548 17726 37550 17778
rect 37602 17726 37604 17778
rect 37548 16884 37604 17726
rect 37548 16818 37604 16828
rect 37772 16660 37828 16670
rect 37772 16658 38052 16660
rect 37772 16606 37774 16658
rect 37826 16606 38052 16658
rect 37772 16604 38052 16606
rect 37772 16594 37828 16604
rect 37212 16098 37268 16110
rect 37212 16046 37214 16098
rect 37266 16046 37268 16098
rect 37212 15988 37268 16046
rect 37660 15988 37716 15998
rect 37212 15986 37716 15988
rect 37212 15934 37662 15986
rect 37714 15934 37716 15986
rect 37212 15932 37716 15934
rect 37212 14530 37268 15932
rect 37660 15922 37716 15932
rect 37212 14478 37214 14530
rect 37266 14478 37268 14530
rect 37212 13636 37268 14478
rect 37772 15874 37828 15886
rect 37772 15822 37774 15874
rect 37826 15822 37828 15874
rect 37772 13970 37828 15822
rect 37772 13918 37774 13970
rect 37826 13918 37828 13970
rect 37772 13906 37828 13918
rect 37212 13076 37268 13580
rect 37884 13188 37940 13198
rect 37660 13076 37716 13086
rect 37212 13074 37716 13076
rect 37212 13022 37662 13074
rect 37714 13022 37716 13074
rect 37212 13020 37716 13022
rect 37212 12962 37268 13020
rect 37212 12910 37214 12962
rect 37266 12910 37268 12962
rect 37212 12898 37268 12910
rect 37212 12740 37268 12750
rect 37212 12646 37268 12684
rect 37324 12628 37380 12638
rect 37324 9266 37380 12572
rect 37436 12404 37492 13020
rect 37660 13010 37716 13020
rect 37772 12740 37828 12778
rect 37772 12674 37828 12684
rect 37436 12348 37828 12404
rect 37772 12290 37828 12348
rect 37884 12402 37940 13132
rect 37884 12350 37886 12402
rect 37938 12350 37940 12402
rect 37884 12338 37940 12350
rect 37772 12238 37774 12290
rect 37826 12238 37828 12290
rect 37772 12226 37828 12238
rect 37548 11954 37604 11966
rect 37548 11902 37550 11954
rect 37602 11902 37604 11954
rect 37548 10724 37604 11902
rect 37548 10658 37604 10668
rect 37324 9214 37326 9266
rect 37378 9214 37380 9266
rect 37324 9202 37380 9214
rect 37548 10498 37604 10510
rect 37548 10446 37550 10498
rect 37602 10446 37604 10498
rect 37100 8306 37156 8316
rect 36988 8036 37044 8046
rect 36988 7942 37044 7980
rect 36988 7476 37044 7486
rect 36988 7382 37044 7420
rect 36988 6468 37044 6478
rect 36988 6374 37044 6412
rect 37548 6132 37604 10446
rect 37772 10052 37828 10062
rect 37772 9958 37828 9996
rect 37772 9268 37828 9278
rect 37772 8370 37828 9212
rect 37884 8818 37940 8830
rect 37884 8766 37886 8818
rect 37938 8766 37940 8818
rect 37884 8484 37940 8766
rect 37884 8418 37940 8428
rect 37772 8318 37774 8370
rect 37826 8318 37828 8370
rect 37772 8306 37828 8318
rect 37772 7476 37828 7486
rect 37548 6066 37604 6076
rect 37660 6692 37716 6702
rect 36764 5794 36932 5796
rect 36764 5742 36766 5794
rect 36818 5742 36932 5794
rect 36764 5740 36932 5742
rect 36764 5730 36820 5740
rect 37436 5684 37492 5694
rect 36652 5516 36820 5572
rect 36204 4610 36260 4620
rect 36764 4226 36820 5516
rect 36988 5348 37044 5358
rect 37044 5292 37156 5348
rect 36988 5282 37044 5292
rect 36988 5124 37044 5134
rect 36876 5122 37044 5124
rect 36876 5070 36990 5122
rect 37042 5070 37044 5122
rect 36876 5068 37044 5070
rect 36876 4564 36932 5068
rect 36988 5058 37044 5068
rect 36876 4498 36932 4508
rect 36764 4174 36766 4226
rect 36818 4174 36820 4226
rect 36764 4162 36820 4174
rect 36428 3668 36484 3678
rect 36428 3574 36484 3612
rect 35980 3502 35982 3554
rect 36034 3502 36036 3554
rect 35980 3490 36036 3502
rect 37100 3388 37156 5292
rect 35868 3332 36372 3388
rect 36316 800 36372 3332
rect 36988 3332 37156 3388
rect 37324 3554 37380 3566
rect 37324 3502 37326 3554
rect 37378 3502 37380 3554
rect 37324 3332 37380 3502
rect 36988 800 37044 3332
rect 37324 3266 37380 3276
rect 33964 700 34132 756
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37436 84 37492 5628
rect 37548 5012 37604 5022
rect 37548 3442 37604 4956
rect 37548 3390 37550 3442
rect 37602 3390 37604 3442
rect 37548 3378 37604 3390
rect 37660 800 37716 6636
rect 37772 6690 37828 7420
rect 37772 6638 37774 6690
rect 37826 6638 37828 6690
rect 37772 6626 37828 6638
rect 37996 6018 38052 16604
rect 38108 16324 38164 20076
rect 38220 20130 38276 20132
rect 38220 20078 38222 20130
rect 38274 20078 38276 20130
rect 38220 20066 38276 20078
rect 38508 18844 38772 18854
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38508 18778 38772 18788
rect 38220 17668 38276 17678
rect 38220 17666 38388 17668
rect 38220 17614 38222 17666
rect 38274 17614 38388 17666
rect 38220 17612 38388 17614
rect 38220 17602 38276 17612
rect 38108 16258 38164 16268
rect 38332 13970 38388 17612
rect 38508 17276 38772 17286
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38508 17210 38772 17220
rect 38892 16212 38948 20132
rect 38892 16146 38948 16156
rect 38508 15708 38772 15718
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38508 15642 38772 15652
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 38332 13918 38334 13970
rect 38386 13918 38388 13970
rect 38332 13906 38388 13918
rect 38508 12572 38772 12582
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38508 12506 38772 12516
rect 38108 11508 38164 11518
rect 38108 11414 38164 11452
rect 38508 11004 38772 11014
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38508 10938 38772 10948
rect 38332 10836 38388 10846
rect 38332 10742 38388 10780
rect 38508 9436 38772 9446
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38508 9370 38772 9380
rect 38108 8148 38164 8158
rect 38108 7586 38164 8092
rect 38508 7868 38772 7878
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38508 7802 38772 7812
rect 38108 7534 38110 7586
rect 38162 7534 38164 7586
rect 38108 7522 38164 7534
rect 38508 6300 38772 6310
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38508 6234 38772 6244
rect 37996 5966 37998 6018
rect 38050 5966 38052 6018
rect 37996 5954 38052 5966
rect 37772 4900 37828 4910
rect 37772 4898 39060 4900
rect 37772 4846 37774 4898
rect 37826 4846 39060 4898
rect 37772 4844 39060 4846
rect 37772 4834 37828 4844
rect 38508 4732 38772 4742
rect 37772 4676 37828 4686
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38508 4666 38772 4676
rect 37772 4450 37828 4620
rect 37772 4398 37774 4450
rect 37826 4398 37828 4450
rect 37772 4386 37828 4398
rect 38108 4340 38164 4350
rect 37884 3442 37940 3454
rect 37884 3390 37886 3442
rect 37938 3390 37940 3442
rect 37884 3332 37940 3390
rect 37884 1428 37940 3276
rect 37884 1362 37940 1372
rect 38108 980 38164 4284
rect 38508 3164 38772 3174
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38508 3098 38772 3108
rect 38108 924 38388 980
rect 38332 800 38388 924
rect 39004 800 39060 4844
rect 39676 3780 39732 3790
rect 39676 800 39732 3724
rect 37436 18 37492 28
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
<< via2 >>
rect 35196 39676 35252 39732
rect 5874 36874 5930 36876
rect 5874 36822 5876 36874
rect 5876 36822 5928 36874
rect 5928 36822 5930 36874
rect 5874 36820 5930 36822
rect 5978 36874 6034 36876
rect 5978 36822 5980 36874
rect 5980 36822 6032 36874
rect 6032 36822 6034 36874
rect 5978 36820 6034 36822
rect 6082 36874 6138 36876
rect 6082 36822 6084 36874
rect 6084 36822 6136 36874
rect 6136 36822 6138 36874
rect 6082 36820 6138 36822
rect 15198 36874 15254 36876
rect 15198 36822 15200 36874
rect 15200 36822 15252 36874
rect 15252 36822 15254 36874
rect 15198 36820 15254 36822
rect 15302 36874 15358 36876
rect 15302 36822 15304 36874
rect 15304 36822 15356 36874
rect 15356 36822 15358 36874
rect 15302 36820 15358 36822
rect 15406 36874 15462 36876
rect 15406 36822 15408 36874
rect 15408 36822 15460 36874
rect 15460 36822 15462 36874
rect 15406 36820 15462 36822
rect 17948 36258 18004 36260
rect 17948 36206 17950 36258
rect 17950 36206 18002 36258
rect 18002 36206 18004 36258
rect 17948 36204 18004 36206
rect 10536 36090 10592 36092
rect 10536 36038 10538 36090
rect 10538 36038 10590 36090
rect 10590 36038 10592 36090
rect 10536 36036 10592 36038
rect 10640 36090 10696 36092
rect 10640 36038 10642 36090
rect 10642 36038 10694 36090
rect 10694 36038 10696 36090
rect 10640 36036 10696 36038
rect 10744 36090 10800 36092
rect 10744 36038 10746 36090
rect 10746 36038 10798 36090
rect 10798 36038 10800 36090
rect 10744 36036 10800 36038
rect 18620 35756 18676 35812
rect 21532 36876 21588 36932
rect 22540 36876 22596 36932
rect 19860 36090 19916 36092
rect 19860 36038 19862 36090
rect 19862 36038 19914 36090
rect 19914 36038 19916 36090
rect 19860 36036 19916 36038
rect 19964 36090 20020 36092
rect 19964 36038 19966 36090
rect 19966 36038 20018 36090
rect 20018 36038 20020 36090
rect 19964 36036 20020 36038
rect 20068 36090 20124 36092
rect 20068 36038 20070 36090
rect 20070 36038 20122 36090
rect 20122 36038 20124 36090
rect 20068 36036 20124 36038
rect 20188 35922 20244 35924
rect 20188 35870 20190 35922
rect 20190 35870 20242 35922
rect 20242 35870 20244 35922
rect 20188 35868 20244 35870
rect 20748 36204 20804 36260
rect 21532 36204 21588 36260
rect 21084 35868 21140 35924
rect 22652 36258 22708 36260
rect 22652 36206 22654 36258
rect 22654 36206 22706 36258
rect 22706 36206 22708 36258
rect 22652 36204 22708 36206
rect 21868 35810 21924 35812
rect 21868 35758 21870 35810
rect 21870 35758 21922 35810
rect 21922 35758 21924 35810
rect 21868 35756 21924 35758
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 24108 35810 24164 35812
rect 24108 35758 24110 35810
rect 24110 35758 24162 35810
rect 24162 35758 24164 35810
rect 24108 35756 24164 35758
rect 24522 36874 24578 36876
rect 24522 36822 24524 36874
rect 24524 36822 24576 36874
rect 24576 36822 24578 36874
rect 24522 36820 24578 36822
rect 24626 36874 24682 36876
rect 24626 36822 24628 36874
rect 24628 36822 24680 36874
rect 24680 36822 24682 36874
rect 24626 36820 24682 36822
rect 24730 36874 24786 36876
rect 24730 36822 24732 36874
rect 24732 36822 24784 36874
rect 24784 36822 24786 36874
rect 24730 36820 24786 36822
rect 24892 36652 24948 36708
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 23436 34860 23492 34916
rect 25340 34914 25396 34916
rect 25340 34862 25342 34914
rect 25342 34862 25394 34914
rect 25394 34862 25396 34914
rect 25340 34860 25396 34862
rect 24780 34802 24836 34804
rect 24780 34750 24782 34802
rect 24782 34750 24834 34802
rect 24834 34750 24836 34802
rect 24780 34748 24836 34750
rect 26124 36652 26180 36708
rect 27132 36370 27188 36372
rect 27132 36318 27134 36370
rect 27134 36318 27186 36370
rect 27186 36318 27188 36370
rect 27132 36316 27188 36318
rect 27580 36652 27636 36708
rect 26124 35756 26180 35812
rect 26684 34802 26740 34804
rect 26684 34750 26686 34802
rect 26686 34750 26738 34802
rect 26738 34750 26740 34802
rect 26684 34748 26740 34750
rect 28812 36652 28868 36708
rect 28924 36316 28980 36372
rect 29184 36090 29240 36092
rect 29184 36038 29186 36090
rect 29186 36038 29238 36090
rect 29238 36038 29240 36090
rect 29184 36036 29240 36038
rect 29288 36090 29344 36092
rect 29288 36038 29290 36090
rect 29290 36038 29342 36090
rect 29342 36038 29344 36090
rect 29288 36036 29344 36038
rect 29392 36090 29448 36092
rect 29392 36038 29394 36090
rect 29394 36038 29446 36090
rect 29446 36038 29448 36090
rect 29392 36036 29448 36038
rect 29708 36482 29764 36484
rect 29708 36430 29710 36482
rect 29710 36430 29762 36482
rect 29762 36430 29764 36482
rect 29708 36428 29764 36430
rect 30940 36652 30996 36708
rect 30268 36428 30324 36484
rect 30716 36482 30772 36484
rect 30716 36430 30718 36482
rect 30718 36430 30770 36482
rect 30770 36430 30772 36482
rect 30716 36428 30772 36430
rect 32956 36876 33012 36932
rect 33628 36876 33684 36932
rect 32284 36540 32340 36596
rect 32620 36652 32676 36708
rect 30716 36204 30772 36260
rect 32172 36258 32228 36260
rect 32172 36206 32174 36258
rect 32174 36206 32226 36258
rect 32226 36206 32228 36258
rect 32172 36204 32228 36206
rect 31948 35922 32004 35924
rect 31948 35870 31950 35922
rect 31950 35870 32002 35922
rect 32002 35870 32004 35922
rect 31948 35868 32004 35870
rect 32396 35756 32452 35812
rect 10536 34522 10592 34524
rect 10536 34470 10538 34522
rect 10538 34470 10590 34522
rect 10590 34470 10592 34522
rect 10536 34468 10592 34470
rect 10640 34522 10696 34524
rect 10640 34470 10642 34522
rect 10642 34470 10694 34522
rect 10694 34470 10696 34522
rect 10640 34468 10696 34470
rect 10744 34522 10800 34524
rect 10744 34470 10746 34522
rect 10746 34470 10798 34522
rect 10798 34470 10800 34522
rect 10744 34468 10800 34470
rect 19860 34522 19916 34524
rect 19860 34470 19862 34522
rect 19862 34470 19914 34522
rect 19914 34470 19916 34522
rect 19860 34468 19916 34470
rect 19964 34522 20020 34524
rect 19964 34470 19966 34522
rect 19966 34470 20018 34522
rect 20018 34470 20020 34522
rect 19964 34468 20020 34470
rect 20068 34522 20124 34524
rect 20068 34470 20070 34522
rect 20070 34470 20122 34522
rect 20122 34470 20124 34522
rect 20068 34468 20124 34470
rect 29184 34522 29240 34524
rect 29184 34470 29186 34522
rect 29186 34470 29238 34522
rect 29238 34470 29240 34522
rect 29184 34468 29240 34470
rect 29288 34522 29344 34524
rect 29288 34470 29290 34522
rect 29290 34470 29342 34522
rect 29342 34470 29344 34522
rect 29288 34468 29344 34470
rect 29392 34522 29448 34524
rect 29392 34470 29394 34522
rect 29394 34470 29446 34522
rect 29446 34470 29448 34522
rect 29392 34468 29448 34470
rect 5874 33738 5930 33740
rect 5874 33686 5876 33738
rect 5876 33686 5928 33738
rect 5928 33686 5930 33738
rect 5874 33684 5930 33686
rect 5978 33738 6034 33740
rect 5978 33686 5980 33738
rect 5980 33686 6032 33738
rect 6032 33686 6034 33738
rect 5978 33684 6034 33686
rect 6082 33738 6138 33740
rect 6082 33686 6084 33738
rect 6084 33686 6136 33738
rect 6136 33686 6138 33738
rect 6082 33684 6138 33686
rect 15198 33738 15254 33740
rect 15198 33686 15200 33738
rect 15200 33686 15252 33738
rect 15252 33686 15254 33738
rect 15198 33684 15254 33686
rect 15302 33738 15358 33740
rect 15302 33686 15304 33738
rect 15304 33686 15356 33738
rect 15356 33686 15358 33738
rect 15302 33684 15358 33686
rect 15406 33738 15462 33740
rect 15406 33686 15408 33738
rect 15408 33686 15460 33738
rect 15460 33686 15462 33738
rect 15406 33684 15462 33686
rect 24522 33738 24578 33740
rect 24522 33686 24524 33738
rect 24524 33686 24576 33738
rect 24576 33686 24578 33738
rect 24522 33684 24578 33686
rect 24626 33738 24682 33740
rect 24626 33686 24628 33738
rect 24628 33686 24680 33738
rect 24680 33686 24682 33738
rect 24626 33684 24682 33686
rect 24730 33738 24786 33740
rect 24730 33686 24732 33738
rect 24732 33686 24784 33738
rect 24784 33686 24786 33738
rect 24730 33684 24786 33686
rect 10536 32954 10592 32956
rect 10536 32902 10538 32954
rect 10538 32902 10590 32954
rect 10590 32902 10592 32954
rect 10536 32900 10592 32902
rect 10640 32954 10696 32956
rect 10640 32902 10642 32954
rect 10642 32902 10694 32954
rect 10694 32902 10696 32954
rect 10640 32900 10696 32902
rect 10744 32954 10800 32956
rect 10744 32902 10746 32954
rect 10746 32902 10798 32954
rect 10798 32902 10800 32954
rect 10744 32900 10800 32902
rect 19860 32954 19916 32956
rect 19860 32902 19862 32954
rect 19862 32902 19914 32954
rect 19914 32902 19916 32954
rect 19860 32900 19916 32902
rect 19964 32954 20020 32956
rect 19964 32902 19966 32954
rect 19966 32902 20018 32954
rect 20018 32902 20020 32954
rect 19964 32900 20020 32902
rect 20068 32954 20124 32956
rect 20068 32902 20070 32954
rect 20070 32902 20122 32954
rect 20122 32902 20124 32954
rect 20068 32900 20124 32902
rect 29184 32954 29240 32956
rect 29184 32902 29186 32954
rect 29186 32902 29238 32954
rect 29238 32902 29240 32954
rect 29184 32900 29240 32902
rect 29288 32954 29344 32956
rect 29288 32902 29290 32954
rect 29290 32902 29342 32954
rect 29342 32902 29344 32954
rect 29288 32900 29344 32902
rect 29392 32954 29448 32956
rect 29392 32902 29394 32954
rect 29394 32902 29446 32954
rect 29446 32902 29448 32954
rect 29392 32900 29448 32902
rect 5874 32170 5930 32172
rect 5874 32118 5876 32170
rect 5876 32118 5928 32170
rect 5928 32118 5930 32170
rect 5874 32116 5930 32118
rect 5978 32170 6034 32172
rect 5978 32118 5980 32170
rect 5980 32118 6032 32170
rect 6032 32118 6034 32170
rect 5978 32116 6034 32118
rect 6082 32170 6138 32172
rect 6082 32118 6084 32170
rect 6084 32118 6136 32170
rect 6136 32118 6138 32170
rect 6082 32116 6138 32118
rect 15198 32170 15254 32172
rect 15198 32118 15200 32170
rect 15200 32118 15252 32170
rect 15252 32118 15254 32170
rect 15198 32116 15254 32118
rect 15302 32170 15358 32172
rect 15302 32118 15304 32170
rect 15304 32118 15356 32170
rect 15356 32118 15358 32170
rect 15302 32116 15358 32118
rect 15406 32170 15462 32172
rect 15406 32118 15408 32170
rect 15408 32118 15460 32170
rect 15460 32118 15462 32170
rect 15406 32116 15462 32118
rect 24522 32170 24578 32172
rect 24522 32118 24524 32170
rect 24524 32118 24576 32170
rect 24576 32118 24578 32170
rect 24522 32116 24578 32118
rect 24626 32170 24682 32172
rect 24626 32118 24628 32170
rect 24628 32118 24680 32170
rect 24680 32118 24682 32170
rect 24626 32116 24682 32118
rect 24730 32170 24786 32172
rect 24730 32118 24732 32170
rect 24732 32118 24784 32170
rect 24784 32118 24786 32170
rect 24730 32116 24786 32118
rect 10536 31386 10592 31388
rect 10536 31334 10538 31386
rect 10538 31334 10590 31386
rect 10590 31334 10592 31386
rect 10536 31332 10592 31334
rect 10640 31386 10696 31388
rect 10640 31334 10642 31386
rect 10642 31334 10694 31386
rect 10694 31334 10696 31386
rect 10640 31332 10696 31334
rect 10744 31386 10800 31388
rect 10744 31334 10746 31386
rect 10746 31334 10798 31386
rect 10798 31334 10800 31386
rect 10744 31332 10800 31334
rect 19860 31386 19916 31388
rect 19860 31334 19862 31386
rect 19862 31334 19914 31386
rect 19914 31334 19916 31386
rect 19860 31332 19916 31334
rect 19964 31386 20020 31388
rect 19964 31334 19966 31386
rect 19966 31334 20018 31386
rect 20018 31334 20020 31386
rect 19964 31332 20020 31334
rect 20068 31386 20124 31388
rect 20068 31334 20070 31386
rect 20070 31334 20122 31386
rect 20122 31334 20124 31386
rect 20068 31332 20124 31334
rect 29184 31386 29240 31388
rect 29184 31334 29186 31386
rect 29186 31334 29238 31386
rect 29238 31334 29240 31386
rect 29184 31332 29240 31334
rect 29288 31386 29344 31388
rect 29288 31334 29290 31386
rect 29290 31334 29342 31386
rect 29342 31334 29344 31386
rect 29288 31332 29344 31334
rect 29392 31386 29448 31388
rect 29392 31334 29394 31386
rect 29394 31334 29446 31386
rect 29446 31334 29448 31386
rect 29392 31332 29448 31334
rect 33846 36874 33902 36876
rect 33846 36822 33848 36874
rect 33848 36822 33900 36874
rect 33900 36822 33902 36874
rect 33846 36820 33902 36822
rect 33950 36874 34006 36876
rect 33950 36822 33952 36874
rect 33952 36822 34004 36874
rect 34004 36822 34006 36874
rect 33950 36820 34006 36822
rect 34054 36874 34110 36876
rect 34054 36822 34056 36874
rect 34056 36822 34108 36874
rect 34108 36822 34110 36874
rect 34054 36820 34110 36822
rect 34188 36316 34244 36372
rect 33740 35868 33796 35924
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 34412 36594 34468 36596
rect 34412 36542 34414 36594
rect 34414 36542 34466 36594
rect 34466 36542 34468 36594
rect 34412 36540 34468 36542
rect 34524 35698 34580 35700
rect 34524 35646 34526 35698
rect 34526 35646 34578 35698
rect 34578 35646 34580 35698
rect 34524 35644 34580 35646
rect 33516 34802 33572 34804
rect 33516 34750 33518 34802
rect 33518 34750 33570 34802
rect 33570 34750 33572 34802
rect 33516 34748 33572 34750
rect 35308 36370 35364 36372
rect 35308 36318 35310 36370
rect 35310 36318 35362 36370
rect 35362 36318 35364 36370
rect 35308 36316 35364 36318
rect 34748 35810 34804 35812
rect 34748 35758 34750 35810
rect 34750 35758 34802 35810
rect 34802 35758 34804 35810
rect 34748 35756 34804 35758
rect 35084 35810 35140 35812
rect 35084 35758 35086 35810
rect 35086 35758 35138 35810
rect 35138 35758 35140 35810
rect 35084 35756 35140 35758
rect 34748 35308 34804 35364
rect 34076 34242 34132 34244
rect 34076 34190 34078 34242
rect 34078 34190 34130 34242
rect 34130 34190 34132 34242
rect 34076 34188 34132 34190
rect 33846 33738 33902 33740
rect 33846 33686 33848 33738
rect 33848 33686 33900 33738
rect 33900 33686 33902 33738
rect 33846 33684 33902 33686
rect 33950 33738 34006 33740
rect 33950 33686 33952 33738
rect 33952 33686 34004 33738
rect 34004 33686 34006 33738
rect 33950 33684 34006 33686
rect 34054 33738 34110 33740
rect 34054 33686 34056 33738
rect 34056 33686 34108 33738
rect 34108 33686 34110 33738
rect 34054 33684 34110 33686
rect 31612 31164 31668 31220
rect 32620 33180 32676 33236
rect 5874 30602 5930 30604
rect 5874 30550 5876 30602
rect 5876 30550 5928 30602
rect 5928 30550 5930 30602
rect 5874 30548 5930 30550
rect 5978 30602 6034 30604
rect 5978 30550 5980 30602
rect 5980 30550 6032 30602
rect 6032 30550 6034 30602
rect 5978 30548 6034 30550
rect 6082 30602 6138 30604
rect 6082 30550 6084 30602
rect 6084 30550 6136 30602
rect 6136 30550 6138 30602
rect 6082 30548 6138 30550
rect 15198 30602 15254 30604
rect 15198 30550 15200 30602
rect 15200 30550 15252 30602
rect 15252 30550 15254 30602
rect 15198 30548 15254 30550
rect 15302 30602 15358 30604
rect 15302 30550 15304 30602
rect 15304 30550 15356 30602
rect 15356 30550 15358 30602
rect 15302 30548 15358 30550
rect 15406 30602 15462 30604
rect 15406 30550 15408 30602
rect 15408 30550 15460 30602
rect 15460 30550 15462 30602
rect 15406 30548 15462 30550
rect 24522 30602 24578 30604
rect 24522 30550 24524 30602
rect 24524 30550 24576 30602
rect 24576 30550 24578 30602
rect 24522 30548 24578 30550
rect 24626 30602 24682 30604
rect 24626 30550 24628 30602
rect 24628 30550 24680 30602
rect 24680 30550 24682 30602
rect 24626 30548 24682 30550
rect 24730 30602 24786 30604
rect 24730 30550 24732 30602
rect 24732 30550 24784 30602
rect 24784 30550 24786 30602
rect 24730 30548 24786 30550
rect 9436 29932 9492 29988
rect 5874 29034 5930 29036
rect 5874 28982 5876 29034
rect 5876 28982 5928 29034
rect 5928 28982 5930 29034
rect 5874 28980 5930 28982
rect 5978 29034 6034 29036
rect 5978 28982 5980 29034
rect 5980 28982 6032 29034
rect 6032 28982 6034 29034
rect 5978 28980 6034 28982
rect 6082 29034 6138 29036
rect 6082 28982 6084 29034
rect 6084 28982 6136 29034
rect 6136 28982 6138 29034
rect 6082 28980 6138 28982
rect 8652 28700 8708 28756
rect 5516 27916 5572 27972
rect 1484 25340 1540 25396
rect 2156 25394 2212 25396
rect 2156 25342 2158 25394
rect 2158 25342 2210 25394
rect 2210 25342 2212 25394
rect 2156 25340 2212 25342
rect 1596 24780 1652 24836
rect 2268 24834 2324 24836
rect 2268 24782 2270 24834
rect 2270 24782 2322 24834
rect 2322 24782 2324 24834
rect 2268 24780 2324 24782
rect 4284 26236 4340 26292
rect 3500 25618 3556 25620
rect 3500 25566 3502 25618
rect 3502 25566 3554 25618
rect 3554 25566 3556 25618
rect 3500 25564 3556 25566
rect 4060 24668 4116 24724
rect 1932 23826 1988 23828
rect 1932 23774 1934 23826
rect 1934 23774 1986 23826
rect 1986 23774 1988 23826
rect 1932 23772 1988 23774
rect 3500 23436 3556 23492
rect 3724 23660 3780 23716
rect 4060 22482 4116 22484
rect 4060 22430 4062 22482
rect 4062 22430 4114 22482
rect 4114 22430 4116 22482
rect 4060 22428 4116 22430
rect 3052 21644 3108 21700
rect 4172 21532 4228 21588
rect 3948 21420 4004 21476
rect 3052 20860 3108 20916
rect 3612 20018 3668 20020
rect 3612 19966 3614 20018
rect 3614 19966 3666 20018
rect 3666 19966 3668 20018
rect 3612 19964 3668 19966
rect 3052 19740 3108 19796
rect 2380 18956 2436 19012
rect 2156 16882 2212 16884
rect 2156 16830 2158 16882
rect 2158 16830 2210 16882
rect 2210 16830 2212 16882
rect 2156 16828 2212 16830
rect 1708 14812 1764 14868
rect 1596 11676 1652 11732
rect 1932 13468 1988 13524
rect 2044 13244 2100 13300
rect 4060 21308 4116 21364
rect 5292 26290 5348 26292
rect 5292 26238 5294 26290
rect 5294 26238 5346 26290
rect 5346 26238 5348 26290
rect 5292 26236 5348 26238
rect 7980 27970 8036 27972
rect 7980 27918 7982 27970
rect 7982 27918 8034 27970
rect 8034 27918 8036 27970
rect 7980 27916 8036 27918
rect 5874 27466 5930 27468
rect 5874 27414 5876 27466
rect 5876 27414 5928 27466
rect 5928 27414 5930 27466
rect 5874 27412 5930 27414
rect 5978 27466 6034 27468
rect 5978 27414 5980 27466
rect 5980 27414 6032 27466
rect 6032 27414 6034 27466
rect 5978 27412 6034 27414
rect 6082 27466 6138 27468
rect 6082 27414 6084 27466
rect 6084 27414 6136 27466
rect 6136 27414 6138 27466
rect 6082 27412 6138 27414
rect 6076 26908 6132 26964
rect 5628 26290 5684 26292
rect 5628 26238 5630 26290
rect 5630 26238 5682 26290
rect 5682 26238 5684 26290
rect 5628 26236 5684 26238
rect 4620 25564 4676 25620
rect 5180 25228 5236 25284
rect 8316 27692 8372 27748
rect 6972 26908 7028 26964
rect 5874 25898 5930 25900
rect 5874 25846 5876 25898
rect 5876 25846 5928 25898
rect 5928 25846 5930 25898
rect 5874 25844 5930 25846
rect 5978 25898 6034 25900
rect 5978 25846 5980 25898
rect 5980 25846 6032 25898
rect 6032 25846 6034 25898
rect 5978 25844 6034 25846
rect 6082 25898 6138 25900
rect 6082 25846 6084 25898
rect 6084 25846 6136 25898
rect 6136 25846 6138 25898
rect 6082 25844 6138 25846
rect 6300 25394 6356 25396
rect 6300 25342 6302 25394
rect 6302 25342 6354 25394
rect 6354 25342 6356 25394
rect 6300 25340 6356 25342
rect 5628 25228 5684 25284
rect 4732 23324 4788 23380
rect 5292 24722 5348 24724
rect 5292 24670 5294 24722
rect 5294 24670 5346 24722
rect 5346 24670 5348 24722
rect 5292 24668 5348 24670
rect 5874 24330 5930 24332
rect 5874 24278 5876 24330
rect 5876 24278 5928 24330
rect 5928 24278 5930 24330
rect 5874 24276 5930 24278
rect 5978 24330 6034 24332
rect 5978 24278 5980 24330
rect 5980 24278 6032 24330
rect 6032 24278 6034 24330
rect 5978 24276 6034 24278
rect 6082 24330 6138 24332
rect 6082 24278 6084 24330
rect 6084 24278 6136 24330
rect 6136 24278 6138 24330
rect 6082 24276 6138 24278
rect 5740 23826 5796 23828
rect 5740 23774 5742 23826
rect 5742 23774 5794 23826
rect 5794 23774 5796 23826
rect 5740 23772 5796 23774
rect 6300 23772 6356 23828
rect 5852 23714 5908 23716
rect 5852 23662 5854 23714
rect 5854 23662 5906 23714
rect 5906 23662 5908 23714
rect 5852 23660 5908 23662
rect 4956 23100 5012 23156
rect 5964 23436 6020 23492
rect 6636 23826 6692 23828
rect 6636 23774 6638 23826
rect 6638 23774 6690 23826
rect 6690 23774 6692 23826
rect 6636 23772 6692 23774
rect 8428 26460 8484 26516
rect 8092 25452 8148 25508
rect 7084 23436 7140 23492
rect 6412 23154 6468 23156
rect 6412 23102 6414 23154
rect 6414 23102 6466 23154
rect 6466 23102 6468 23154
rect 6412 23100 6468 23102
rect 5874 22762 5930 22764
rect 5874 22710 5876 22762
rect 5876 22710 5928 22762
rect 5928 22710 5930 22762
rect 5874 22708 5930 22710
rect 5978 22762 6034 22764
rect 5978 22710 5980 22762
rect 5980 22710 6032 22762
rect 6032 22710 6034 22762
rect 5978 22708 6034 22710
rect 6082 22762 6138 22764
rect 6082 22710 6084 22762
rect 6084 22710 6136 22762
rect 6136 22710 6138 22762
rect 6082 22708 6138 22710
rect 5404 21586 5460 21588
rect 5404 21534 5406 21586
rect 5406 21534 5458 21586
rect 5458 21534 5460 21586
rect 5404 21532 5460 21534
rect 4284 20972 4340 21028
rect 6076 21420 6132 21476
rect 5964 21308 6020 21364
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 5964 20802 6020 20804
rect 5964 20750 5966 20802
rect 5966 20750 6018 20802
rect 6018 20750 6020 20802
rect 5964 20748 6020 20750
rect 3724 18620 3780 18676
rect 3052 18284 3108 18340
rect 3948 18396 4004 18452
rect 4060 18172 4116 18228
rect 3052 17554 3108 17556
rect 3052 17502 3054 17554
rect 3054 17502 3106 17554
rect 3106 17502 3108 17554
rect 3052 17500 3108 17502
rect 2604 16940 2660 16996
rect 3500 16940 3556 16996
rect 3052 16716 3108 16772
rect 2940 16604 2996 16660
rect 2268 14588 2324 14644
rect 2268 11116 2324 11172
rect 2380 11676 2436 11732
rect 3388 11900 3444 11956
rect 2492 10722 2548 10724
rect 2492 10670 2494 10722
rect 2494 10670 2546 10722
rect 2546 10670 2548 10722
rect 2492 10668 2548 10670
rect 6972 20748 7028 20804
rect 10444 29932 10500 29988
rect 10536 29818 10592 29820
rect 10536 29766 10538 29818
rect 10538 29766 10590 29818
rect 10590 29766 10592 29818
rect 10536 29764 10592 29766
rect 10640 29818 10696 29820
rect 10640 29766 10642 29818
rect 10642 29766 10694 29818
rect 10694 29766 10696 29818
rect 10640 29764 10696 29766
rect 10744 29818 10800 29820
rect 10744 29766 10746 29818
rect 10746 29766 10798 29818
rect 10798 29766 10800 29818
rect 10744 29764 10800 29766
rect 9660 28754 9716 28756
rect 9660 28702 9662 28754
rect 9662 28702 9714 28754
rect 9714 28702 9716 28754
rect 9660 28700 9716 28702
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 10668 27746 10724 27748
rect 10668 27694 10670 27746
rect 10670 27694 10722 27746
rect 10722 27694 10724 27746
rect 10668 27692 10724 27694
rect 9996 27356 10052 27412
rect 9100 26796 9156 26852
rect 8988 25228 9044 25284
rect 7644 22540 7700 22596
rect 8428 22428 8484 22484
rect 7756 21532 7812 21588
rect 8092 20748 8148 20804
rect 7532 20188 7588 20244
rect 5964 19964 6020 20020
rect 5068 16828 5124 16884
rect 4060 16044 4116 16100
rect 4732 15932 4788 15988
rect 3612 14642 3668 14644
rect 3612 14590 3614 14642
rect 3614 14590 3666 14642
rect 3666 14590 3668 14642
rect 3612 14588 3668 14590
rect 8540 21810 8596 21812
rect 8540 21758 8542 21810
rect 8542 21758 8594 21810
rect 8594 21758 8596 21810
rect 8540 21756 8596 21758
rect 7756 19794 7812 19796
rect 7756 19742 7758 19794
rect 7758 19742 7810 19794
rect 7810 19742 7812 19794
rect 7756 19740 7812 19742
rect 5874 19626 5930 19628
rect 5874 19574 5876 19626
rect 5876 19574 5928 19626
rect 5928 19574 5930 19626
rect 5874 19572 5930 19574
rect 5978 19626 6034 19628
rect 5978 19574 5980 19626
rect 5980 19574 6032 19626
rect 6032 19574 6034 19626
rect 5978 19572 6034 19574
rect 6082 19626 6138 19628
rect 6082 19574 6084 19626
rect 6084 19574 6136 19626
rect 6136 19574 6138 19626
rect 6082 19572 6138 19574
rect 5852 19010 5908 19012
rect 5852 18958 5854 19010
rect 5854 18958 5906 19010
rect 5906 18958 5908 19010
rect 5852 18956 5908 18958
rect 5852 18450 5908 18452
rect 5852 18398 5854 18450
rect 5854 18398 5906 18450
rect 5906 18398 5908 18450
rect 5852 18396 5908 18398
rect 5874 18058 5930 18060
rect 5874 18006 5876 18058
rect 5876 18006 5928 18058
rect 5928 18006 5930 18058
rect 5874 18004 5930 18006
rect 5978 18058 6034 18060
rect 5978 18006 5980 18058
rect 5980 18006 6032 18058
rect 6032 18006 6034 18058
rect 5978 18004 6034 18006
rect 6082 18058 6138 18060
rect 6082 18006 6084 18058
rect 6084 18006 6136 18058
rect 6136 18006 6138 18058
rect 6082 18004 6138 18006
rect 5516 17554 5572 17556
rect 5516 17502 5518 17554
rect 5518 17502 5570 17554
rect 5570 17502 5572 17554
rect 5516 17500 5572 17502
rect 5964 16882 6020 16884
rect 5964 16830 5966 16882
rect 5966 16830 6018 16882
rect 6018 16830 6020 16882
rect 5964 16828 6020 16830
rect 5628 16658 5684 16660
rect 5628 16606 5630 16658
rect 5630 16606 5682 16658
rect 5682 16606 5684 16658
rect 5628 16604 5684 16606
rect 5068 15874 5124 15876
rect 5068 15822 5070 15874
rect 5070 15822 5122 15874
rect 5122 15822 5124 15874
rect 5068 15820 5124 15822
rect 7756 18396 7812 18452
rect 9548 25452 9604 25508
rect 10536 26682 10592 26684
rect 10536 26630 10538 26682
rect 10538 26630 10590 26682
rect 10590 26630 10592 26682
rect 10536 26628 10592 26630
rect 10640 26682 10696 26684
rect 10640 26630 10642 26682
rect 10642 26630 10694 26682
rect 10694 26630 10696 26682
rect 10640 26628 10696 26630
rect 10744 26682 10800 26684
rect 10744 26630 10746 26682
rect 10746 26630 10798 26682
rect 10798 26630 10800 26682
rect 10744 26628 10800 26630
rect 10892 26460 10948 26516
rect 10108 25340 10164 25396
rect 10536 25114 10592 25116
rect 10536 25062 10538 25114
rect 10538 25062 10590 25114
rect 10590 25062 10592 25114
rect 10536 25060 10592 25062
rect 10640 25114 10696 25116
rect 10640 25062 10642 25114
rect 10642 25062 10694 25114
rect 10694 25062 10696 25114
rect 10640 25060 10696 25062
rect 10744 25114 10800 25116
rect 10744 25062 10746 25114
rect 10746 25062 10798 25114
rect 10798 25062 10800 25114
rect 10744 25060 10800 25062
rect 12460 29484 12516 29540
rect 12236 29036 12292 29092
rect 12124 28700 12180 28756
rect 11788 27858 11844 27860
rect 11788 27806 11790 27858
rect 11790 27806 11842 27858
rect 11842 27806 11844 27858
rect 11788 27804 11844 27806
rect 11452 26908 11508 26964
rect 11676 26962 11732 26964
rect 11676 26910 11678 26962
rect 11678 26910 11730 26962
rect 11730 26910 11732 26962
rect 11676 26908 11732 26910
rect 11116 25116 11172 25172
rect 11900 25116 11956 25172
rect 11004 25004 11060 25060
rect 10332 24722 10388 24724
rect 10332 24670 10334 24722
rect 10334 24670 10386 24722
rect 10386 24670 10388 24722
rect 10332 24668 10388 24670
rect 11004 24722 11060 24724
rect 11004 24670 11006 24722
rect 11006 24670 11058 24722
rect 11058 24670 11060 24722
rect 11004 24668 11060 24670
rect 11452 24722 11508 24724
rect 11452 24670 11454 24722
rect 11454 24670 11506 24722
rect 11506 24670 11508 24722
rect 11452 24668 11508 24670
rect 9212 22370 9268 22372
rect 9212 22318 9214 22370
rect 9214 22318 9266 22370
rect 9266 22318 9268 22370
rect 9212 22316 9268 22318
rect 10536 23546 10592 23548
rect 10536 23494 10538 23546
rect 10538 23494 10590 23546
rect 10590 23494 10592 23546
rect 10536 23492 10592 23494
rect 10640 23546 10696 23548
rect 10640 23494 10642 23546
rect 10642 23494 10694 23546
rect 10694 23494 10696 23546
rect 10640 23492 10696 23494
rect 10744 23546 10800 23548
rect 10744 23494 10746 23546
rect 10746 23494 10798 23546
rect 10798 23494 10800 23546
rect 10744 23492 10800 23494
rect 10332 23042 10388 23044
rect 10332 22990 10334 23042
rect 10334 22990 10386 23042
rect 10386 22990 10388 23042
rect 10332 22988 10388 22990
rect 10332 22316 10388 22372
rect 9884 22092 9940 22148
rect 9660 21810 9716 21812
rect 9660 21758 9662 21810
rect 9662 21758 9714 21810
rect 9714 21758 9716 21810
rect 9660 21756 9716 21758
rect 9100 21698 9156 21700
rect 9100 21646 9102 21698
rect 9102 21646 9154 21698
rect 9154 21646 9156 21698
rect 9100 21644 9156 21646
rect 9548 20748 9604 20804
rect 9996 21420 10052 21476
rect 8652 18172 8708 18228
rect 8764 20188 8820 20244
rect 7980 17612 8036 17668
rect 6972 17388 7028 17444
rect 6860 16716 6916 16772
rect 7532 16716 7588 16772
rect 5874 16490 5930 16492
rect 5874 16438 5876 16490
rect 5876 16438 5928 16490
rect 5928 16438 5930 16490
rect 5874 16436 5930 16438
rect 5978 16490 6034 16492
rect 5978 16438 5980 16490
rect 5980 16438 6032 16490
rect 6032 16438 6034 16490
rect 5978 16436 6034 16438
rect 6082 16490 6138 16492
rect 6082 16438 6084 16490
rect 6084 16438 6136 16490
rect 6136 16438 6138 16490
rect 6082 16436 6138 16438
rect 8092 16156 8148 16212
rect 4956 14700 5012 14756
rect 4508 13244 4564 13300
rect 5628 15986 5684 15988
rect 5628 15934 5630 15986
rect 5630 15934 5682 15986
rect 5682 15934 5684 15986
rect 5628 15932 5684 15934
rect 5292 15820 5348 15876
rect 6412 15874 6468 15876
rect 6412 15822 6414 15874
rect 6414 15822 6466 15874
rect 6466 15822 6468 15874
rect 6412 15820 6468 15822
rect 4732 10722 4788 10724
rect 4732 10670 4734 10722
rect 4734 10670 4786 10722
rect 4786 10670 4788 10722
rect 4732 10668 4788 10670
rect 4732 9996 4788 10052
rect 3052 8876 3108 8932
rect 2268 8316 2324 8372
rect 3612 8370 3668 8372
rect 3612 8318 3614 8370
rect 3614 8318 3666 8370
rect 3666 8318 3668 8370
rect 3612 8316 3668 8318
rect 4956 9884 5012 9940
rect 5292 10444 5348 10500
rect 7084 15260 7140 15316
rect 5874 14922 5930 14924
rect 5874 14870 5876 14922
rect 5876 14870 5928 14922
rect 5928 14870 5930 14922
rect 5874 14868 5930 14870
rect 5978 14922 6034 14924
rect 5978 14870 5980 14922
rect 5980 14870 6032 14922
rect 6032 14870 6034 14922
rect 5978 14868 6034 14870
rect 6082 14922 6138 14924
rect 6082 14870 6084 14922
rect 6084 14870 6136 14922
rect 6136 14870 6138 14922
rect 6082 14868 6138 14870
rect 7756 15820 7812 15876
rect 8316 16098 8372 16100
rect 8316 16046 8318 16098
rect 8318 16046 8370 16098
rect 8370 16046 8372 16098
rect 8316 16044 8372 16046
rect 5740 13468 5796 13524
rect 5874 13354 5930 13356
rect 5874 13302 5876 13354
rect 5876 13302 5928 13354
rect 5928 13302 5930 13354
rect 5874 13300 5930 13302
rect 5978 13354 6034 13356
rect 5978 13302 5980 13354
rect 5980 13302 6032 13354
rect 6032 13302 6034 13354
rect 5978 13300 6034 13302
rect 6082 13354 6138 13356
rect 6082 13302 6084 13354
rect 6084 13302 6136 13354
rect 6136 13302 6138 13354
rect 6082 13300 6138 13302
rect 5964 12796 6020 12852
rect 5628 12178 5684 12180
rect 5628 12126 5630 12178
rect 5630 12126 5682 12178
rect 5682 12126 5684 12178
rect 5628 12124 5684 12126
rect 5516 11228 5572 11284
rect 5964 11900 6020 11956
rect 5874 11786 5930 11788
rect 5874 11734 5876 11786
rect 5876 11734 5928 11786
rect 5928 11734 5930 11786
rect 5874 11732 5930 11734
rect 5978 11786 6034 11788
rect 5978 11734 5980 11786
rect 5980 11734 6032 11786
rect 6032 11734 6034 11786
rect 5978 11732 6034 11734
rect 6082 11786 6138 11788
rect 6082 11734 6084 11786
rect 6084 11734 6136 11786
rect 6136 11734 6138 11786
rect 6082 11732 6138 11734
rect 5404 9884 5460 9940
rect 5180 8092 5236 8148
rect 5292 5964 5348 6020
rect 5874 10218 5930 10220
rect 5874 10166 5876 10218
rect 5876 10166 5928 10218
rect 5928 10166 5930 10218
rect 5874 10164 5930 10166
rect 5978 10218 6034 10220
rect 5978 10166 5980 10218
rect 5980 10166 6032 10218
rect 6032 10166 6034 10218
rect 5978 10164 6034 10166
rect 6082 10218 6138 10220
rect 6082 10166 6084 10218
rect 6084 10166 6136 10218
rect 6136 10166 6138 10218
rect 6082 10164 6138 10166
rect 6412 11116 6468 11172
rect 6524 9996 6580 10052
rect 5628 8876 5684 8932
rect 5874 8650 5930 8652
rect 5874 8598 5876 8650
rect 5876 8598 5928 8650
rect 5928 8598 5930 8650
rect 5874 8596 5930 8598
rect 5978 8650 6034 8652
rect 5978 8598 5980 8650
rect 5980 8598 6032 8650
rect 6032 8598 6034 8650
rect 5978 8596 6034 8598
rect 6082 8650 6138 8652
rect 6082 8598 6084 8650
rect 6084 8598 6136 8650
rect 6136 8598 6138 8650
rect 6082 8596 6138 8598
rect 6076 8146 6132 8148
rect 6076 8094 6078 8146
rect 6078 8094 6130 8146
rect 6130 8094 6132 8146
rect 6076 8092 6132 8094
rect 6860 12850 6916 12852
rect 6860 12798 6862 12850
rect 6862 12798 6914 12850
rect 6914 12798 6916 12850
rect 6860 12796 6916 12798
rect 7308 12124 7364 12180
rect 6860 11788 6916 11844
rect 7868 11788 7924 11844
rect 7532 11282 7588 11284
rect 7532 11230 7534 11282
rect 7534 11230 7586 11282
rect 7586 11230 7588 11282
rect 7532 11228 7588 11230
rect 6748 10444 6804 10500
rect 6636 7644 6692 7700
rect 7084 8930 7140 8932
rect 7084 8878 7086 8930
rect 7086 8878 7138 8930
rect 7138 8878 7140 8930
rect 7084 8876 7140 8878
rect 7308 8370 7364 8372
rect 7308 8318 7310 8370
rect 7310 8318 7362 8370
rect 7362 8318 7364 8370
rect 7308 8316 7364 8318
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 8316 12290 8372 12292
rect 8316 12238 8318 12290
rect 8318 12238 8370 12290
rect 8370 12238 8372 12290
rect 8316 12236 8372 12238
rect 8092 12124 8148 12180
rect 8092 11676 8148 11732
rect 8204 10780 8260 10836
rect 10108 21084 10164 21140
rect 10536 21978 10592 21980
rect 10536 21926 10538 21978
rect 10538 21926 10590 21978
rect 10590 21926 10592 21978
rect 10536 21924 10592 21926
rect 10640 21978 10696 21980
rect 10640 21926 10642 21978
rect 10642 21926 10694 21978
rect 10694 21926 10696 21978
rect 10640 21924 10696 21926
rect 10744 21978 10800 21980
rect 10744 21926 10746 21978
rect 10746 21926 10798 21978
rect 10798 21926 10800 21978
rect 10744 21924 10800 21926
rect 12348 27356 12404 27412
rect 13356 29538 13412 29540
rect 13356 29486 13358 29538
rect 13358 29486 13410 29538
rect 13410 29486 13412 29538
rect 13356 29484 13412 29486
rect 14476 29036 14532 29092
rect 13020 28476 13076 28532
rect 12572 27804 12628 27860
rect 12572 27020 12628 27076
rect 15198 29034 15254 29036
rect 15198 28982 15200 29034
rect 15200 28982 15252 29034
rect 15252 28982 15254 29034
rect 15198 28980 15254 28982
rect 15302 29034 15358 29036
rect 15302 28982 15304 29034
rect 15304 28982 15356 29034
rect 15356 28982 15358 29034
rect 15302 28980 15358 28982
rect 15406 29034 15462 29036
rect 15406 28982 15408 29034
rect 15408 28982 15460 29034
rect 15460 28982 15462 29034
rect 15406 28980 15462 28982
rect 15260 28754 15316 28756
rect 15260 28702 15262 28754
rect 15262 28702 15314 28754
rect 15314 28702 15316 28754
rect 15260 28700 15316 28702
rect 15708 28700 15764 28756
rect 15036 28476 15092 28532
rect 13244 27692 13300 27748
rect 13468 26962 13524 26964
rect 13468 26910 13470 26962
rect 13470 26910 13522 26962
rect 13522 26910 13524 26962
rect 13468 26908 13524 26910
rect 14588 27074 14644 27076
rect 14588 27022 14590 27074
rect 14590 27022 14642 27074
rect 14642 27022 14644 27074
rect 14588 27020 14644 27022
rect 15372 28028 15428 28084
rect 15198 27466 15254 27468
rect 15198 27414 15200 27466
rect 15200 27414 15252 27466
rect 15252 27414 15254 27466
rect 15198 27412 15254 27414
rect 15302 27466 15358 27468
rect 15302 27414 15304 27466
rect 15304 27414 15356 27466
rect 15356 27414 15358 27466
rect 15302 27412 15358 27414
rect 15406 27466 15462 27468
rect 15406 27414 15408 27466
rect 15408 27414 15460 27466
rect 15460 27414 15462 27466
rect 15406 27412 15462 27414
rect 19860 29818 19916 29820
rect 19860 29766 19862 29818
rect 19862 29766 19914 29818
rect 19914 29766 19916 29818
rect 19860 29764 19916 29766
rect 19964 29818 20020 29820
rect 19964 29766 19966 29818
rect 19966 29766 20018 29818
rect 20018 29766 20020 29818
rect 19964 29764 20020 29766
rect 20068 29818 20124 29820
rect 20068 29766 20070 29818
rect 20070 29766 20122 29818
rect 20122 29766 20124 29818
rect 20068 29764 20124 29766
rect 29184 29818 29240 29820
rect 29184 29766 29186 29818
rect 29186 29766 29238 29818
rect 29238 29766 29240 29818
rect 29184 29764 29240 29766
rect 29288 29818 29344 29820
rect 29288 29766 29290 29818
rect 29290 29766 29342 29818
rect 29342 29766 29344 29818
rect 29288 29764 29344 29766
rect 29392 29818 29448 29820
rect 29392 29766 29394 29818
rect 29394 29766 29446 29818
rect 29446 29766 29448 29818
rect 29392 29764 29448 29766
rect 15820 27692 15876 27748
rect 16044 28476 16100 28532
rect 14700 26460 14756 26516
rect 24522 29034 24578 29036
rect 24522 28982 24524 29034
rect 24524 28982 24576 29034
rect 24576 28982 24578 29034
rect 24522 28980 24578 28982
rect 24626 29034 24682 29036
rect 24626 28982 24628 29034
rect 24628 28982 24680 29034
rect 24680 28982 24682 29034
rect 24626 28980 24682 28982
rect 24730 29034 24786 29036
rect 24730 28982 24732 29034
rect 24732 28982 24784 29034
rect 24784 28982 24786 29034
rect 24730 28980 24786 28982
rect 18060 28754 18116 28756
rect 18060 28702 18062 28754
rect 18062 28702 18114 28754
rect 18114 28702 18116 28754
rect 18060 28700 18116 28702
rect 16268 28028 16324 28084
rect 16380 26514 16436 26516
rect 16380 26462 16382 26514
rect 16382 26462 16434 26514
rect 16434 26462 16436 26514
rect 16380 26460 16436 26462
rect 19068 28530 19124 28532
rect 19068 28478 19070 28530
rect 19070 28478 19122 28530
rect 19122 28478 19124 28530
rect 19068 28476 19124 28478
rect 26012 28476 26068 28532
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 18284 27916 18340 27972
rect 19628 27970 19684 27972
rect 19628 27918 19630 27970
rect 19630 27918 19682 27970
rect 19682 27918 19684 27970
rect 19628 27916 19684 27918
rect 21084 27916 21140 27972
rect 16604 26460 16660 26516
rect 13692 26124 13748 26180
rect 14140 26348 14196 26404
rect 15260 26402 15316 26404
rect 15260 26350 15262 26402
rect 15262 26350 15314 26402
rect 15314 26350 15316 26402
rect 15260 26348 15316 26350
rect 16268 26178 16324 26180
rect 16268 26126 16270 26178
rect 16270 26126 16322 26178
rect 16322 26126 16324 26178
rect 16268 26124 16324 26126
rect 15198 25898 15254 25900
rect 15198 25846 15200 25898
rect 15200 25846 15252 25898
rect 15252 25846 15254 25898
rect 15198 25844 15254 25846
rect 15302 25898 15358 25900
rect 15302 25846 15304 25898
rect 15304 25846 15356 25898
rect 15356 25846 15358 25898
rect 15302 25844 15358 25846
rect 15406 25898 15462 25900
rect 15406 25846 15408 25898
rect 15408 25846 15460 25898
rect 15460 25846 15462 25898
rect 15406 25844 15462 25846
rect 16716 25788 16772 25844
rect 13692 25004 13748 25060
rect 12572 24668 12628 24724
rect 12460 23996 12516 24052
rect 11452 23772 11508 23828
rect 12572 22988 12628 23044
rect 13468 24050 13524 24052
rect 13468 23998 13470 24050
rect 13470 23998 13522 24050
rect 13522 23998 13524 24050
rect 13468 23996 13524 23998
rect 12684 23436 12740 23492
rect 12348 22370 12404 22372
rect 12348 22318 12350 22370
rect 12350 22318 12402 22370
rect 12402 22318 12404 22370
rect 12348 22316 12404 22318
rect 12684 21756 12740 21812
rect 11564 21474 11620 21476
rect 11564 21422 11566 21474
rect 11566 21422 11618 21474
rect 11618 21422 11620 21474
rect 11564 21420 11620 21422
rect 12460 21084 12516 21140
rect 11900 20524 11956 20580
rect 10536 20410 10592 20412
rect 10536 20358 10538 20410
rect 10538 20358 10590 20410
rect 10590 20358 10592 20410
rect 10536 20356 10592 20358
rect 10640 20410 10696 20412
rect 10640 20358 10642 20410
rect 10642 20358 10694 20410
rect 10694 20358 10696 20410
rect 10640 20356 10696 20358
rect 10744 20410 10800 20412
rect 10744 20358 10746 20410
rect 10746 20358 10798 20410
rect 10798 20358 10800 20410
rect 10744 20356 10800 20358
rect 11564 20188 11620 20244
rect 11004 19404 11060 19460
rect 11452 19122 11508 19124
rect 11452 19070 11454 19122
rect 11454 19070 11506 19122
rect 11506 19070 11508 19122
rect 11452 19068 11508 19070
rect 11116 18956 11172 19012
rect 10536 18842 10592 18844
rect 10536 18790 10538 18842
rect 10538 18790 10590 18842
rect 10590 18790 10592 18842
rect 10536 18788 10592 18790
rect 10640 18842 10696 18844
rect 10640 18790 10642 18842
rect 10642 18790 10694 18842
rect 10694 18790 10696 18842
rect 10640 18788 10696 18790
rect 10744 18842 10800 18844
rect 10744 18790 10746 18842
rect 10746 18790 10798 18842
rect 10798 18790 10800 18842
rect 10744 18788 10800 18790
rect 10332 18508 10388 18564
rect 8988 18338 9044 18340
rect 8988 18286 8990 18338
rect 8990 18286 9042 18338
rect 9042 18286 9044 18338
rect 8988 18284 9044 18286
rect 10108 18338 10164 18340
rect 10108 18286 10110 18338
rect 10110 18286 10162 18338
rect 10162 18286 10164 18338
rect 10108 18284 10164 18286
rect 11788 18956 11844 19012
rect 11004 18562 11060 18564
rect 11004 18510 11006 18562
rect 11006 18510 11058 18562
rect 11058 18510 11060 18562
rect 11004 18508 11060 18510
rect 12012 20748 12068 20804
rect 12796 20524 12852 20580
rect 8540 15820 8596 15876
rect 9996 16882 10052 16884
rect 9996 16830 9998 16882
rect 9998 16830 10050 16882
rect 10050 16830 10052 16882
rect 9996 16828 10052 16830
rect 10536 17274 10592 17276
rect 10536 17222 10538 17274
rect 10538 17222 10590 17274
rect 10590 17222 10592 17274
rect 10536 17220 10592 17222
rect 10640 17274 10696 17276
rect 10640 17222 10642 17274
rect 10642 17222 10694 17274
rect 10694 17222 10696 17274
rect 10640 17220 10696 17222
rect 10744 17274 10800 17276
rect 10744 17222 10746 17274
rect 10746 17222 10798 17274
rect 10798 17222 10800 17274
rect 10744 17220 10800 17222
rect 10780 16994 10836 16996
rect 10780 16942 10782 16994
rect 10782 16942 10834 16994
rect 10834 16942 10836 16994
rect 10780 16940 10836 16942
rect 10332 16716 10388 16772
rect 9884 16156 9940 16212
rect 11788 17388 11844 17444
rect 12348 19068 12404 19124
rect 12124 17052 12180 17108
rect 11564 16940 11620 16996
rect 11340 16882 11396 16884
rect 11340 16830 11342 16882
rect 11342 16830 11394 16882
rect 11394 16830 11396 16882
rect 11340 16828 11396 16830
rect 10536 15706 10592 15708
rect 10536 15654 10538 15706
rect 10538 15654 10590 15706
rect 10590 15654 10592 15706
rect 10536 15652 10592 15654
rect 10640 15706 10696 15708
rect 10640 15654 10642 15706
rect 10642 15654 10694 15706
rect 10694 15654 10696 15706
rect 10640 15652 10696 15654
rect 10744 15706 10800 15708
rect 10744 15654 10746 15706
rect 10746 15654 10798 15706
rect 10798 15654 10800 15706
rect 10744 15652 10800 15654
rect 9100 15372 9156 15428
rect 8428 10556 8484 10612
rect 11452 15260 11508 15316
rect 10108 15148 10164 15204
rect 7756 7308 7812 7364
rect 8764 10834 8820 10836
rect 8764 10782 8766 10834
rect 8766 10782 8818 10834
rect 8818 10782 8820 10834
rect 8764 10780 8820 10782
rect 8764 10556 8820 10612
rect 8764 8540 8820 8596
rect 8988 10108 9044 10164
rect 8876 8316 8932 8372
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 9548 12460 9604 12516
rect 9772 12684 9828 12740
rect 9660 11228 9716 11284
rect 10556 12738 10612 12740
rect 10556 12686 10558 12738
rect 10558 12686 10610 12738
rect 10610 12686 10612 12738
rect 10556 12684 10612 12686
rect 10536 12570 10592 12572
rect 10332 12460 10388 12516
rect 10536 12518 10538 12570
rect 10538 12518 10590 12570
rect 10590 12518 10592 12570
rect 10536 12516 10592 12518
rect 10640 12570 10696 12572
rect 10640 12518 10642 12570
rect 10642 12518 10694 12570
rect 10694 12518 10696 12570
rect 10640 12516 10696 12518
rect 10744 12570 10800 12572
rect 10744 12518 10746 12570
rect 10746 12518 10798 12570
rect 10798 12518 10800 12570
rect 10744 12516 10800 12518
rect 10108 12236 10164 12292
rect 9884 11788 9940 11844
rect 9212 9996 9268 10052
rect 9660 10108 9716 10164
rect 10108 11116 10164 11172
rect 10668 11676 10724 11732
rect 10536 11002 10592 11004
rect 10536 10950 10538 11002
rect 10538 10950 10590 11002
rect 10590 10950 10592 11002
rect 10536 10948 10592 10950
rect 10640 11002 10696 11004
rect 10640 10950 10642 11002
rect 10642 10950 10694 11002
rect 10694 10950 10696 11002
rect 10640 10948 10696 10950
rect 10744 11002 10800 11004
rect 10744 10950 10746 11002
rect 10746 10950 10798 11002
rect 10798 10950 10800 11002
rect 10744 10948 10800 10950
rect 10536 9434 10592 9436
rect 10536 9382 10538 9434
rect 10538 9382 10590 9434
rect 10590 9382 10592 9434
rect 10536 9380 10592 9382
rect 10640 9434 10696 9436
rect 10640 9382 10642 9434
rect 10642 9382 10694 9434
rect 10694 9382 10696 9434
rect 10640 9380 10696 9382
rect 10744 9434 10800 9436
rect 10744 9382 10746 9434
rect 10746 9382 10798 9434
rect 10798 9382 10800 9434
rect 10744 9380 10800 9382
rect 9100 8316 9156 8372
rect 10332 8540 10388 8596
rect 6860 6018 6916 6020
rect 6860 5966 6862 6018
rect 6862 5966 6914 6018
rect 6914 5966 6916 6018
rect 6860 5964 6916 5966
rect 11004 11170 11060 11172
rect 11004 11118 11006 11170
rect 11006 11118 11058 11170
rect 11058 11118 11060 11170
rect 11004 11116 11060 11118
rect 11116 10108 11172 10164
rect 11564 11676 11620 11732
rect 12124 16716 12180 16772
rect 12124 15260 12180 15316
rect 11788 10498 11844 10500
rect 11788 10446 11790 10498
rect 11790 10446 11842 10498
rect 11842 10446 11844 10498
rect 11788 10444 11844 10446
rect 12236 11676 12292 11732
rect 13244 20860 13300 20916
rect 14028 22988 14084 23044
rect 13692 21756 13748 21812
rect 13916 20914 13972 20916
rect 13916 20862 13918 20914
rect 13918 20862 13970 20914
rect 13970 20862 13972 20914
rect 13916 20860 13972 20862
rect 15198 24330 15254 24332
rect 15198 24278 15200 24330
rect 15200 24278 15252 24330
rect 15252 24278 15254 24330
rect 15198 24276 15254 24278
rect 15302 24330 15358 24332
rect 15302 24278 15304 24330
rect 15304 24278 15356 24330
rect 15356 24278 15358 24330
rect 15302 24276 15358 24278
rect 15406 24330 15462 24332
rect 15406 24278 15408 24330
rect 15408 24278 15460 24330
rect 15460 24278 15462 24330
rect 15406 24276 15462 24278
rect 16044 23436 16100 23492
rect 14700 23154 14756 23156
rect 14700 23102 14702 23154
rect 14702 23102 14754 23154
rect 14754 23102 14756 23154
rect 14700 23100 14756 23102
rect 15372 23100 15428 23156
rect 15198 22762 15254 22764
rect 15198 22710 15200 22762
rect 15200 22710 15252 22762
rect 15252 22710 15254 22762
rect 15198 22708 15254 22710
rect 15302 22762 15358 22764
rect 15302 22710 15304 22762
rect 15304 22710 15356 22762
rect 15356 22710 15358 22762
rect 15302 22708 15358 22710
rect 15406 22762 15462 22764
rect 15406 22710 15408 22762
rect 15408 22710 15460 22762
rect 15460 22710 15462 22762
rect 15406 22708 15462 22710
rect 14588 22092 14644 22148
rect 15484 22092 15540 22148
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 15036 20972 15092 21028
rect 14812 20860 14868 20916
rect 13580 20578 13636 20580
rect 13580 20526 13582 20578
rect 13582 20526 13634 20578
rect 13634 20526 13636 20578
rect 13580 20524 13636 20526
rect 13356 19458 13412 19460
rect 13356 19406 13358 19458
rect 13358 19406 13410 19458
rect 13410 19406 13412 19458
rect 13356 19404 13412 19406
rect 16716 23436 16772 23492
rect 18508 26460 18564 26516
rect 17836 26124 17892 26180
rect 18620 25788 18676 25844
rect 18844 25228 18900 25284
rect 17164 23436 17220 23492
rect 19860 26682 19916 26684
rect 19860 26630 19862 26682
rect 19862 26630 19914 26682
rect 19914 26630 19916 26682
rect 19860 26628 19916 26630
rect 19964 26682 20020 26684
rect 19964 26630 19966 26682
rect 19966 26630 20018 26682
rect 20018 26630 20020 26682
rect 19964 26628 20020 26630
rect 20068 26682 20124 26684
rect 20068 26630 20070 26682
rect 20070 26630 20122 26682
rect 20122 26630 20124 26682
rect 20068 26628 20124 26630
rect 22316 27970 22372 27972
rect 22316 27918 22318 27970
rect 22318 27918 22370 27970
rect 22370 27918 22372 27970
rect 22316 27916 22372 27918
rect 24220 27692 24276 27748
rect 19404 26178 19460 26180
rect 19404 26126 19406 26178
rect 19406 26126 19458 26178
rect 19458 26126 19460 26178
rect 19404 26124 19460 26126
rect 19292 24834 19348 24836
rect 19292 24782 19294 24834
rect 19294 24782 19346 24834
rect 19346 24782 19348 24834
rect 19292 24780 19348 24782
rect 21644 25564 21700 25620
rect 20860 25394 20916 25396
rect 20860 25342 20862 25394
rect 20862 25342 20914 25394
rect 20914 25342 20916 25394
rect 20860 25340 20916 25342
rect 19860 25114 19916 25116
rect 19860 25062 19862 25114
rect 19862 25062 19914 25114
rect 19914 25062 19916 25114
rect 19860 25060 19916 25062
rect 19964 25114 20020 25116
rect 19964 25062 19966 25114
rect 19966 25062 20018 25114
rect 20018 25062 20020 25114
rect 19964 25060 20020 25062
rect 20068 25114 20124 25116
rect 20068 25062 20070 25114
rect 20070 25062 20122 25114
rect 20122 25062 20124 25114
rect 20068 25060 20124 25062
rect 20300 25228 20356 25284
rect 21532 25228 21588 25284
rect 21308 24780 21364 24836
rect 19860 23546 19916 23548
rect 19860 23494 19862 23546
rect 19862 23494 19914 23546
rect 19914 23494 19916 23546
rect 19860 23492 19916 23494
rect 19964 23546 20020 23548
rect 19964 23494 19966 23546
rect 19966 23494 20018 23546
rect 20018 23494 20020 23546
rect 19964 23492 20020 23494
rect 20068 23546 20124 23548
rect 20068 23494 20070 23546
rect 20070 23494 20122 23546
rect 20122 23494 20124 23546
rect 20068 23492 20124 23494
rect 17388 23042 17444 23044
rect 17388 22990 17390 23042
rect 17390 22990 17442 23042
rect 17442 22990 17444 23042
rect 17388 22988 17444 22990
rect 19516 23212 19572 23268
rect 19292 22316 19348 22372
rect 17836 21644 17892 21700
rect 18508 21698 18564 21700
rect 18508 21646 18510 21698
rect 18510 21646 18562 21698
rect 18562 21646 18564 21698
rect 18508 21644 18564 21646
rect 16380 20802 16436 20804
rect 16380 20750 16382 20802
rect 16382 20750 16434 20802
rect 16434 20750 16436 20802
rect 16380 20748 16436 20750
rect 16716 20524 16772 20580
rect 16380 20242 16436 20244
rect 16380 20190 16382 20242
rect 16382 20190 16434 20242
rect 16434 20190 16436 20242
rect 16380 20188 16436 20190
rect 15036 19852 15092 19908
rect 15198 19626 15254 19628
rect 15198 19574 15200 19626
rect 15200 19574 15252 19626
rect 15252 19574 15254 19626
rect 15198 19572 15254 19574
rect 15302 19626 15358 19628
rect 15302 19574 15304 19626
rect 15304 19574 15356 19626
rect 15356 19574 15358 19626
rect 15302 19572 15358 19574
rect 15406 19626 15462 19628
rect 15406 19574 15408 19626
rect 15408 19574 15460 19626
rect 15460 19574 15462 19626
rect 15406 19572 15462 19574
rect 14140 19010 14196 19012
rect 14140 18958 14142 19010
rect 14142 18958 14194 19010
rect 14194 18958 14196 19010
rect 14140 18956 14196 18958
rect 13804 18620 13860 18676
rect 14812 17836 14868 17892
rect 12908 16716 12964 16772
rect 12796 15426 12852 15428
rect 12796 15374 12798 15426
rect 12798 15374 12850 15426
rect 12850 15374 12852 15426
rect 12796 15372 12852 15374
rect 13916 17666 13972 17668
rect 13916 17614 13918 17666
rect 13918 17614 13970 17666
rect 13970 17614 13972 17666
rect 13916 17612 13972 17614
rect 14028 17106 14084 17108
rect 14028 17054 14030 17106
rect 14030 17054 14082 17106
rect 14082 17054 14084 17106
rect 14028 17052 14084 17054
rect 13580 16828 13636 16884
rect 13580 16044 13636 16100
rect 14140 16098 14196 16100
rect 14140 16046 14142 16098
rect 14142 16046 14194 16098
rect 14194 16046 14196 16098
rect 14140 16044 14196 16046
rect 13580 15372 13636 15428
rect 16156 19964 16212 20020
rect 15198 18058 15254 18060
rect 15198 18006 15200 18058
rect 15200 18006 15252 18058
rect 15252 18006 15254 18058
rect 15198 18004 15254 18006
rect 15302 18058 15358 18060
rect 15302 18006 15304 18058
rect 15304 18006 15356 18058
rect 15356 18006 15358 18058
rect 15302 18004 15358 18006
rect 15406 18058 15462 18060
rect 15406 18006 15408 18058
rect 15408 18006 15460 18058
rect 15460 18006 15462 18058
rect 15406 18004 15462 18006
rect 15484 17052 15540 17108
rect 15198 16490 15254 16492
rect 15198 16438 15200 16490
rect 15200 16438 15252 16490
rect 15252 16438 15254 16490
rect 15198 16436 15254 16438
rect 15302 16490 15358 16492
rect 15302 16438 15304 16490
rect 15304 16438 15356 16490
rect 15356 16438 15358 16490
rect 15302 16436 15358 16438
rect 15406 16490 15462 16492
rect 15406 16438 15408 16490
rect 15408 16438 15460 16490
rect 15460 16438 15462 16490
rect 15406 16436 15462 16438
rect 12460 12348 12516 12404
rect 12124 11282 12180 11284
rect 12124 11230 12126 11282
rect 12126 11230 12178 11282
rect 12178 11230 12180 11282
rect 12124 11228 12180 11230
rect 12236 11116 12292 11172
rect 13020 14476 13076 14532
rect 13804 14530 13860 14532
rect 13804 14478 13806 14530
rect 13806 14478 13858 14530
rect 13858 14478 13860 14530
rect 13804 14476 13860 14478
rect 12908 11170 12964 11172
rect 12908 11118 12910 11170
rect 12910 11118 12962 11170
rect 12962 11118 12964 11170
rect 12908 11116 12964 11118
rect 12460 10556 12516 10612
rect 11788 9324 11844 9380
rect 11900 9996 11956 10052
rect 11228 9042 11284 9044
rect 11228 8990 11230 9042
rect 11230 8990 11282 9042
rect 11282 8990 11284 9042
rect 11228 8988 11284 8990
rect 10536 7866 10592 7868
rect 10536 7814 10538 7866
rect 10538 7814 10590 7866
rect 10590 7814 10592 7866
rect 10536 7812 10592 7814
rect 10640 7866 10696 7868
rect 10640 7814 10642 7866
rect 10642 7814 10694 7866
rect 10694 7814 10696 7866
rect 10640 7812 10696 7814
rect 10744 7866 10800 7868
rect 10744 7814 10746 7866
rect 10746 7814 10798 7866
rect 10798 7814 10800 7866
rect 10744 7812 10800 7814
rect 10668 7644 10724 7700
rect 10556 7362 10612 7364
rect 10556 7310 10558 7362
rect 10558 7310 10610 7362
rect 10610 7310 10612 7362
rect 10556 7308 10612 7310
rect 11676 7308 11732 7364
rect 11788 8316 11844 8372
rect 10536 6298 10592 6300
rect 10536 6246 10538 6298
rect 10538 6246 10590 6298
rect 10590 6246 10592 6298
rect 10536 6244 10592 6246
rect 10640 6298 10696 6300
rect 10640 6246 10642 6298
rect 10642 6246 10694 6298
rect 10694 6246 10696 6298
rect 10640 6244 10696 6246
rect 10744 6298 10800 6300
rect 10744 6246 10746 6298
rect 10746 6246 10798 6298
rect 10798 6246 10800 6298
rect 10744 6244 10800 6246
rect 13916 12348 13972 12404
rect 13804 10722 13860 10724
rect 13804 10670 13806 10722
rect 13806 10670 13858 10722
rect 13858 10670 13860 10722
rect 13804 10668 13860 10670
rect 13580 10556 13636 10612
rect 13916 10332 13972 10388
rect 12460 10108 12516 10164
rect 15148 15202 15204 15204
rect 15148 15150 15150 15202
rect 15150 15150 15202 15202
rect 15202 15150 15204 15202
rect 15148 15148 15204 15150
rect 15372 15148 15428 15204
rect 15198 14922 15254 14924
rect 15198 14870 15200 14922
rect 15200 14870 15252 14922
rect 15252 14870 15254 14922
rect 15198 14868 15254 14870
rect 15302 14922 15358 14924
rect 15302 14870 15304 14922
rect 15304 14870 15356 14922
rect 15356 14870 15358 14922
rect 15302 14868 15358 14870
rect 15406 14922 15462 14924
rect 15406 14870 15408 14922
rect 15408 14870 15460 14922
rect 15460 14870 15462 14922
rect 15406 14868 15462 14870
rect 14812 14476 14868 14532
rect 15198 13354 15254 13356
rect 15198 13302 15200 13354
rect 15200 13302 15252 13354
rect 15252 13302 15254 13354
rect 15198 13300 15254 13302
rect 15302 13354 15358 13356
rect 15302 13302 15304 13354
rect 15304 13302 15356 13354
rect 15356 13302 15358 13354
rect 15302 13300 15358 13302
rect 15406 13354 15462 13356
rect 15406 13302 15408 13354
rect 15408 13302 15460 13354
rect 15460 13302 15462 13354
rect 15406 13300 15462 13302
rect 15198 11786 15254 11788
rect 15198 11734 15200 11786
rect 15200 11734 15252 11786
rect 15252 11734 15254 11786
rect 15198 11732 15254 11734
rect 15302 11786 15358 11788
rect 15302 11734 15304 11786
rect 15304 11734 15356 11786
rect 15356 11734 15358 11786
rect 15302 11732 15358 11734
rect 15406 11786 15462 11788
rect 15406 11734 15408 11786
rect 15408 11734 15460 11786
rect 15460 11734 15462 11786
rect 15406 11732 15462 11734
rect 17612 20188 17668 20244
rect 17276 20018 17332 20020
rect 17276 19966 17278 20018
rect 17278 19966 17330 20018
rect 17330 19966 17332 20018
rect 17276 19964 17332 19966
rect 16716 17052 16772 17108
rect 16828 18284 16884 18340
rect 15708 15260 15764 15316
rect 17948 21196 18004 21252
rect 19404 21196 19460 21252
rect 20412 23266 20468 23268
rect 20412 23214 20414 23266
rect 20414 23214 20466 23266
rect 20466 23214 20468 23266
rect 20412 23212 20468 23214
rect 21868 24892 21924 24948
rect 24522 27466 24578 27468
rect 24522 27414 24524 27466
rect 24524 27414 24576 27466
rect 24576 27414 24578 27466
rect 24522 27412 24578 27414
rect 24626 27466 24682 27468
rect 24626 27414 24628 27466
rect 24628 27414 24680 27466
rect 24680 27414 24682 27466
rect 24626 27412 24682 27414
rect 24730 27466 24786 27468
rect 24730 27414 24732 27466
rect 24732 27414 24784 27466
rect 24784 27414 24786 27466
rect 24730 27412 24786 27414
rect 25788 27468 25844 27524
rect 24668 26290 24724 26292
rect 24668 26238 24670 26290
rect 24670 26238 24722 26290
rect 24722 26238 24724 26290
rect 24668 26236 24724 26238
rect 25340 26290 25396 26292
rect 25340 26238 25342 26290
rect 25342 26238 25394 26290
rect 25394 26238 25396 26290
rect 25340 26236 25396 26238
rect 24522 25898 24578 25900
rect 24522 25846 24524 25898
rect 24524 25846 24576 25898
rect 24576 25846 24578 25898
rect 24522 25844 24578 25846
rect 24626 25898 24682 25900
rect 24626 25846 24628 25898
rect 24628 25846 24680 25898
rect 24680 25846 24682 25898
rect 24626 25844 24682 25846
rect 24730 25898 24786 25900
rect 24730 25846 24732 25898
rect 24732 25846 24784 25898
rect 24784 25846 24786 25898
rect 24730 25844 24786 25846
rect 22428 25618 22484 25620
rect 22428 25566 22430 25618
rect 22430 25566 22482 25618
rect 22482 25566 22484 25618
rect 22428 25564 22484 25566
rect 23996 25564 24052 25620
rect 23548 25394 23604 25396
rect 23548 25342 23550 25394
rect 23550 25342 23602 25394
rect 23602 25342 23604 25394
rect 23548 25340 23604 25342
rect 22204 24722 22260 24724
rect 22204 24670 22206 24722
rect 22206 24670 22258 24722
rect 22258 24670 22260 24722
rect 22204 24668 22260 24670
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 19740 22146 19796 22148
rect 19740 22094 19742 22146
rect 19742 22094 19794 22146
rect 19794 22094 19796 22146
rect 19740 22092 19796 22094
rect 19860 21978 19916 21980
rect 19860 21926 19862 21978
rect 19862 21926 19914 21978
rect 19914 21926 19916 21978
rect 19860 21924 19916 21926
rect 19964 21978 20020 21980
rect 19964 21926 19966 21978
rect 19966 21926 20018 21978
rect 20018 21926 20020 21978
rect 19964 21924 20020 21926
rect 20068 21978 20124 21980
rect 20068 21926 20070 21978
rect 20070 21926 20122 21978
rect 20122 21926 20124 21978
rect 20068 21924 20124 21926
rect 19860 20410 19916 20412
rect 19860 20358 19862 20410
rect 19862 20358 19914 20410
rect 19914 20358 19916 20410
rect 19860 20356 19916 20358
rect 19964 20410 20020 20412
rect 19964 20358 19966 20410
rect 19966 20358 20018 20410
rect 20018 20358 20020 20410
rect 19964 20356 20020 20358
rect 20068 20410 20124 20412
rect 20068 20358 20070 20410
rect 20070 20358 20122 20410
rect 20122 20358 20124 20410
rect 20068 20356 20124 20358
rect 20636 21532 20692 21588
rect 21308 21532 21364 21588
rect 23436 24668 23492 24724
rect 25228 24892 25284 24948
rect 25564 25618 25620 25620
rect 25564 25566 25566 25618
rect 25566 25566 25618 25618
rect 25618 25566 25620 25618
rect 25564 25564 25620 25566
rect 25340 24668 25396 24724
rect 24522 24330 24578 24332
rect 24522 24278 24524 24330
rect 24524 24278 24576 24330
rect 24576 24278 24578 24330
rect 24522 24276 24578 24278
rect 24626 24330 24682 24332
rect 24626 24278 24628 24330
rect 24628 24278 24680 24330
rect 24680 24278 24682 24330
rect 24626 24276 24682 24278
rect 24730 24330 24786 24332
rect 24730 24278 24732 24330
rect 24732 24278 24784 24330
rect 24784 24278 24786 24330
rect 24730 24276 24786 24278
rect 24780 24108 24836 24164
rect 24220 23378 24276 23380
rect 24220 23326 24222 23378
rect 24222 23326 24274 23378
rect 24274 23326 24276 23378
rect 24220 23324 24276 23326
rect 25564 23884 25620 23940
rect 26572 24108 26628 24164
rect 27132 28700 27188 28756
rect 28028 28530 28084 28532
rect 28028 28478 28030 28530
rect 28030 28478 28082 28530
rect 28082 28478 28084 28530
rect 28028 28476 28084 28478
rect 29932 28812 29988 28868
rect 28476 27692 28532 27748
rect 28812 28476 28868 28532
rect 27020 27468 27076 27524
rect 27580 26908 27636 26964
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 29596 28252 29652 28308
rect 29148 26962 29204 26964
rect 29148 26910 29150 26962
rect 29150 26910 29202 26962
rect 29202 26910 29204 26962
rect 29148 26908 29204 26910
rect 29184 26682 29240 26684
rect 29184 26630 29186 26682
rect 29186 26630 29238 26682
rect 29238 26630 29240 26682
rect 29184 26628 29240 26630
rect 29288 26682 29344 26684
rect 29288 26630 29290 26682
rect 29290 26630 29342 26682
rect 29342 26630 29344 26682
rect 29288 26628 29344 26630
rect 29392 26682 29448 26684
rect 29392 26630 29394 26682
rect 29394 26630 29446 26682
rect 29446 26630 29448 26682
rect 29392 26628 29448 26630
rect 30156 28754 30212 28756
rect 30156 28702 30158 28754
rect 30158 28702 30210 28754
rect 30210 28702 30212 28754
rect 30156 28700 30212 28702
rect 32060 28812 32116 28868
rect 31164 28530 31220 28532
rect 31164 28478 31166 28530
rect 31166 28478 31218 28530
rect 31218 28478 31220 28530
rect 31164 28476 31220 28478
rect 31052 28252 31108 28308
rect 29708 27020 29764 27076
rect 29260 25506 29316 25508
rect 29260 25454 29262 25506
rect 29262 25454 29314 25506
rect 29314 25454 29316 25506
rect 29260 25452 29316 25454
rect 26684 24722 26740 24724
rect 26684 24670 26686 24722
rect 26686 24670 26738 24722
rect 26738 24670 26740 24722
rect 26684 24668 26740 24670
rect 26236 23884 26292 23940
rect 26460 23772 26516 23828
rect 21868 23100 21924 23156
rect 27132 23996 27188 24052
rect 31164 26850 31220 26852
rect 31164 26798 31166 26850
rect 31166 26798 31218 26850
rect 31218 26798 31220 26850
rect 31164 26796 31220 26798
rect 30156 26684 30212 26740
rect 29184 25114 29240 25116
rect 29184 25062 29186 25114
rect 29186 25062 29238 25114
rect 29238 25062 29240 25114
rect 29184 25060 29240 25062
rect 29288 25114 29344 25116
rect 29288 25062 29290 25114
rect 29290 25062 29342 25114
rect 29342 25062 29344 25114
rect 29288 25060 29344 25062
rect 29392 25114 29448 25116
rect 29392 25062 29394 25114
rect 29394 25062 29446 25114
rect 29446 25062 29448 25114
rect 29392 25060 29448 25062
rect 29596 24946 29652 24948
rect 29596 24894 29598 24946
rect 29598 24894 29650 24946
rect 29650 24894 29652 24946
rect 29596 24892 29652 24894
rect 34076 33234 34132 33236
rect 34076 33182 34078 33234
rect 34078 33182 34130 33234
rect 34130 33182 34132 33234
rect 34076 33180 34132 33182
rect 33846 32170 33902 32172
rect 33846 32118 33848 32170
rect 33848 32118 33900 32170
rect 33900 32118 33902 32170
rect 33846 32116 33902 32118
rect 33950 32170 34006 32172
rect 33950 32118 33952 32170
rect 33952 32118 34004 32170
rect 34004 32118 34006 32170
rect 33950 32116 34006 32118
rect 34054 32170 34110 32172
rect 34054 32118 34056 32170
rect 34056 32118 34108 32170
rect 34108 32118 34110 32170
rect 34054 32116 34110 32118
rect 33846 30602 33902 30604
rect 33846 30550 33848 30602
rect 33848 30550 33900 30602
rect 33900 30550 33902 30602
rect 33846 30548 33902 30550
rect 33950 30602 34006 30604
rect 33950 30550 33952 30602
rect 33952 30550 34004 30602
rect 34004 30550 34006 30602
rect 33950 30548 34006 30550
rect 34054 30602 34110 30604
rect 34054 30550 34056 30602
rect 34056 30550 34108 30602
rect 34108 30550 34110 30602
rect 34054 30548 34110 30550
rect 33516 29372 33572 29428
rect 32732 28364 32788 28420
rect 32956 27020 33012 27076
rect 33180 28476 33236 28532
rect 33404 28140 33460 28196
rect 33180 26796 33236 26852
rect 33068 26236 33124 26292
rect 33068 25506 33124 25508
rect 33068 25454 33070 25506
rect 33070 25454 33122 25506
rect 33122 25454 33124 25506
rect 33068 25452 33124 25454
rect 30492 24946 30548 24948
rect 30492 24894 30494 24946
rect 30494 24894 30546 24946
rect 30546 24894 30548 24946
rect 30492 24892 30548 24894
rect 34524 33516 34580 33572
rect 34412 31052 34468 31108
rect 34300 29372 34356 29428
rect 33846 29034 33902 29036
rect 33846 28982 33848 29034
rect 33848 28982 33900 29034
rect 33900 28982 33902 29034
rect 33846 28980 33902 28982
rect 33950 29034 34006 29036
rect 33950 28982 33952 29034
rect 33952 28982 34004 29034
rect 34004 28982 34006 29034
rect 33950 28980 34006 28982
rect 34054 29034 34110 29036
rect 34054 28982 34056 29034
rect 34056 28982 34108 29034
rect 34108 28982 34110 29034
rect 34054 28980 34110 28982
rect 33846 27466 33902 27468
rect 33846 27414 33848 27466
rect 33848 27414 33900 27466
rect 33900 27414 33902 27466
rect 33846 27412 33902 27414
rect 33950 27466 34006 27468
rect 33950 27414 33952 27466
rect 33952 27414 34004 27466
rect 34004 27414 34006 27466
rect 33950 27412 34006 27414
rect 34054 27466 34110 27468
rect 34054 27414 34056 27466
rect 34056 27414 34108 27466
rect 34108 27414 34110 27466
rect 34054 27412 34110 27414
rect 34412 28140 34468 28196
rect 34188 26684 34244 26740
rect 34076 26236 34132 26292
rect 33846 25898 33902 25900
rect 33846 25846 33848 25898
rect 33848 25846 33900 25898
rect 33900 25846 33902 25898
rect 33846 25844 33902 25846
rect 33950 25898 34006 25900
rect 33950 25846 33952 25898
rect 33952 25846 34004 25898
rect 34004 25846 34006 25898
rect 33950 25844 34006 25846
rect 34054 25898 34110 25900
rect 34054 25846 34056 25898
rect 34056 25846 34108 25898
rect 34108 25846 34110 25898
rect 34054 25844 34110 25846
rect 33852 25228 33908 25284
rect 31948 24668 32004 24724
rect 33404 24722 33460 24724
rect 33404 24670 33406 24722
rect 33406 24670 33458 24722
rect 33458 24670 33460 24722
rect 33404 24668 33460 24670
rect 27580 23884 27636 23940
rect 27244 23826 27300 23828
rect 27244 23774 27246 23826
rect 27246 23774 27298 23826
rect 27298 23774 27300 23826
rect 27244 23772 27300 23774
rect 28252 23938 28308 23940
rect 28252 23886 28254 23938
rect 28254 23886 28306 23938
rect 28306 23886 28308 23938
rect 28252 23884 28308 23886
rect 27020 23714 27076 23716
rect 27020 23662 27022 23714
rect 27022 23662 27074 23714
rect 27074 23662 27076 23714
rect 27020 23660 27076 23662
rect 24522 22762 24578 22764
rect 24522 22710 24524 22762
rect 24524 22710 24576 22762
rect 24576 22710 24578 22762
rect 24522 22708 24578 22710
rect 24626 22762 24682 22764
rect 24626 22710 24628 22762
rect 24628 22710 24680 22762
rect 24680 22710 24682 22762
rect 24626 22708 24682 22710
rect 24730 22762 24786 22764
rect 24730 22710 24732 22762
rect 24732 22710 24784 22762
rect 24784 22710 24786 22762
rect 24730 22708 24786 22710
rect 25788 22764 25844 22820
rect 21756 22370 21812 22372
rect 21756 22318 21758 22370
rect 21758 22318 21810 22370
rect 21810 22318 21812 22370
rect 21756 22316 21812 22318
rect 22204 22428 22260 22484
rect 22764 22204 22820 22260
rect 23772 22092 23828 22148
rect 21532 20188 21588 20244
rect 21756 21420 21812 21476
rect 24668 21474 24724 21476
rect 24668 21422 24670 21474
rect 24670 21422 24722 21474
rect 24722 21422 24724 21474
rect 24668 21420 24724 21422
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 22316 20524 22372 20580
rect 22988 20578 23044 20580
rect 22988 20526 22990 20578
rect 22990 20526 23042 20578
rect 23042 20526 23044 20578
rect 22988 20524 23044 20526
rect 22092 19906 22148 19908
rect 22092 19854 22094 19906
rect 22094 19854 22146 19906
rect 22146 19854 22148 19906
rect 22092 19852 22148 19854
rect 23436 20132 23492 20188
rect 23212 19906 23268 19908
rect 23212 19854 23214 19906
rect 23214 19854 23266 19906
rect 23266 19854 23268 19906
rect 23212 19852 23268 19854
rect 22988 19180 23044 19236
rect 17388 18956 17444 19012
rect 19860 18842 19916 18844
rect 19860 18790 19862 18842
rect 19862 18790 19914 18842
rect 19914 18790 19916 18842
rect 19860 18788 19916 18790
rect 19964 18842 20020 18844
rect 19964 18790 19966 18842
rect 19966 18790 20018 18842
rect 20018 18790 20020 18842
rect 19964 18788 20020 18790
rect 20068 18842 20124 18844
rect 20068 18790 20070 18842
rect 20070 18790 20122 18842
rect 20122 18790 20124 18842
rect 20068 18788 20124 18790
rect 17052 18396 17108 18452
rect 18956 18450 19012 18452
rect 18956 18398 18958 18450
rect 18958 18398 19010 18450
rect 19010 18398 19012 18450
rect 18956 18396 19012 18398
rect 17612 18338 17668 18340
rect 17612 18286 17614 18338
rect 17614 18286 17666 18338
rect 17666 18286 17668 18338
rect 17612 18284 17668 18286
rect 18060 18338 18116 18340
rect 18060 18286 18062 18338
rect 18062 18286 18114 18338
rect 18114 18286 18116 18338
rect 18060 18284 18116 18286
rect 16940 17836 16996 17892
rect 17948 17836 18004 17892
rect 20636 18284 20692 18340
rect 19404 17612 19460 17668
rect 16380 16098 16436 16100
rect 16380 16046 16382 16098
rect 16382 16046 16434 16098
rect 16434 16046 16436 16098
rect 16380 16044 16436 16046
rect 16044 15314 16100 15316
rect 16044 15262 16046 15314
rect 16046 15262 16098 15314
rect 16098 15262 16100 15314
rect 16044 15260 16100 15262
rect 16380 15148 16436 15204
rect 16828 14642 16884 14644
rect 16828 14590 16830 14642
rect 16830 14590 16882 14642
rect 16882 14590 16884 14642
rect 16828 14588 16884 14590
rect 16380 12236 16436 12292
rect 15708 11564 15764 11620
rect 14028 9884 14084 9940
rect 14924 10556 14980 10612
rect 14364 9324 14420 9380
rect 15596 10444 15652 10500
rect 15198 10218 15254 10220
rect 15198 10166 15200 10218
rect 15200 10166 15252 10218
rect 15252 10166 15254 10218
rect 15198 10164 15254 10166
rect 15302 10218 15358 10220
rect 15302 10166 15304 10218
rect 15304 10166 15356 10218
rect 15356 10166 15358 10218
rect 15302 10164 15358 10166
rect 15406 10218 15462 10220
rect 15406 10166 15408 10218
rect 15408 10166 15460 10218
rect 15460 10166 15462 10218
rect 15406 10164 15462 10166
rect 18956 16156 19012 16212
rect 19292 15932 19348 15988
rect 17836 15260 17892 15316
rect 17500 15202 17556 15204
rect 17500 15150 17502 15202
rect 17502 15150 17554 15202
rect 17554 15150 17556 15202
rect 17500 15148 17556 15150
rect 17164 14812 17220 14868
rect 17276 14588 17332 14644
rect 17052 12908 17108 12964
rect 16940 12124 16996 12180
rect 16940 11564 16996 11620
rect 15932 10332 15988 10388
rect 15036 9042 15092 9044
rect 15036 8990 15038 9042
rect 15038 8990 15090 9042
rect 15090 8990 15092 9042
rect 15036 8988 15092 8990
rect 15198 8650 15254 8652
rect 15198 8598 15200 8650
rect 15200 8598 15252 8650
rect 15252 8598 15254 8650
rect 15198 8596 15254 8598
rect 15302 8650 15358 8652
rect 15302 8598 15304 8650
rect 15304 8598 15356 8650
rect 15356 8598 15358 8650
rect 15302 8596 15358 8598
rect 15406 8650 15462 8652
rect 15406 8598 15408 8650
rect 15408 8598 15460 8650
rect 15460 8598 15462 8650
rect 15406 8596 15462 8598
rect 16492 10610 16548 10612
rect 16492 10558 16494 10610
rect 16494 10558 16546 10610
rect 16546 10558 16548 10610
rect 16492 10556 16548 10558
rect 17724 12290 17780 12292
rect 17724 12238 17726 12290
rect 17726 12238 17778 12290
rect 17778 12238 17780 12290
rect 17724 12236 17780 12238
rect 17948 13020 18004 13076
rect 17948 12850 18004 12852
rect 17948 12798 17950 12850
rect 17950 12798 18002 12850
rect 18002 12798 18004 12850
rect 17948 12796 18004 12798
rect 17388 10892 17444 10948
rect 17948 12012 18004 12068
rect 17388 10722 17444 10724
rect 17388 10670 17390 10722
rect 17390 10670 17442 10722
rect 17442 10670 17444 10722
rect 17388 10668 17444 10670
rect 19292 14588 19348 14644
rect 18620 13020 18676 13076
rect 18284 12908 18340 12964
rect 18172 11116 18228 11172
rect 17612 10444 17668 10500
rect 18284 10668 18340 10724
rect 14700 7420 14756 7476
rect 15708 7420 15764 7476
rect 13356 7362 13412 7364
rect 13356 7310 13358 7362
rect 13358 7310 13410 7362
rect 13410 7310 13412 7362
rect 13356 7308 13412 7310
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 18844 12124 18900 12180
rect 18732 12066 18788 12068
rect 18732 12014 18734 12066
rect 18734 12014 18786 12066
rect 18786 12014 18788 12066
rect 18732 12012 18788 12014
rect 19068 11564 19124 11620
rect 19292 11228 19348 11284
rect 20188 17666 20244 17668
rect 20188 17614 20190 17666
rect 20190 17614 20242 17666
rect 20242 17614 20244 17666
rect 20188 17612 20244 17614
rect 19860 17274 19916 17276
rect 19860 17222 19862 17274
rect 19862 17222 19914 17274
rect 19914 17222 19916 17274
rect 19860 17220 19916 17222
rect 19964 17274 20020 17276
rect 19964 17222 19966 17274
rect 19966 17222 20018 17274
rect 20018 17222 20020 17274
rect 19964 17220 20020 17222
rect 20068 17274 20124 17276
rect 20068 17222 20070 17274
rect 20070 17222 20122 17274
rect 20122 17222 20124 17274
rect 20068 17220 20124 17222
rect 21980 17164 22036 17220
rect 20636 16882 20692 16884
rect 20636 16830 20638 16882
rect 20638 16830 20690 16882
rect 20690 16830 20692 16882
rect 20636 16828 20692 16830
rect 21084 16044 21140 16100
rect 21532 16828 21588 16884
rect 20076 15986 20132 15988
rect 20076 15934 20078 15986
rect 20078 15934 20130 15986
rect 20130 15934 20132 15986
rect 20076 15932 20132 15934
rect 19516 15148 19572 15204
rect 19516 14476 19572 14532
rect 19516 11564 19572 11620
rect 19860 15706 19916 15708
rect 19860 15654 19862 15706
rect 19862 15654 19914 15706
rect 19914 15654 19916 15706
rect 19860 15652 19916 15654
rect 19964 15706 20020 15708
rect 19964 15654 19966 15706
rect 19966 15654 20018 15706
rect 20018 15654 20020 15706
rect 19964 15652 20020 15654
rect 20068 15706 20124 15708
rect 20068 15654 20070 15706
rect 20070 15654 20122 15706
rect 20122 15654 20124 15706
rect 20068 15652 20124 15654
rect 20412 15260 20468 15316
rect 19964 14642 20020 14644
rect 19964 14590 19966 14642
rect 19966 14590 20018 14642
rect 20018 14590 20020 14642
rect 19964 14588 20020 14590
rect 20748 14252 20804 14308
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 20412 13244 20468 13300
rect 19860 12570 19916 12572
rect 19860 12518 19862 12570
rect 19862 12518 19914 12570
rect 19914 12518 19916 12570
rect 19860 12516 19916 12518
rect 19964 12570 20020 12572
rect 19964 12518 19966 12570
rect 19966 12518 20018 12570
rect 20018 12518 20020 12570
rect 19964 12516 20020 12518
rect 20068 12570 20124 12572
rect 20068 12518 20070 12570
rect 20070 12518 20122 12570
rect 20122 12518 20124 12570
rect 20068 12516 20124 12518
rect 19628 11228 19684 11284
rect 19628 10892 19684 10948
rect 19292 9938 19348 9940
rect 19292 9886 19294 9938
rect 19294 9886 19346 9938
rect 19346 9886 19348 9938
rect 19292 9884 19348 9886
rect 20188 11452 20244 11508
rect 19860 11002 19916 11004
rect 19860 10950 19862 11002
rect 19862 10950 19914 11002
rect 19914 10950 19916 11002
rect 19860 10948 19916 10950
rect 19964 11002 20020 11004
rect 19964 10950 19966 11002
rect 19966 10950 20018 11002
rect 20018 10950 20020 11002
rect 19964 10948 20020 10950
rect 20068 11002 20124 11004
rect 20068 10950 20070 11002
rect 20070 10950 20122 11002
rect 20122 10950 20124 11002
rect 20068 10948 20124 10950
rect 20188 10722 20244 10724
rect 20188 10670 20190 10722
rect 20190 10670 20242 10722
rect 20242 10670 20244 10722
rect 20188 10668 20244 10670
rect 19740 10444 19796 10500
rect 20636 11170 20692 11172
rect 20636 11118 20638 11170
rect 20638 11118 20690 11170
rect 20690 11118 20692 11170
rect 20636 11116 20692 11118
rect 20300 9996 20356 10052
rect 21308 13916 21364 13972
rect 21644 16210 21700 16212
rect 21644 16158 21646 16210
rect 21646 16158 21698 16210
rect 21698 16158 21700 16210
rect 21644 16156 21700 16158
rect 22204 16828 22260 16884
rect 23212 18338 23268 18340
rect 23212 18286 23214 18338
rect 23214 18286 23266 18338
rect 23266 18286 23268 18338
rect 23212 18284 23268 18286
rect 22876 17836 22932 17892
rect 22876 17052 22932 17108
rect 23436 16716 23492 16772
rect 23100 16044 23156 16100
rect 22764 15538 22820 15540
rect 22764 15486 22766 15538
rect 22766 15486 22818 15538
rect 22818 15486 22820 15538
rect 22764 15484 22820 15486
rect 22652 15372 22708 15428
rect 23660 15484 23716 15540
rect 24220 20578 24276 20580
rect 24220 20526 24222 20578
rect 24222 20526 24274 20578
rect 24274 20526 24276 20578
rect 24220 20524 24276 20526
rect 25564 22146 25620 22148
rect 25564 22094 25566 22146
rect 25566 22094 25618 22146
rect 25618 22094 25620 22146
rect 25564 22092 25620 22094
rect 25340 21586 25396 21588
rect 25340 21534 25342 21586
rect 25342 21534 25394 21586
rect 25394 21534 25396 21586
rect 25340 21532 25396 21534
rect 26460 22482 26516 22484
rect 26460 22430 26462 22482
rect 26462 22430 26514 22482
rect 26514 22430 26516 22482
rect 26460 22428 26516 22430
rect 27468 22258 27524 22260
rect 27468 22206 27470 22258
rect 27470 22206 27522 22258
rect 27522 22206 27524 22258
rect 27468 22204 27524 22206
rect 26908 21532 26964 21588
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 26012 19794 26068 19796
rect 26012 19742 26014 19794
rect 26014 19742 26066 19794
rect 26066 19742 26068 19794
rect 26012 19740 26068 19742
rect 24522 19626 24578 19628
rect 24522 19574 24524 19626
rect 24524 19574 24576 19626
rect 24576 19574 24578 19626
rect 24522 19572 24578 19574
rect 24626 19626 24682 19628
rect 24626 19574 24628 19626
rect 24628 19574 24680 19626
rect 24680 19574 24682 19626
rect 24626 19572 24682 19574
rect 24730 19626 24786 19628
rect 24730 19574 24732 19626
rect 24732 19574 24784 19626
rect 24784 19574 24786 19626
rect 24730 19572 24786 19574
rect 23884 18338 23940 18340
rect 23884 18286 23886 18338
rect 23886 18286 23938 18338
rect 23938 18286 23940 18338
rect 23884 18284 23940 18286
rect 24522 18058 24578 18060
rect 24522 18006 24524 18058
rect 24524 18006 24576 18058
rect 24576 18006 24578 18058
rect 24522 18004 24578 18006
rect 24626 18058 24682 18060
rect 24626 18006 24628 18058
rect 24628 18006 24680 18058
rect 24680 18006 24682 18058
rect 24626 18004 24682 18006
rect 24730 18058 24786 18060
rect 24730 18006 24732 18058
rect 24732 18006 24784 18058
rect 24784 18006 24786 18058
rect 24730 18004 24786 18006
rect 29184 23546 29240 23548
rect 29184 23494 29186 23546
rect 29186 23494 29238 23546
rect 29238 23494 29240 23546
rect 29184 23492 29240 23494
rect 29288 23546 29344 23548
rect 29288 23494 29290 23546
rect 29290 23494 29342 23546
rect 29342 23494 29344 23546
rect 29288 23492 29344 23494
rect 29392 23546 29448 23548
rect 29392 23494 29394 23546
rect 29394 23494 29446 23546
rect 29446 23494 29448 23546
rect 29392 23492 29448 23494
rect 28364 23324 28420 23380
rect 28812 22876 28868 22932
rect 28588 22316 28644 22372
rect 27580 21420 27636 21476
rect 29260 22204 29316 22260
rect 32956 24050 33012 24052
rect 32956 23998 32958 24050
rect 32958 23998 33010 24050
rect 33010 23998 33012 24050
rect 32956 23996 33012 23998
rect 30380 23884 30436 23940
rect 31164 23660 31220 23716
rect 33180 23154 33236 23156
rect 33180 23102 33182 23154
rect 33182 23102 33234 23154
rect 33234 23102 33236 23154
rect 33180 23100 33236 23102
rect 30156 22764 30212 22820
rect 29484 22316 29540 22372
rect 29372 22092 29428 22148
rect 29820 22204 29876 22260
rect 29184 21978 29240 21980
rect 29184 21926 29186 21978
rect 29186 21926 29238 21978
rect 29238 21926 29240 21978
rect 29184 21924 29240 21926
rect 29288 21978 29344 21980
rect 29288 21926 29290 21978
rect 29290 21926 29342 21978
rect 29342 21926 29344 21978
rect 29288 21924 29344 21926
rect 29392 21978 29448 21980
rect 29392 21926 29394 21978
rect 29394 21926 29446 21978
rect 29446 21926 29448 21978
rect 29392 21924 29448 21926
rect 28476 21420 28532 21476
rect 29596 21586 29652 21588
rect 29596 21534 29598 21586
rect 29598 21534 29650 21586
rect 29650 21534 29652 21586
rect 29596 21532 29652 21534
rect 28924 20748 28980 20804
rect 26796 20636 26852 20692
rect 28252 20690 28308 20692
rect 28252 20638 28254 20690
rect 28254 20638 28306 20690
rect 28306 20638 28308 20690
rect 28252 20636 28308 20638
rect 28588 20690 28644 20692
rect 28588 20638 28590 20690
rect 28590 20638 28642 20690
rect 28642 20638 28644 20690
rect 28588 20636 28644 20638
rect 27356 20524 27412 20580
rect 30828 22258 30884 22260
rect 30828 22206 30830 22258
rect 30830 22206 30882 22258
rect 30882 22206 30884 22258
rect 30828 22204 30884 22206
rect 31164 22092 31220 22148
rect 32060 21644 32116 21700
rect 33068 21698 33124 21700
rect 33068 21646 33070 21698
rect 33070 21646 33122 21698
rect 33122 21646 33124 21698
rect 33068 21644 33124 21646
rect 31724 21420 31780 21476
rect 29184 20410 29240 20412
rect 29184 20358 29186 20410
rect 29186 20358 29238 20410
rect 29238 20358 29240 20410
rect 29184 20356 29240 20358
rect 29288 20410 29344 20412
rect 29288 20358 29290 20410
rect 29290 20358 29342 20410
rect 29342 20358 29344 20410
rect 29288 20356 29344 20358
rect 29392 20410 29448 20412
rect 29392 20358 29394 20410
rect 29394 20358 29446 20410
rect 29446 20358 29448 20410
rect 29392 20356 29448 20358
rect 26572 18956 26628 19012
rect 26908 19852 26964 19908
rect 26460 18844 26516 18900
rect 23884 17164 23940 17220
rect 24668 17164 24724 17220
rect 24108 16994 24164 16996
rect 24108 16942 24110 16994
rect 24110 16942 24162 16994
rect 24162 16942 24164 16994
rect 24108 16940 24164 16942
rect 25564 17164 25620 17220
rect 26012 16882 26068 16884
rect 26012 16830 26014 16882
rect 26014 16830 26066 16882
rect 26066 16830 26068 16882
rect 26012 16828 26068 16830
rect 24220 15874 24276 15876
rect 24220 15822 24222 15874
rect 24222 15822 24274 15874
rect 24274 15822 24276 15874
rect 24220 15820 24276 15822
rect 24108 15426 24164 15428
rect 24108 15374 24110 15426
rect 24110 15374 24162 15426
rect 24162 15374 24164 15426
rect 24108 15372 24164 15374
rect 23772 15148 23828 15204
rect 23660 14306 23716 14308
rect 23660 14254 23662 14306
rect 23662 14254 23714 14306
rect 23714 14254 23716 14306
rect 23660 14252 23716 14254
rect 24522 16490 24578 16492
rect 24522 16438 24524 16490
rect 24524 16438 24576 16490
rect 24576 16438 24578 16490
rect 24522 16436 24578 16438
rect 24626 16490 24682 16492
rect 24626 16438 24628 16490
rect 24628 16438 24680 16490
rect 24680 16438 24682 16490
rect 24626 16436 24682 16438
rect 24730 16490 24786 16492
rect 24730 16438 24732 16490
rect 24732 16438 24784 16490
rect 24784 16438 24786 16490
rect 24730 16436 24786 16438
rect 24522 14922 24578 14924
rect 24522 14870 24524 14922
rect 24524 14870 24576 14922
rect 24576 14870 24578 14922
rect 24522 14868 24578 14870
rect 24626 14922 24682 14924
rect 24626 14870 24628 14922
rect 24628 14870 24680 14922
rect 24680 14870 24682 14922
rect 24626 14868 24682 14870
rect 24730 14922 24786 14924
rect 24730 14870 24732 14922
rect 24732 14870 24784 14922
rect 24784 14870 24786 14922
rect 24730 14868 24786 14870
rect 22316 13916 22372 13972
rect 20972 13132 21028 13188
rect 21084 12908 21140 12964
rect 21532 12850 21588 12852
rect 21532 12798 21534 12850
rect 21534 12798 21586 12850
rect 21586 12798 21588 12850
rect 21532 12796 21588 12798
rect 22204 13074 22260 13076
rect 22204 13022 22206 13074
rect 22206 13022 22258 13074
rect 22258 13022 22260 13074
rect 22204 13020 22260 13022
rect 21756 12572 21812 12628
rect 21532 12236 21588 12292
rect 23212 13468 23268 13524
rect 22876 13132 22932 13188
rect 22428 12796 22484 12852
rect 22428 11452 22484 11508
rect 21980 10498 22036 10500
rect 21980 10446 21982 10498
rect 21982 10446 22034 10498
rect 22034 10446 22036 10498
rect 21980 10444 22036 10446
rect 23324 13244 23380 13300
rect 23212 12962 23268 12964
rect 23212 12910 23214 12962
rect 23214 12910 23266 12962
rect 23266 12910 23268 12962
rect 23212 12908 23268 12910
rect 23324 12796 23380 12852
rect 22988 11564 23044 11620
rect 23548 11282 23604 11284
rect 23548 11230 23550 11282
rect 23550 11230 23602 11282
rect 23602 11230 23604 11282
rect 23548 11228 23604 11230
rect 24522 13354 24578 13356
rect 24522 13302 24524 13354
rect 24524 13302 24576 13354
rect 24576 13302 24578 13354
rect 24522 13300 24578 13302
rect 24626 13354 24682 13356
rect 24626 13302 24628 13354
rect 24628 13302 24680 13354
rect 24680 13302 24682 13354
rect 24626 13300 24682 13302
rect 24730 13354 24786 13356
rect 24730 13302 24732 13354
rect 24732 13302 24784 13354
rect 24784 13302 24786 13354
rect 24730 13300 24786 13302
rect 24556 12290 24612 12292
rect 24556 12238 24558 12290
rect 24558 12238 24610 12290
rect 24610 12238 24612 12290
rect 24556 12236 24612 12238
rect 25228 13468 25284 13524
rect 24892 12012 24948 12068
rect 25116 12572 25172 12628
rect 24522 11786 24578 11788
rect 24522 11734 24524 11786
rect 24524 11734 24576 11786
rect 24576 11734 24578 11786
rect 24522 11732 24578 11734
rect 24626 11786 24682 11788
rect 24626 11734 24628 11786
rect 24628 11734 24680 11786
rect 24680 11734 24682 11786
rect 24626 11732 24682 11734
rect 24730 11786 24786 11788
rect 24730 11734 24732 11786
rect 24732 11734 24784 11786
rect 24784 11734 24786 11786
rect 24730 11732 24786 11734
rect 25564 12236 25620 12292
rect 25788 13468 25844 13524
rect 26348 16828 26404 16884
rect 27916 19234 27972 19236
rect 27916 19182 27918 19234
rect 27918 19182 27970 19234
rect 27970 19182 27972 19234
rect 27916 19180 27972 19182
rect 27356 18956 27412 19012
rect 27580 17164 27636 17220
rect 26684 16828 26740 16884
rect 26572 14028 26628 14084
rect 26124 13356 26180 13412
rect 25788 12124 25844 12180
rect 26124 11564 26180 11620
rect 23884 10444 23940 10500
rect 26236 10498 26292 10500
rect 26236 10446 26238 10498
rect 26238 10446 26290 10498
rect 26290 10446 26292 10498
rect 26236 10444 26292 10446
rect 24522 10218 24578 10220
rect 24522 10166 24524 10218
rect 24524 10166 24576 10218
rect 24576 10166 24578 10218
rect 24522 10164 24578 10166
rect 24626 10218 24682 10220
rect 24626 10166 24628 10218
rect 24628 10166 24680 10218
rect 24680 10166 24682 10218
rect 24626 10164 24682 10166
rect 24730 10218 24786 10220
rect 24730 10166 24732 10218
rect 24732 10166 24784 10218
rect 24784 10166 24786 10218
rect 24730 10164 24786 10166
rect 23548 9996 23604 10052
rect 19860 9434 19916 9436
rect 19860 9382 19862 9434
rect 19862 9382 19914 9434
rect 19914 9382 19916 9434
rect 19860 9380 19916 9382
rect 19964 9434 20020 9436
rect 19964 9382 19966 9434
rect 19966 9382 20018 9434
rect 20018 9382 20020 9434
rect 19964 9380 20020 9382
rect 20068 9434 20124 9436
rect 20068 9382 20070 9434
rect 20070 9382 20122 9434
rect 20122 9382 20124 9434
rect 20068 9380 20124 9382
rect 24522 8650 24578 8652
rect 24522 8598 24524 8650
rect 24524 8598 24576 8650
rect 24576 8598 24578 8650
rect 24522 8596 24578 8598
rect 24626 8650 24682 8652
rect 24626 8598 24628 8650
rect 24628 8598 24680 8650
rect 24680 8598 24682 8650
rect 24626 8596 24682 8598
rect 24730 8650 24786 8652
rect 24730 8598 24732 8650
rect 24732 8598 24784 8650
rect 24784 8598 24786 8650
rect 24730 8596 24786 8598
rect 19860 7866 19916 7868
rect 19860 7814 19862 7866
rect 19862 7814 19914 7866
rect 19914 7814 19916 7866
rect 19860 7812 19916 7814
rect 19964 7866 20020 7868
rect 19964 7814 19966 7866
rect 19966 7814 20018 7866
rect 20018 7814 20020 7866
rect 19964 7812 20020 7814
rect 20068 7866 20124 7868
rect 20068 7814 20070 7866
rect 20070 7814 20122 7866
rect 20122 7814 20124 7866
rect 20068 7812 20124 7814
rect 19860 6298 19916 6300
rect 19860 6246 19862 6298
rect 19862 6246 19914 6298
rect 19914 6246 19916 6298
rect 19860 6244 19916 6246
rect 19964 6298 20020 6300
rect 19964 6246 19966 6298
rect 19966 6246 20018 6298
rect 20018 6246 20020 6298
rect 19964 6244 20020 6246
rect 20068 6298 20124 6300
rect 20068 6246 20070 6298
rect 20070 6246 20122 6298
rect 20122 6246 20124 6298
rect 20068 6244 20124 6246
rect 5874 5514 5930 5516
rect 5874 5462 5876 5514
rect 5876 5462 5928 5514
rect 5928 5462 5930 5514
rect 5874 5460 5930 5462
rect 5978 5514 6034 5516
rect 5978 5462 5980 5514
rect 5980 5462 6032 5514
rect 6032 5462 6034 5514
rect 5978 5460 6034 5462
rect 6082 5514 6138 5516
rect 6082 5462 6084 5514
rect 6084 5462 6136 5514
rect 6136 5462 6138 5514
rect 6082 5460 6138 5462
rect 15198 5514 15254 5516
rect 15198 5462 15200 5514
rect 15200 5462 15252 5514
rect 15252 5462 15254 5514
rect 15198 5460 15254 5462
rect 15302 5514 15358 5516
rect 15302 5462 15304 5514
rect 15304 5462 15356 5514
rect 15356 5462 15358 5514
rect 15302 5460 15358 5462
rect 15406 5514 15462 5516
rect 15406 5462 15408 5514
rect 15408 5462 15460 5514
rect 15460 5462 15462 5514
rect 15406 5460 15462 5462
rect 10536 4730 10592 4732
rect 10536 4678 10538 4730
rect 10538 4678 10590 4730
rect 10590 4678 10592 4730
rect 10536 4676 10592 4678
rect 10640 4730 10696 4732
rect 10640 4678 10642 4730
rect 10642 4678 10694 4730
rect 10694 4678 10696 4730
rect 10640 4676 10696 4678
rect 10744 4730 10800 4732
rect 10744 4678 10746 4730
rect 10746 4678 10798 4730
rect 10798 4678 10800 4730
rect 10744 4676 10800 4678
rect 19860 4730 19916 4732
rect 19860 4678 19862 4730
rect 19862 4678 19914 4730
rect 19914 4678 19916 4730
rect 19860 4676 19916 4678
rect 19964 4730 20020 4732
rect 19964 4678 19966 4730
rect 19966 4678 20018 4730
rect 20018 4678 20020 4730
rect 19964 4676 20020 4678
rect 20068 4730 20124 4732
rect 20068 4678 20070 4730
rect 20070 4678 20122 4730
rect 20122 4678 20124 4730
rect 20068 4676 20124 4678
rect 5874 3946 5930 3948
rect 5874 3894 5876 3946
rect 5876 3894 5928 3946
rect 5928 3894 5930 3946
rect 5874 3892 5930 3894
rect 5978 3946 6034 3948
rect 5978 3894 5980 3946
rect 5980 3894 6032 3946
rect 6032 3894 6034 3946
rect 5978 3892 6034 3894
rect 6082 3946 6138 3948
rect 6082 3894 6084 3946
rect 6084 3894 6136 3946
rect 6136 3894 6138 3946
rect 6082 3892 6138 3894
rect 15198 3946 15254 3948
rect 15198 3894 15200 3946
rect 15200 3894 15252 3946
rect 15252 3894 15254 3946
rect 15198 3892 15254 3894
rect 15302 3946 15358 3948
rect 15302 3894 15304 3946
rect 15304 3894 15356 3946
rect 15356 3894 15358 3946
rect 15302 3892 15358 3894
rect 15406 3946 15462 3948
rect 15406 3894 15408 3946
rect 15408 3894 15460 3946
rect 15460 3894 15462 3946
rect 15406 3892 15462 3894
rect 10536 3162 10592 3164
rect 10536 3110 10538 3162
rect 10538 3110 10590 3162
rect 10590 3110 10592 3162
rect 10536 3108 10592 3110
rect 10640 3162 10696 3164
rect 10640 3110 10642 3162
rect 10642 3110 10694 3162
rect 10694 3110 10696 3162
rect 10640 3108 10696 3110
rect 10744 3162 10800 3164
rect 10744 3110 10746 3162
rect 10746 3110 10798 3162
rect 10798 3110 10800 3162
rect 10744 3108 10800 3110
rect 19860 3162 19916 3164
rect 19860 3110 19862 3162
rect 19862 3110 19914 3162
rect 19914 3110 19916 3162
rect 19860 3108 19916 3110
rect 19964 3162 20020 3164
rect 19964 3110 19966 3162
rect 19966 3110 20018 3162
rect 20018 3110 20020 3162
rect 19964 3108 20020 3110
rect 20068 3162 20124 3164
rect 20068 3110 20070 3162
rect 20070 3110 20122 3162
rect 20122 3110 20124 3162
rect 20068 3108 20124 3110
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 26684 13468 26740 13524
rect 26348 6524 26404 6580
rect 26460 11564 26516 11620
rect 26572 11116 26628 11172
rect 28252 18172 28308 18228
rect 27692 15874 27748 15876
rect 27692 15822 27694 15874
rect 27694 15822 27746 15874
rect 27746 15822 27748 15874
rect 27692 15820 27748 15822
rect 27356 14028 27412 14084
rect 26908 11676 26964 11732
rect 27244 12012 27300 12068
rect 27580 12236 27636 12292
rect 27580 11564 27636 11620
rect 27244 10444 27300 10500
rect 26796 8876 26852 8932
rect 27020 10332 27076 10388
rect 29148 20018 29204 20020
rect 29148 19966 29150 20018
rect 29150 19966 29202 20018
rect 29202 19966 29204 20018
rect 29148 19964 29204 19966
rect 31052 20802 31108 20804
rect 31052 20750 31054 20802
rect 31054 20750 31106 20802
rect 31106 20750 31108 20802
rect 31052 20748 31108 20750
rect 30380 20690 30436 20692
rect 30380 20638 30382 20690
rect 30382 20638 30434 20690
rect 30434 20638 30436 20690
rect 30380 20636 30436 20638
rect 29820 20076 29876 20132
rect 30604 20130 30660 20132
rect 30604 20078 30606 20130
rect 30606 20078 30658 20130
rect 30658 20078 30660 20130
rect 30604 20076 30660 20078
rect 30940 19906 30996 19908
rect 30940 19854 30942 19906
rect 30942 19854 30994 19906
rect 30994 19854 30996 19906
rect 30940 19852 30996 19854
rect 29820 19292 29876 19348
rect 30380 19292 30436 19348
rect 28588 19234 28644 19236
rect 28588 19182 28590 19234
rect 28590 19182 28642 19234
rect 28642 19182 28644 19234
rect 28588 19180 28644 19182
rect 29260 19234 29316 19236
rect 29260 19182 29262 19234
rect 29262 19182 29314 19234
rect 29314 19182 29316 19234
rect 29260 19180 29316 19182
rect 29184 18842 29240 18844
rect 29184 18790 29186 18842
rect 29186 18790 29238 18842
rect 29238 18790 29240 18842
rect 29184 18788 29240 18790
rect 29288 18842 29344 18844
rect 29288 18790 29290 18842
rect 29290 18790 29342 18842
rect 29342 18790 29344 18842
rect 29288 18788 29344 18790
rect 29392 18842 29448 18844
rect 29392 18790 29394 18842
rect 29394 18790 29446 18842
rect 29446 18790 29448 18842
rect 29392 18788 29448 18790
rect 29184 17274 29240 17276
rect 29184 17222 29186 17274
rect 29186 17222 29238 17274
rect 29238 17222 29240 17274
rect 29184 17220 29240 17222
rect 29288 17274 29344 17276
rect 29288 17222 29290 17274
rect 29290 17222 29342 17274
rect 29342 17222 29344 17274
rect 29288 17220 29344 17222
rect 29392 17274 29448 17276
rect 29392 17222 29394 17274
rect 29394 17222 29446 17274
rect 29446 17222 29448 17274
rect 29392 17220 29448 17222
rect 29932 18226 29988 18228
rect 29932 18174 29934 18226
rect 29934 18174 29986 18226
rect 29986 18174 29988 18226
rect 29932 18172 29988 18174
rect 29820 17442 29876 17444
rect 29820 17390 29822 17442
rect 29822 17390 29874 17442
rect 29874 17390 29876 17442
rect 29820 17388 29876 17390
rect 29708 16828 29764 16884
rect 29708 16658 29764 16660
rect 29708 16606 29710 16658
rect 29710 16606 29762 16658
rect 29762 16606 29764 16658
rect 29708 16604 29764 16606
rect 30940 17052 30996 17108
rect 30492 16828 30548 16884
rect 29184 15706 29240 15708
rect 29184 15654 29186 15706
rect 29186 15654 29238 15706
rect 29238 15654 29240 15706
rect 29184 15652 29240 15654
rect 29288 15706 29344 15708
rect 29288 15654 29290 15706
rect 29290 15654 29342 15706
rect 29342 15654 29344 15706
rect 29288 15652 29344 15654
rect 29392 15706 29448 15708
rect 29392 15654 29394 15706
rect 29394 15654 29446 15706
rect 29446 15654 29448 15706
rect 29392 15652 29448 15654
rect 29036 15260 29092 15316
rect 29372 15148 29428 15204
rect 29036 14530 29092 14532
rect 29036 14478 29038 14530
rect 29038 14478 29090 14530
rect 29090 14478 29092 14530
rect 29036 14476 29092 14478
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 28588 13356 28644 13412
rect 29184 12570 29240 12572
rect 29184 12518 29186 12570
rect 29186 12518 29238 12570
rect 29238 12518 29240 12570
rect 29184 12516 29240 12518
rect 29288 12570 29344 12572
rect 29288 12518 29290 12570
rect 29290 12518 29342 12570
rect 29342 12518 29344 12570
rect 29288 12516 29344 12518
rect 29392 12570 29448 12572
rect 29392 12518 29394 12570
rect 29394 12518 29446 12570
rect 29446 12518 29448 12570
rect 29392 12516 29448 12518
rect 29036 12124 29092 12180
rect 30380 12738 30436 12740
rect 30380 12686 30382 12738
rect 30382 12686 30434 12738
rect 30434 12686 30436 12738
rect 30380 12684 30436 12686
rect 30156 12124 30212 12180
rect 30604 16044 30660 16100
rect 30828 16268 30884 16324
rect 31500 16268 31556 16324
rect 31276 16098 31332 16100
rect 31276 16046 31278 16098
rect 31278 16046 31330 16098
rect 31330 16046 31332 16098
rect 31276 16044 31332 16046
rect 30604 15148 30660 15204
rect 31500 14028 31556 14084
rect 31388 13468 31444 13524
rect 30716 13132 30772 13188
rect 30268 11676 30324 11732
rect 29708 11564 29764 11620
rect 29596 11116 29652 11172
rect 29184 11002 29240 11004
rect 29184 10950 29186 11002
rect 29186 10950 29238 11002
rect 29238 10950 29240 11002
rect 29184 10948 29240 10950
rect 29288 11002 29344 11004
rect 29288 10950 29290 11002
rect 29290 10950 29342 11002
rect 29342 10950 29344 11002
rect 29288 10948 29344 10950
rect 29392 11002 29448 11004
rect 29392 10950 29394 11002
rect 29394 10950 29446 11002
rect 29446 10950 29448 11002
rect 29392 10948 29448 10950
rect 28252 9660 28308 9716
rect 29596 9772 29652 9828
rect 29184 9434 29240 9436
rect 29184 9382 29186 9434
rect 29186 9382 29238 9434
rect 29238 9382 29240 9434
rect 29184 9380 29240 9382
rect 29288 9434 29344 9436
rect 29288 9382 29290 9434
rect 29290 9382 29342 9434
rect 29342 9382 29344 9434
rect 29288 9380 29344 9382
rect 29392 9434 29448 9436
rect 29392 9382 29394 9434
rect 29394 9382 29446 9434
rect 29446 9382 29448 9434
rect 29392 9380 29448 9382
rect 27580 8988 27636 9044
rect 28924 8930 28980 8932
rect 28924 8878 28926 8930
rect 28926 8878 28978 8930
rect 28978 8878 28980 8930
rect 28924 8876 28980 8878
rect 27916 8540 27972 8596
rect 27692 8428 27748 8484
rect 27356 7420 27412 7476
rect 27244 6860 27300 6916
rect 26684 6636 26740 6692
rect 26572 5964 26628 6020
rect 24522 5514 24578 5516
rect 24522 5462 24524 5514
rect 24524 5462 24576 5514
rect 24576 5462 24578 5514
rect 24522 5460 24578 5462
rect 24626 5514 24682 5516
rect 24626 5462 24628 5514
rect 24628 5462 24680 5514
rect 24680 5462 24682 5514
rect 24626 5460 24682 5462
rect 24730 5514 24786 5516
rect 24730 5462 24732 5514
rect 24732 5462 24784 5514
rect 24784 5462 24786 5514
rect 24730 5460 24786 5462
rect 26460 5628 26516 5684
rect 26348 4844 26404 4900
rect 26124 4450 26180 4452
rect 26124 4398 26126 4450
rect 26126 4398 26178 4450
rect 26178 4398 26180 4450
rect 26124 4396 26180 4398
rect 27692 6690 27748 6692
rect 27692 6638 27694 6690
rect 27694 6638 27746 6690
rect 27746 6638 27748 6690
rect 27692 6636 27748 6638
rect 29184 7866 29240 7868
rect 29184 7814 29186 7866
rect 29186 7814 29238 7866
rect 29238 7814 29240 7866
rect 29184 7812 29240 7814
rect 29288 7866 29344 7868
rect 29288 7814 29290 7866
rect 29290 7814 29342 7866
rect 29342 7814 29344 7866
rect 29288 7812 29344 7814
rect 29392 7866 29448 7868
rect 29392 7814 29394 7866
rect 29394 7814 29446 7866
rect 29446 7814 29448 7866
rect 29392 7812 29448 7814
rect 29820 8258 29876 8260
rect 29820 8206 29822 8258
rect 29822 8206 29874 8258
rect 29874 8206 29876 8258
rect 29820 8204 29876 8206
rect 30044 8034 30100 8036
rect 30044 7982 30046 8034
rect 30046 7982 30098 8034
rect 30098 7982 30100 8034
rect 30044 7980 30100 7982
rect 28700 7362 28756 7364
rect 28700 7310 28702 7362
rect 28702 7310 28754 7362
rect 28754 7310 28756 7362
rect 28700 7308 28756 7310
rect 28588 6972 28644 7028
rect 27692 6130 27748 6132
rect 27692 6078 27694 6130
rect 27694 6078 27746 6130
rect 27746 6078 27748 6130
rect 27692 6076 27748 6078
rect 26908 5292 26964 5348
rect 26684 4562 26740 4564
rect 26684 4510 26686 4562
rect 26686 4510 26738 4562
rect 26738 4510 26740 4562
rect 26684 4508 26740 4510
rect 24522 3946 24578 3948
rect 24522 3894 24524 3946
rect 24524 3894 24576 3946
rect 24576 3894 24578 3946
rect 24522 3892 24578 3894
rect 24626 3946 24682 3948
rect 24626 3894 24628 3946
rect 24628 3894 24680 3946
rect 24680 3894 24682 3946
rect 24626 3892 24682 3894
rect 24730 3946 24786 3948
rect 24730 3894 24732 3946
rect 24732 3894 24784 3946
rect 24784 3894 24786 3946
rect 24730 3892 24786 3894
rect 27132 5404 27188 5460
rect 28028 6018 28084 6020
rect 28028 5966 28030 6018
rect 28030 5966 28082 6018
rect 28082 5966 28084 6018
rect 28028 5964 28084 5966
rect 27468 5628 27524 5684
rect 27692 5740 27748 5796
rect 27244 4620 27300 4676
rect 27132 4396 27188 4452
rect 27132 4060 27188 4116
rect 26124 3442 26180 3444
rect 26124 3390 26126 3442
rect 26126 3390 26178 3442
rect 26178 3390 26180 3442
rect 26124 3388 26180 3390
rect 27692 3724 27748 3780
rect 27580 3388 27636 3444
rect 28812 6748 28868 6804
rect 28364 6018 28420 6020
rect 28364 5966 28366 6018
rect 28366 5966 28418 6018
rect 28418 5966 28420 6018
rect 28364 5964 28420 5966
rect 29260 6636 29316 6692
rect 28252 4508 28308 4564
rect 28364 4620 28420 4676
rect 28028 3500 28084 3556
rect 28700 4844 28756 4900
rect 29184 6298 29240 6300
rect 29184 6246 29186 6298
rect 29186 6246 29238 6298
rect 29238 6246 29240 6298
rect 29184 6244 29240 6246
rect 29288 6298 29344 6300
rect 29288 6246 29290 6298
rect 29290 6246 29342 6298
rect 29342 6246 29344 6298
rect 29288 6244 29344 6246
rect 29392 6298 29448 6300
rect 29392 6246 29394 6298
rect 29394 6246 29446 6298
rect 29446 6246 29448 6298
rect 29392 6244 29448 6246
rect 29372 5292 29428 5348
rect 29596 5964 29652 6020
rect 29708 5906 29764 5908
rect 29708 5854 29710 5906
rect 29710 5854 29762 5906
rect 29762 5854 29764 5906
rect 29708 5852 29764 5854
rect 29260 4898 29316 4900
rect 29260 4846 29262 4898
rect 29262 4846 29314 4898
rect 29314 4846 29316 4898
rect 29260 4844 29316 4846
rect 29184 4730 29240 4732
rect 29184 4678 29186 4730
rect 29186 4678 29238 4730
rect 29238 4678 29240 4730
rect 29184 4676 29240 4678
rect 29288 4730 29344 4732
rect 29288 4678 29290 4730
rect 29290 4678 29342 4730
rect 29342 4678 29344 4730
rect 29288 4676 29344 4678
rect 29392 4730 29448 4732
rect 29392 4678 29394 4730
rect 29394 4678 29446 4730
rect 29446 4678 29448 4730
rect 29392 4676 29448 4678
rect 29036 4562 29092 4564
rect 29036 4510 29038 4562
rect 29038 4510 29090 4562
rect 29090 4510 29092 4562
rect 29036 4508 29092 4510
rect 29372 4338 29428 4340
rect 29372 4286 29374 4338
rect 29374 4286 29426 4338
rect 29426 4286 29428 4338
rect 29372 4284 29428 4286
rect 29036 4172 29092 4228
rect 30940 12124 30996 12180
rect 31052 11170 31108 11172
rect 31052 11118 31054 11170
rect 31054 11118 31106 11170
rect 31106 11118 31108 11170
rect 31052 11116 31108 11118
rect 31276 10556 31332 10612
rect 31164 9154 31220 9156
rect 31164 9102 31166 9154
rect 31166 9102 31218 9154
rect 31218 9102 31220 9154
rect 31164 9100 31220 9102
rect 30940 8764 30996 8820
rect 34188 24722 34244 24724
rect 34188 24670 34190 24722
rect 34190 24670 34242 24722
rect 34242 24670 34244 24722
rect 34188 24668 34244 24670
rect 33846 24330 33902 24332
rect 33846 24278 33848 24330
rect 33848 24278 33900 24330
rect 33900 24278 33902 24330
rect 33846 24276 33902 24278
rect 33950 24330 34006 24332
rect 33950 24278 33952 24330
rect 33952 24278 34004 24330
rect 34004 24278 34006 24330
rect 33950 24276 34006 24278
rect 34054 24330 34110 24332
rect 34054 24278 34056 24330
rect 34056 24278 34108 24330
rect 34108 24278 34110 24330
rect 34054 24276 34110 24278
rect 34188 23996 34244 24052
rect 33964 22876 34020 22932
rect 33846 22762 33902 22764
rect 33846 22710 33848 22762
rect 33848 22710 33900 22762
rect 33900 22710 33902 22762
rect 33846 22708 33902 22710
rect 33950 22762 34006 22764
rect 33950 22710 33952 22762
rect 33952 22710 34004 22762
rect 34004 22710 34006 22762
rect 33950 22708 34006 22710
rect 34054 22762 34110 22764
rect 34054 22710 34056 22762
rect 34056 22710 34108 22762
rect 34108 22710 34110 22762
rect 34054 22708 34110 22710
rect 33404 21420 33460 21476
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 33180 20748 33236 20804
rect 31948 19740 32004 19796
rect 33068 20636 33124 20692
rect 33292 20188 33348 20244
rect 31948 16994 32004 16996
rect 31948 16942 31950 16994
rect 31950 16942 32002 16994
rect 32002 16942 32004 16994
rect 31948 16940 32004 16942
rect 32956 19234 33012 19236
rect 32956 19182 32958 19234
rect 32958 19182 33010 19234
rect 33010 19182 33012 19234
rect 32956 19180 33012 19182
rect 32732 19010 32788 19012
rect 32732 18958 32734 19010
rect 32734 18958 32786 19010
rect 32786 18958 32788 19010
rect 32732 18956 32788 18958
rect 32172 16940 32228 16996
rect 33068 17388 33124 17444
rect 32732 16828 32788 16884
rect 33846 19626 33902 19628
rect 33846 19574 33848 19626
rect 33848 19574 33900 19626
rect 33900 19574 33902 19626
rect 33846 19572 33902 19574
rect 33950 19626 34006 19628
rect 33950 19574 33952 19626
rect 33952 19574 34004 19626
rect 34004 19574 34006 19626
rect 33950 19572 34006 19574
rect 34054 19626 34110 19628
rect 34054 19574 34056 19626
rect 34056 19574 34108 19626
rect 34108 19574 34110 19626
rect 34054 19572 34110 19574
rect 33516 19234 33572 19236
rect 33516 19182 33518 19234
rect 33518 19182 33570 19234
rect 33570 19182 33572 19234
rect 33516 19180 33572 19182
rect 35644 35756 35700 35812
rect 35196 35084 35252 35140
rect 35644 35138 35700 35140
rect 35644 35086 35646 35138
rect 35646 35086 35698 35138
rect 35698 35086 35700 35138
rect 35644 35084 35700 35086
rect 35196 34300 35252 34356
rect 34972 33628 35028 33684
rect 34748 28028 34804 28084
rect 34860 31052 34916 31108
rect 34636 27020 34692 27076
rect 34524 26236 34580 26292
rect 34524 23100 34580 23156
rect 34860 26460 34916 26516
rect 37548 39004 37604 39060
rect 36092 34188 36148 34244
rect 35420 33292 35476 33348
rect 35420 32284 35476 32340
rect 35084 30156 35140 30212
rect 35420 31388 35476 31444
rect 35420 28476 35476 28532
rect 35308 28364 35364 28420
rect 34972 25228 35028 25284
rect 35196 24722 35252 24724
rect 35196 24670 35198 24722
rect 35198 24670 35250 24722
rect 35250 24670 35252 24722
rect 35196 24668 35252 24670
rect 35420 24556 35476 24612
rect 34636 21532 34692 21588
rect 35980 25340 36036 25396
rect 36428 36316 36484 36372
rect 36652 35868 36708 35924
rect 36988 35868 37044 35924
rect 37100 35308 37156 35364
rect 36316 33180 36372 33236
rect 36204 31276 36260 31332
rect 37324 33404 37380 33460
rect 37100 33346 37156 33348
rect 37100 33294 37102 33346
rect 37102 33294 37154 33346
rect 37154 33294 37156 33346
rect 37100 33292 37156 33294
rect 36428 31388 36484 31444
rect 36316 29820 36372 29876
rect 36428 26290 36484 26292
rect 36428 26238 36430 26290
rect 36430 26238 36482 26290
rect 36482 26238 36484 26290
rect 36428 26236 36484 26238
rect 36876 32732 36932 32788
rect 36764 29650 36820 29652
rect 36764 29598 36766 29650
rect 36766 29598 36818 29650
rect 36818 29598 36820 29650
rect 36764 29596 36820 29598
rect 36876 27020 36932 27076
rect 37772 38332 37828 38388
rect 37660 36988 37716 37044
rect 37772 34972 37828 35028
rect 37884 34748 37940 34804
rect 38220 37660 38276 37716
rect 37772 33516 37828 33572
rect 37100 31612 37156 31668
rect 37212 31218 37268 31220
rect 37212 31166 37214 31218
rect 37214 31166 37266 31218
rect 37266 31166 37268 31218
rect 37212 31164 37268 31166
rect 37548 31554 37604 31556
rect 37548 31502 37550 31554
rect 37550 31502 37602 31554
rect 37602 31502 37604 31554
rect 37548 31500 37604 31502
rect 37660 30940 37716 30996
rect 37548 30268 37604 30324
rect 38508 36090 38564 36092
rect 38508 36038 38510 36090
rect 38510 36038 38562 36090
rect 38562 36038 38564 36090
rect 38508 36036 38564 36038
rect 38612 36090 38668 36092
rect 38612 36038 38614 36090
rect 38614 36038 38666 36090
rect 38666 36038 38668 36090
rect 38612 36036 38668 36038
rect 38716 36090 38772 36092
rect 38716 36038 38718 36090
rect 38718 36038 38770 36090
rect 38770 36038 38772 36090
rect 38716 36036 38772 36038
rect 38220 33458 38276 33460
rect 38220 33406 38222 33458
rect 38222 33406 38274 33458
rect 38274 33406 38276 33458
rect 38220 33404 38276 33406
rect 38332 35644 38388 35700
rect 37884 33180 37940 33236
rect 38508 34522 38564 34524
rect 38508 34470 38510 34522
rect 38510 34470 38562 34522
rect 38562 34470 38564 34522
rect 38508 34468 38564 34470
rect 38612 34522 38668 34524
rect 38612 34470 38614 34522
rect 38614 34470 38666 34522
rect 38666 34470 38668 34522
rect 38612 34468 38668 34470
rect 38716 34522 38772 34524
rect 38716 34470 38718 34522
rect 38718 34470 38770 34522
rect 38770 34470 38772 34522
rect 38716 34468 38772 34470
rect 38508 32954 38564 32956
rect 38508 32902 38510 32954
rect 38510 32902 38562 32954
rect 38562 32902 38564 32954
rect 38508 32900 38564 32902
rect 38612 32954 38668 32956
rect 38612 32902 38614 32954
rect 38614 32902 38666 32954
rect 38666 32902 38668 32954
rect 38612 32900 38668 32902
rect 38716 32954 38772 32956
rect 38716 32902 38718 32954
rect 38718 32902 38770 32954
rect 38770 32902 38772 32954
rect 38716 32900 38772 32902
rect 37884 31276 37940 31332
rect 38220 31500 38276 31556
rect 38508 31386 38564 31388
rect 38508 31334 38510 31386
rect 38510 31334 38562 31386
rect 38562 31334 38564 31386
rect 38508 31332 38564 31334
rect 38612 31386 38668 31388
rect 38612 31334 38614 31386
rect 38614 31334 38666 31386
rect 38666 31334 38668 31386
rect 38612 31332 38668 31334
rect 38716 31386 38772 31388
rect 38716 31334 38718 31386
rect 38718 31334 38770 31386
rect 38770 31334 38772 31386
rect 38716 31332 38772 31334
rect 37772 30156 37828 30212
rect 37884 29820 37940 29876
rect 38508 29818 38564 29820
rect 38508 29766 38510 29818
rect 38510 29766 38562 29818
rect 38562 29766 38564 29818
rect 38508 29764 38564 29766
rect 38612 29818 38668 29820
rect 38612 29766 38614 29818
rect 38614 29766 38666 29818
rect 38666 29766 38668 29818
rect 38612 29764 38668 29766
rect 38716 29818 38772 29820
rect 38716 29766 38718 29818
rect 38718 29766 38770 29818
rect 38770 29766 38772 29818
rect 38716 29764 38772 29766
rect 38220 29596 38276 29652
rect 37212 28924 37268 28980
rect 37660 28642 37716 28644
rect 37660 28590 37662 28642
rect 37662 28590 37714 28642
rect 37714 28590 37716 28642
rect 37660 28588 37716 28590
rect 38220 28924 38276 28980
rect 38108 28642 38164 28644
rect 38108 28590 38110 28642
rect 38110 28590 38162 28642
rect 38162 28590 38164 28642
rect 38108 28588 38164 28590
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 37884 28082 37940 28084
rect 37884 28030 37886 28082
rect 37886 28030 37938 28082
rect 37938 28030 37940 28082
rect 37884 28028 37940 28030
rect 37660 27580 37716 27636
rect 38220 27580 38276 27636
rect 36988 25394 37044 25396
rect 36988 25342 36990 25394
rect 36990 25342 37042 25394
rect 37042 25342 37044 25394
rect 36988 25340 37044 25342
rect 36204 24892 36260 24948
rect 36092 24668 36148 24724
rect 36988 24050 37044 24052
rect 36988 23998 36990 24050
rect 36990 23998 37042 24050
rect 37042 23998 37044 24050
rect 36988 23996 37044 23998
rect 38220 26796 38276 26852
rect 37884 26514 37940 26516
rect 37884 26462 37886 26514
rect 37886 26462 37938 26514
rect 37938 26462 37940 26514
rect 37884 26460 37940 26462
rect 37772 26236 37828 26292
rect 38508 26682 38564 26684
rect 38508 26630 38510 26682
rect 38510 26630 38562 26682
rect 38562 26630 38564 26682
rect 38508 26628 38564 26630
rect 38612 26682 38668 26684
rect 38612 26630 38614 26682
rect 38614 26630 38666 26682
rect 38666 26630 38668 26682
rect 38612 26628 38668 26630
rect 38716 26682 38772 26684
rect 38716 26630 38718 26682
rect 38718 26630 38770 26682
rect 38770 26630 38772 26682
rect 38716 26628 38772 26630
rect 37548 25564 37604 25620
rect 38508 25114 38564 25116
rect 38508 25062 38510 25114
rect 38510 25062 38562 25114
rect 38562 25062 38564 25114
rect 38508 25060 38564 25062
rect 38612 25114 38668 25116
rect 38612 25062 38614 25114
rect 38614 25062 38666 25114
rect 38666 25062 38668 25114
rect 38612 25060 38668 25062
rect 38716 25114 38772 25116
rect 38716 25062 38718 25114
rect 38718 25062 38770 25114
rect 38770 25062 38772 25114
rect 38716 25060 38772 25062
rect 38220 24946 38276 24948
rect 38220 24894 38222 24946
rect 38222 24894 38274 24946
rect 38274 24894 38276 24946
rect 38220 24892 38276 24894
rect 37212 23996 37268 24052
rect 36092 23378 36148 23380
rect 36092 23326 36094 23378
rect 36094 23326 36146 23378
rect 36146 23326 36148 23378
rect 36092 23324 36148 23326
rect 36988 23324 37044 23380
rect 38220 24556 38276 24612
rect 38508 23546 38564 23548
rect 38508 23494 38510 23546
rect 38510 23494 38562 23546
rect 38562 23494 38564 23546
rect 38508 23492 38564 23494
rect 38612 23546 38668 23548
rect 38612 23494 38614 23546
rect 38614 23494 38666 23546
rect 38666 23494 38668 23546
rect 38612 23492 38668 23494
rect 38716 23546 38772 23548
rect 38716 23494 38718 23546
rect 38718 23494 38770 23546
rect 38770 23494 38772 23546
rect 38716 23492 38772 23494
rect 38508 21978 38564 21980
rect 38508 21926 38510 21978
rect 38510 21926 38562 21978
rect 38562 21926 38564 21978
rect 38508 21924 38564 21926
rect 38612 21978 38668 21980
rect 38612 21926 38614 21978
rect 38614 21926 38666 21978
rect 38666 21926 38668 21978
rect 38612 21924 38668 21926
rect 38716 21978 38772 21980
rect 38716 21926 38718 21978
rect 38718 21926 38770 21978
rect 38770 21926 38772 21978
rect 38716 21924 38772 21926
rect 34972 20188 35028 20244
rect 38508 20410 38564 20412
rect 38508 20358 38510 20410
rect 38510 20358 38562 20410
rect 38562 20358 38564 20410
rect 38508 20356 38564 20358
rect 38612 20410 38668 20412
rect 38612 20358 38614 20410
rect 38614 20358 38666 20410
rect 38666 20358 38668 20410
rect 38612 20356 38668 20358
rect 38716 20410 38772 20412
rect 38716 20358 38718 20410
rect 38718 20358 38770 20410
rect 38770 20358 38772 20410
rect 38716 20356 38772 20358
rect 34860 20076 34916 20132
rect 34412 19964 34468 20020
rect 34300 18508 34356 18564
rect 35084 19180 35140 19236
rect 33846 18058 33902 18060
rect 33846 18006 33848 18058
rect 33848 18006 33900 18058
rect 33900 18006 33902 18058
rect 33846 18004 33902 18006
rect 33950 18058 34006 18060
rect 33950 18006 33952 18058
rect 33952 18006 34004 18058
rect 34004 18006 34006 18058
rect 33950 18004 34006 18006
rect 34054 18058 34110 18060
rect 34054 18006 34056 18058
rect 34056 18006 34108 18058
rect 34108 18006 34110 18058
rect 34054 18004 34110 18006
rect 33516 17052 33572 17108
rect 31612 13020 31668 13076
rect 31724 15260 31780 15316
rect 31836 13858 31892 13860
rect 31836 13806 31838 13858
rect 31838 13806 31890 13858
rect 31890 13806 31892 13858
rect 31836 13804 31892 13806
rect 33846 16490 33902 16492
rect 33846 16438 33848 16490
rect 33848 16438 33900 16490
rect 33900 16438 33902 16490
rect 33846 16436 33902 16438
rect 33950 16490 34006 16492
rect 33950 16438 33952 16490
rect 33952 16438 34004 16490
rect 34004 16438 34006 16490
rect 33950 16436 34006 16438
rect 34054 16490 34110 16492
rect 34054 16438 34056 16490
rect 34056 16438 34108 16490
rect 34108 16438 34110 16490
rect 34054 16436 34110 16438
rect 33740 15932 33796 15988
rect 32956 15202 33012 15204
rect 32956 15150 32958 15202
rect 32958 15150 33010 15202
rect 33010 15150 33012 15202
rect 32956 15148 33012 15150
rect 34972 17052 35028 17108
rect 34636 16940 34692 16996
rect 34300 16882 34356 16884
rect 34300 16830 34302 16882
rect 34302 16830 34354 16882
rect 34354 16830 34356 16882
rect 34300 16828 34356 16830
rect 34748 16882 34804 16884
rect 34748 16830 34750 16882
rect 34750 16830 34802 16882
rect 34802 16830 34804 16882
rect 34748 16828 34804 16830
rect 34636 15260 34692 15316
rect 32284 15090 32340 15092
rect 32284 15038 32286 15090
rect 32286 15038 32338 15090
rect 32338 15038 32340 15090
rect 32284 15036 32340 15038
rect 33292 15036 33348 15092
rect 32844 14530 32900 14532
rect 32844 14478 32846 14530
rect 32846 14478 32898 14530
rect 32898 14478 32900 14530
rect 32844 14476 32900 14478
rect 32172 14306 32228 14308
rect 32172 14254 32174 14306
rect 32174 14254 32226 14306
rect 32226 14254 32228 14306
rect 32172 14252 32228 14254
rect 32732 13916 32788 13972
rect 32620 13132 32676 13188
rect 31948 12796 32004 12852
rect 32396 11564 32452 11620
rect 31612 10108 31668 10164
rect 31500 9212 31556 9268
rect 30604 6972 30660 7028
rect 30492 6748 30548 6804
rect 30380 5292 30436 5348
rect 30156 4956 30212 5012
rect 30492 4844 30548 4900
rect 30604 4620 30660 4676
rect 29708 3724 29764 3780
rect 29596 3612 29652 3668
rect 29184 3162 29240 3164
rect 29184 3110 29186 3162
rect 29186 3110 29238 3162
rect 29238 3110 29240 3162
rect 29184 3108 29240 3110
rect 29288 3162 29344 3164
rect 29288 3110 29290 3162
rect 29290 3110 29342 3162
rect 29342 3110 29344 3162
rect 29288 3108 29344 3110
rect 29392 3162 29448 3164
rect 29392 3110 29394 3162
rect 29394 3110 29446 3162
rect 29446 3110 29448 3162
rect 29392 3108 29448 3110
rect 30492 3666 30548 3668
rect 30492 3614 30494 3666
rect 30494 3614 30546 3666
rect 30546 3614 30548 3666
rect 30492 3612 30548 3614
rect 31500 6972 31556 7028
rect 31948 9714 32004 9716
rect 31948 9662 31950 9714
rect 31950 9662 32002 9714
rect 32002 9662 32004 9714
rect 31948 9660 32004 9662
rect 31836 7196 31892 7252
rect 32172 6972 32228 7028
rect 31948 5852 32004 5908
rect 31948 5180 32004 5236
rect 32508 10668 32564 10724
rect 32396 8540 32452 8596
rect 33068 14252 33124 14308
rect 32956 13692 33012 13748
rect 33846 14922 33902 14924
rect 33846 14870 33848 14922
rect 33848 14870 33900 14922
rect 33900 14870 33902 14922
rect 33846 14868 33902 14870
rect 33950 14922 34006 14924
rect 33950 14870 33952 14922
rect 33952 14870 34004 14922
rect 34004 14870 34006 14922
rect 33950 14868 34006 14870
rect 34054 14922 34110 14924
rect 34054 14870 34056 14922
rect 34056 14870 34108 14922
rect 34108 14870 34110 14922
rect 34054 14868 34110 14870
rect 33404 13916 33460 13972
rect 33740 13858 33796 13860
rect 33740 13806 33742 13858
rect 33742 13806 33794 13858
rect 33794 13806 33796 13858
rect 33740 13804 33796 13806
rect 33292 13580 33348 13636
rect 33628 13580 33684 13636
rect 33292 12684 33348 12740
rect 33964 13580 34020 13636
rect 33846 13354 33902 13356
rect 33846 13302 33848 13354
rect 33848 13302 33900 13354
rect 33900 13302 33902 13354
rect 33846 13300 33902 13302
rect 33950 13354 34006 13356
rect 33950 13302 33952 13354
rect 33952 13302 34004 13354
rect 34004 13302 34006 13354
rect 33950 13300 34006 13302
rect 34054 13354 34110 13356
rect 34054 13302 34056 13354
rect 34056 13302 34108 13354
rect 34108 13302 34110 13354
rect 34054 13300 34110 13302
rect 32956 9212 33012 9268
rect 32732 8876 32788 8932
rect 32060 5068 32116 5124
rect 30940 4338 30996 4340
rect 30940 4286 30942 4338
rect 30942 4286 30994 4338
rect 30994 4286 30996 4338
rect 30940 4284 30996 4286
rect 31612 4172 31668 4228
rect 30940 3724 30996 3780
rect 32284 4732 32340 4788
rect 32172 3554 32228 3556
rect 32172 3502 32174 3554
rect 32174 3502 32226 3554
rect 32226 3502 32228 3554
rect 32172 3500 32228 3502
rect 32956 8540 33012 8596
rect 32844 7308 32900 7364
rect 32956 6076 33012 6132
rect 33068 7196 33124 7252
rect 33846 11786 33902 11788
rect 33846 11734 33848 11786
rect 33848 11734 33900 11786
rect 33900 11734 33902 11786
rect 33846 11732 33902 11734
rect 33950 11786 34006 11788
rect 33950 11734 33952 11786
rect 33952 11734 34004 11786
rect 34004 11734 34006 11786
rect 33950 11732 34006 11734
rect 34054 11786 34110 11788
rect 34054 11734 34056 11786
rect 34056 11734 34108 11786
rect 34108 11734 34110 11786
rect 34054 11732 34110 11734
rect 34636 13746 34692 13748
rect 34636 13694 34638 13746
rect 34638 13694 34690 13746
rect 34690 13694 34692 13746
rect 34636 13692 34692 13694
rect 34636 13468 34692 13524
rect 34524 13074 34580 13076
rect 34524 13022 34526 13074
rect 34526 13022 34578 13074
rect 34578 13022 34580 13074
rect 34524 13020 34580 13022
rect 34188 11228 34244 11284
rect 34300 11116 34356 11172
rect 33628 10610 33684 10612
rect 33628 10558 33630 10610
rect 33630 10558 33682 10610
rect 33682 10558 33684 10610
rect 33628 10556 33684 10558
rect 33292 10108 33348 10164
rect 33846 10218 33902 10220
rect 33846 10166 33848 10218
rect 33848 10166 33900 10218
rect 33900 10166 33902 10218
rect 33846 10164 33902 10166
rect 33950 10218 34006 10220
rect 33950 10166 33952 10218
rect 33952 10166 34004 10218
rect 34004 10166 34006 10218
rect 33950 10164 34006 10166
rect 34054 10218 34110 10220
rect 34054 10166 34056 10218
rect 34056 10166 34108 10218
rect 34108 10166 34110 10218
rect 34054 10164 34110 10166
rect 34076 9996 34132 10052
rect 33852 9938 33908 9940
rect 33852 9886 33854 9938
rect 33854 9886 33906 9938
rect 33906 9886 33908 9938
rect 33852 9884 33908 9886
rect 33404 9548 33460 9604
rect 33628 9154 33684 9156
rect 33628 9102 33630 9154
rect 33630 9102 33682 9154
rect 33682 9102 33684 9154
rect 33628 9100 33684 9102
rect 34524 11564 34580 11620
rect 34524 11282 34580 11284
rect 34524 11230 34526 11282
rect 34526 11230 34578 11282
rect 34578 11230 34580 11282
rect 34524 11228 34580 11230
rect 33846 8650 33902 8652
rect 33628 8540 33684 8596
rect 33846 8598 33848 8650
rect 33848 8598 33900 8650
rect 33900 8598 33902 8650
rect 33846 8596 33902 8598
rect 33950 8650 34006 8652
rect 33950 8598 33952 8650
rect 33952 8598 34004 8650
rect 34004 8598 34006 8650
rect 33950 8596 34006 8598
rect 34054 8650 34110 8652
rect 34054 8598 34056 8650
rect 34056 8598 34108 8650
rect 34108 8598 34110 8650
rect 34054 8596 34110 8598
rect 33292 6860 33348 6916
rect 33404 6412 33460 6468
rect 33180 5404 33236 5460
rect 33068 3442 33124 3444
rect 33068 3390 33070 3442
rect 33070 3390 33122 3442
rect 33122 3390 33124 3442
rect 33068 3388 33124 3390
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 34076 6860 34132 6916
rect 34748 9884 34804 9940
rect 34748 9714 34804 9716
rect 34748 9662 34750 9714
rect 34750 9662 34802 9714
rect 34802 9662 34804 9714
rect 34748 9660 34804 9662
rect 34972 9436 35028 9492
rect 34748 9042 34804 9044
rect 34748 8990 34750 9042
rect 34750 8990 34802 9042
rect 34802 8990 34804 9042
rect 34748 8988 34804 8990
rect 33852 5740 33908 5796
rect 33846 5514 33902 5516
rect 33846 5462 33848 5514
rect 33848 5462 33900 5514
rect 33900 5462 33902 5514
rect 33846 5460 33902 5462
rect 33950 5514 34006 5516
rect 33950 5462 33952 5514
rect 33952 5462 34004 5514
rect 34004 5462 34006 5514
rect 33950 5460 34006 5462
rect 34054 5514 34110 5516
rect 34054 5462 34056 5514
rect 34056 5462 34108 5514
rect 34108 5462 34110 5514
rect 34054 5460 34110 5462
rect 33516 4226 33572 4228
rect 33516 4174 33518 4226
rect 33518 4174 33570 4226
rect 33570 4174 33572 4226
rect 33516 4172 33572 4174
rect 34188 4172 34244 4228
rect 33846 3946 33902 3948
rect 33846 3894 33848 3946
rect 33848 3894 33900 3946
rect 33900 3894 33902 3946
rect 33846 3892 33902 3894
rect 33950 3946 34006 3948
rect 33950 3894 33952 3946
rect 33952 3894 34004 3946
rect 34004 3894 34006 3946
rect 33950 3892 34006 3894
rect 34054 3946 34110 3948
rect 34054 3894 34056 3946
rect 34056 3894 34108 3946
rect 34108 3894 34110 3946
rect 34054 3892 34110 3894
rect 37436 20076 37492 20132
rect 36092 18396 36148 18452
rect 35980 18284 36036 18340
rect 35868 18172 35924 18228
rect 35196 13468 35252 13524
rect 35532 12850 35588 12852
rect 35532 12798 35534 12850
rect 35534 12798 35586 12850
rect 35586 12798 35588 12850
rect 35532 12796 35588 12798
rect 35196 11170 35252 11172
rect 35196 11118 35198 11170
rect 35198 11118 35250 11170
rect 35250 11118 35252 11170
rect 35196 11116 35252 11118
rect 35420 10444 35476 10500
rect 35532 8876 35588 8932
rect 36764 18508 36820 18564
rect 36652 18226 36708 18228
rect 36652 18174 36654 18226
rect 36654 18174 36706 18226
rect 36706 18174 36708 18226
rect 36652 18172 36708 18174
rect 35980 15148 36036 15204
rect 35980 13132 36036 13188
rect 35980 12684 36036 12740
rect 35756 11116 35812 11172
rect 36204 16828 36260 16884
rect 35756 9826 35812 9828
rect 35756 9774 35758 9826
rect 35758 9774 35810 9826
rect 35810 9774 35812 9826
rect 35756 9772 35812 9774
rect 35980 10220 36036 10276
rect 36428 15314 36484 15316
rect 36428 15262 36430 15314
rect 36430 15262 36482 15314
rect 36482 15262 36484 15314
rect 36428 15260 36484 15262
rect 36540 14028 36596 14084
rect 36428 10780 36484 10836
rect 36876 18450 36932 18452
rect 36876 18398 36878 18450
rect 36878 18398 36930 18450
rect 36930 18398 36932 18450
rect 36876 18396 36932 18398
rect 36988 15986 37044 15988
rect 36988 15934 36990 15986
rect 36990 15934 37042 15986
rect 37042 15934 37044 15986
rect 36988 15932 37044 15934
rect 36652 10386 36708 10388
rect 36652 10334 36654 10386
rect 36654 10334 36706 10386
rect 36706 10334 36708 10386
rect 36652 10332 36708 10334
rect 36540 10220 36596 10276
rect 35196 7868 35252 7924
rect 35084 7532 35140 7588
rect 34972 7362 35028 7364
rect 34972 7310 34974 7362
rect 34974 7310 35026 7362
rect 35026 7310 35028 7362
rect 34972 7308 35028 7310
rect 34748 6860 34804 6916
rect 33964 1036 34020 1092
rect 34524 5180 34580 5236
rect 34636 4060 34692 4116
rect 34972 6578 35028 6580
rect 34972 6526 34974 6578
rect 34974 6526 35026 6578
rect 35026 6526 35028 6578
rect 34972 6524 35028 6526
rect 34748 3388 34804 3444
rect 34972 3612 35028 3668
rect 35868 5964 35924 6020
rect 35644 5068 35700 5124
rect 35196 3724 35252 3780
rect 35084 2716 35140 2772
rect 36092 8316 36148 8372
rect 35980 4620 36036 4676
rect 36316 8204 36372 8260
rect 36652 7586 36708 7588
rect 36652 7534 36654 7586
rect 36654 7534 36706 7586
rect 36706 7534 36708 7586
rect 36652 7532 36708 7534
rect 36428 6860 36484 6916
rect 36316 5628 36372 5684
rect 36988 11394 37044 11396
rect 36988 11342 36990 11394
rect 36990 11342 37042 11394
rect 37042 11342 37044 11394
rect 36988 11340 37044 11342
rect 36988 10108 37044 10164
rect 36988 9602 37044 9604
rect 36988 9550 36990 9602
rect 36990 9550 37042 9602
rect 37042 9550 37044 9602
rect 36988 9548 37044 9550
rect 37884 18338 37940 18340
rect 37884 18286 37886 18338
rect 37886 18286 37938 18338
rect 37938 18286 37940 18338
rect 37884 18284 37940 18286
rect 37548 16828 37604 16884
rect 37212 13580 37268 13636
rect 37884 13132 37940 13188
rect 37212 12738 37268 12740
rect 37212 12686 37214 12738
rect 37214 12686 37266 12738
rect 37266 12686 37268 12738
rect 37212 12684 37268 12686
rect 37324 12572 37380 12628
rect 37772 12738 37828 12740
rect 37772 12686 37774 12738
rect 37774 12686 37826 12738
rect 37826 12686 37828 12738
rect 37772 12684 37828 12686
rect 37548 10668 37604 10724
rect 37100 8316 37156 8372
rect 36988 8034 37044 8036
rect 36988 7982 36990 8034
rect 36990 7982 37042 8034
rect 37042 7982 37044 8034
rect 36988 7980 37044 7982
rect 36988 7474 37044 7476
rect 36988 7422 36990 7474
rect 36990 7422 37042 7474
rect 37042 7422 37044 7474
rect 36988 7420 37044 7422
rect 36988 6466 37044 6468
rect 36988 6414 36990 6466
rect 36990 6414 37042 6466
rect 37042 6414 37044 6466
rect 36988 6412 37044 6414
rect 37772 10050 37828 10052
rect 37772 9998 37774 10050
rect 37774 9998 37826 10050
rect 37826 9998 37828 10050
rect 37772 9996 37828 9998
rect 37772 9212 37828 9268
rect 37884 8428 37940 8484
rect 37772 7420 37828 7476
rect 37548 6076 37604 6132
rect 37660 6636 37716 6692
rect 37436 5628 37492 5684
rect 36204 4620 36260 4676
rect 36988 5292 37044 5348
rect 36876 4508 36932 4564
rect 36428 3666 36484 3668
rect 36428 3614 36430 3666
rect 36430 3614 36482 3666
rect 36482 3614 36484 3666
rect 36428 3612 36484 3614
rect 37324 3276 37380 3332
rect 37548 4956 37604 5012
rect 38508 18842 38564 18844
rect 38508 18790 38510 18842
rect 38510 18790 38562 18842
rect 38562 18790 38564 18842
rect 38508 18788 38564 18790
rect 38612 18842 38668 18844
rect 38612 18790 38614 18842
rect 38614 18790 38666 18842
rect 38666 18790 38668 18842
rect 38612 18788 38668 18790
rect 38716 18842 38772 18844
rect 38716 18790 38718 18842
rect 38718 18790 38770 18842
rect 38770 18790 38772 18842
rect 38716 18788 38772 18790
rect 38108 16268 38164 16324
rect 38508 17274 38564 17276
rect 38508 17222 38510 17274
rect 38510 17222 38562 17274
rect 38562 17222 38564 17274
rect 38508 17220 38564 17222
rect 38612 17274 38668 17276
rect 38612 17222 38614 17274
rect 38614 17222 38666 17274
rect 38666 17222 38668 17274
rect 38612 17220 38668 17222
rect 38716 17274 38772 17276
rect 38716 17222 38718 17274
rect 38718 17222 38770 17274
rect 38770 17222 38772 17274
rect 38716 17220 38772 17222
rect 38892 16156 38948 16212
rect 38508 15706 38564 15708
rect 38508 15654 38510 15706
rect 38510 15654 38562 15706
rect 38562 15654 38564 15706
rect 38508 15652 38564 15654
rect 38612 15706 38668 15708
rect 38612 15654 38614 15706
rect 38614 15654 38666 15706
rect 38666 15654 38668 15706
rect 38612 15652 38668 15654
rect 38716 15706 38772 15708
rect 38716 15654 38718 15706
rect 38718 15654 38770 15706
rect 38770 15654 38772 15706
rect 38716 15652 38772 15654
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 38508 12570 38564 12572
rect 38508 12518 38510 12570
rect 38510 12518 38562 12570
rect 38562 12518 38564 12570
rect 38508 12516 38564 12518
rect 38612 12570 38668 12572
rect 38612 12518 38614 12570
rect 38614 12518 38666 12570
rect 38666 12518 38668 12570
rect 38612 12516 38668 12518
rect 38716 12570 38772 12572
rect 38716 12518 38718 12570
rect 38718 12518 38770 12570
rect 38770 12518 38772 12570
rect 38716 12516 38772 12518
rect 38108 11506 38164 11508
rect 38108 11454 38110 11506
rect 38110 11454 38162 11506
rect 38162 11454 38164 11506
rect 38108 11452 38164 11454
rect 38508 11002 38564 11004
rect 38508 10950 38510 11002
rect 38510 10950 38562 11002
rect 38562 10950 38564 11002
rect 38508 10948 38564 10950
rect 38612 11002 38668 11004
rect 38612 10950 38614 11002
rect 38614 10950 38666 11002
rect 38666 10950 38668 11002
rect 38612 10948 38668 10950
rect 38716 11002 38772 11004
rect 38716 10950 38718 11002
rect 38718 10950 38770 11002
rect 38770 10950 38772 11002
rect 38716 10948 38772 10950
rect 38332 10834 38388 10836
rect 38332 10782 38334 10834
rect 38334 10782 38386 10834
rect 38386 10782 38388 10834
rect 38332 10780 38388 10782
rect 38508 9434 38564 9436
rect 38508 9382 38510 9434
rect 38510 9382 38562 9434
rect 38562 9382 38564 9434
rect 38508 9380 38564 9382
rect 38612 9434 38668 9436
rect 38612 9382 38614 9434
rect 38614 9382 38666 9434
rect 38666 9382 38668 9434
rect 38612 9380 38668 9382
rect 38716 9434 38772 9436
rect 38716 9382 38718 9434
rect 38718 9382 38770 9434
rect 38770 9382 38772 9434
rect 38716 9380 38772 9382
rect 38108 8092 38164 8148
rect 38508 7866 38564 7868
rect 38508 7814 38510 7866
rect 38510 7814 38562 7866
rect 38562 7814 38564 7866
rect 38508 7812 38564 7814
rect 38612 7866 38668 7868
rect 38612 7814 38614 7866
rect 38614 7814 38666 7866
rect 38666 7814 38668 7866
rect 38612 7812 38668 7814
rect 38716 7866 38772 7868
rect 38716 7814 38718 7866
rect 38718 7814 38770 7866
rect 38770 7814 38772 7866
rect 38716 7812 38772 7814
rect 38508 6298 38564 6300
rect 38508 6246 38510 6298
rect 38510 6246 38562 6298
rect 38562 6246 38564 6298
rect 38508 6244 38564 6246
rect 38612 6298 38668 6300
rect 38612 6246 38614 6298
rect 38614 6246 38666 6298
rect 38666 6246 38668 6298
rect 38612 6244 38668 6246
rect 38716 6298 38772 6300
rect 38716 6246 38718 6298
rect 38718 6246 38770 6298
rect 38770 6246 38772 6298
rect 38716 6244 38772 6246
rect 38508 4730 38564 4732
rect 37772 4620 37828 4676
rect 38508 4678 38510 4730
rect 38510 4678 38562 4730
rect 38562 4678 38564 4730
rect 38508 4676 38564 4678
rect 38612 4730 38668 4732
rect 38612 4678 38614 4730
rect 38614 4678 38666 4730
rect 38666 4678 38668 4730
rect 38612 4676 38668 4678
rect 38716 4730 38772 4732
rect 38716 4678 38718 4730
rect 38718 4678 38770 4730
rect 38770 4678 38772 4730
rect 38716 4676 38772 4678
rect 38108 4284 38164 4340
rect 37884 3276 37940 3332
rect 37884 1372 37940 1428
rect 38508 3162 38564 3164
rect 38508 3110 38510 3162
rect 38510 3110 38562 3162
rect 38562 3110 38564 3162
rect 38508 3108 38564 3110
rect 38612 3162 38668 3164
rect 38612 3110 38614 3162
rect 38614 3110 38666 3162
rect 38666 3110 38668 3162
rect 38612 3108 38668 3110
rect 38716 3162 38772 3164
rect 38716 3110 38718 3162
rect 38718 3110 38770 3162
rect 38770 3110 38772 3162
rect 38716 3108 38772 3110
rect 39676 3724 39732 3780
rect 37436 28 37492 84
<< metal3 >>
rect 39200 39732 40000 39760
rect 35186 39676 35196 39732
rect 35252 39676 40000 39732
rect 39200 39648 40000 39676
rect 39200 39060 40000 39088
rect 37538 39004 37548 39060
rect 37604 39004 40000 39060
rect 39200 38976 40000 39004
rect 39200 38388 40000 38416
rect 37762 38332 37772 38388
rect 37828 38332 40000 38388
rect 39200 38304 40000 38332
rect 39200 37716 40000 37744
rect 38210 37660 38220 37716
rect 38276 37660 40000 37716
rect 39200 37632 40000 37660
rect 39200 37044 40000 37072
rect 37650 36988 37660 37044
rect 37716 36988 40000 37044
rect 39200 36960 40000 36988
rect 21522 36876 21532 36932
rect 21588 36876 22540 36932
rect 22596 36876 22606 36932
rect 32946 36876 32956 36932
rect 33012 36876 33628 36932
rect 33684 36876 33694 36932
rect 5864 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6148 36876
rect 15188 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15472 36876
rect 24512 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24796 36876
rect 33836 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34120 36876
rect 24882 36652 24892 36708
rect 24948 36652 26124 36708
rect 26180 36652 26190 36708
rect 27570 36652 27580 36708
rect 27636 36652 28812 36708
rect 28868 36652 28878 36708
rect 30930 36652 30940 36708
rect 30996 36652 32620 36708
rect 32676 36652 32686 36708
rect 32274 36540 32284 36596
rect 32340 36540 34412 36596
rect 34468 36540 34478 36596
rect 29698 36428 29708 36484
rect 29764 36428 30268 36484
rect 30324 36428 30716 36484
rect 30772 36428 30782 36484
rect 39200 36372 40000 36400
rect 27122 36316 27132 36372
rect 27188 36316 28924 36372
rect 28980 36316 28990 36372
rect 34178 36316 34188 36372
rect 34244 36316 35308 36372
rect 35364 36316 35374 36372
rect 36418 36316 36428 36372
rect 36484 36316 40000 36372
rect 39200 36288 40000 36316
rect 17938 36204 17948 36260
rect 18004 36204 20748 36260
rect 20804 36204 20814 36260
rect 21522 36204 21532 36260
rect 21588 36204 22652 36260
rect 22708 36204 22718 36260
rect 30706 36204 30716 36260
rect 30772 36204 32172 36260
rect 32228 36204 32238 36260
rect 10526 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10810 36092
rect 19850 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20134 36092
rect 29174 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29458 36092
rect 38498 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38782 36092
rect 20178 35868 20188 35924
rect 20244 35868 21084 35924
rect 21140 35868 21150 35924
rect 31938 35868 31948 35924
rect 32004 35868 33740 35924
rect 33796 35868 33806 35924
rect 36642 35868 36652 35924
rect 36708 35868 36988 35924
rect 37044 35868 37054 35924
rect 18610 35756 18620 35812
rect 18676 35756 21868 35812
rect 21924 35756 21934 35812
rect 24098 35756 24108 35812
rect 24164 35756 26124 35812
rect 26180 35756 26190 35812
rect 32386 35756 32396 35812
rect 32452 35756 34748 35812
rect 34804 35756 34814 35812
rect 35074 35756 35084 35812
rect 35140 35756 35644 35812
rect 35700 35756 35710 35812
rect 35084 35700 35140 35756
rect 39200 35700 40000 35728
rect 34514 35644 34524 35700
rect 34580 35644 35140 35700
rect 38322 35644 38332 35700
rect 38388 35644 40000 35700
rect 39200 35616 40000 35644
rect 34738 35308 34748 35364
rect 34804 35308 37100 35364
rect 37156 35308 37166 35364
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 35186 35084 35196 35140
rect 35252 35084 35644 35140
rect 35700 35084 35710 35140
rect 39200 35028 40000 35056
rect 37762 34972 37772 35028
rect 37828 34972 40000 35028
rect 39200 34944 40000 34972
rect 23426 34860 23436 34916
rect 23492 34860 25340 34916
rect 25396 34860 25406 34916
rect 24770 34748 24780 34804
rect 24836 34748 26684 34804
rect 26740 34748 26750 34804
rect 33506 34748 33516 34804
rect 33572 34748 37884 34804
rect 37940 34748 37950 34804
rect 10526 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10810 34524
rect 19850 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20134 34524
rect 29174 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29458 34524
rect 38498 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38782 34524
rect 39200 34356 40000 34384
rect 35186 34300 35196 34356
rect 35252 34300 40000 34356
rect 39200 34272 40000 34300
rect 34066 34188 34076 34244
rect 34132 34188 36092 34244
rect 36148 34188 36158 34244
rect 5864 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6148 33740
rect 15188 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15472 33740
rect 24512 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24796 33740
rect 33836 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34120 33740
rect 39200 33684 40000 33712
rect 34962 33628 34972 33684
rect 35028 33628 40000 33684
rect 39200 33600 40000 33628
rect 34514 33516 34524 33572
rect 34580 33516 37772 33572
rect 37828 33516 37838 33572
rect 37314 33404 37324 33460
rect 37380 33404 38220 33460
rect 38276 33404 38286 33460
rect 35410 33292 35420 33348
rect 35476 33292 37100 33348
rect 37156 33292 37166 33348
rect 32610 33180 32620 33236
rect 32676 33180 34076 33236
rect 34132 33180 34142 33236
rect 36306 33180 36316 33236
rect 36372 33180 37884 33236
rect 37940 33180 37950 33236
rect 39200 33012 40000 33040
rect 38892 32956 40000 33012
rect 10526 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10810 32956
rect 19850 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20134 32956
rect 29174 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29458 32956
rect 38498 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38782 32956
rect 38892 32788 38948 32956
rect 39200 32928 40000 32956
rect 36866 32732 36876 32788
rect 36932 32732 38948 32788
rect 39200 32340 40000 32368
rect 35410 32284 35420 32340
rect 35476 32284 40000 32340
rect 39200 32256 40000 32284
rect 5864 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6148 32172
rect 15188 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15472 32172
rect 24512 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24796 32172
rect 33836 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34120 32172
rect 39200 31668 40000 31696
rect 37090 31612 37100 31668
rect 37156 31612 40000 31668
rect 39200 31584 40000 31612
rect 37538 31500 37548 31556
rect 37604 31500 38220 31556
rect 38276 31500 38286 31556
rect 35410 31388 35420 31444
rect 35476 31388 36428 31444
rect 36484 31388 36494 31444
rect 10526 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10810 31388
rect 19850 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20134 31388
rect 29174 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29458 31388
rect 38498 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38782 31388
rect 36194 31276 36204 31332
rect 36260 31276 37884 31332
rect 37940 31276 37950 31332
rect 31602 31164 31612 31220
rect 31668 31164 37212 31220
rect 37268 31164 37278 31220
rect 34402 31052 34412 31108
rect 34468 31052 34860 31108
rect 34916 31052 34926 31108
rect 39200 30996 40000 31024
rect 37650 30940 37660 30996
rect 37716 30940 40000 30996
rect 39200 30912 40000 30940
rect 5864 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6148 30604
rect 15188 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15472 30604
rect 24512 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24796 30604
rect 33836 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34120 30604
rect 39200 30324 40000 30352
rect 37538 30268 37548 30324
rect 37604 30268 40000 30324
rect 39200 30240 40000 30268
rect 35074 30156 35084 30212
rect 35140 30156 37772 30212
rect 37828 30156 37838 30212
rect 9426 29932 9436 29988
rect 9492 29932 10444 29988
rect 10500 29932 10510 29988
rect 36306 29820 36316 29876
rect 36372 29820 37884 29876
rect 37940 29820 37950 29876
rect 10526 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10810 29820
rect 19850 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20134 29820
rect 29174 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29458 29820
rect 38498 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38782 29820
rect 39200 29652 40000 29680
rect 36754 29596 36764 29652
rect 36820 29596 38220 29652
rect 38276 29596 40000 29652
rect 39200 29568 40000 29596
rect 12450 29484 12460 29540
rect 12516 29484 13356 29540
rect 13412 29484 13422 29540
rect 33506 29372 33516 29428
rect 33572 29372 34300 29428
rect 34356 29372 34366 29428
rect 12226 29036 12236 29092
rect 12292 29036 14476 29092
rect 14532 29036 14542 29092
rect 5864 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6148 29036
rect 15188 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15472 29036
rect 24512 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24796 29036
rect 33836 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34120 29036
rect 39200 28980 40000 29008
rect 37202 28924 37212 28980
rect 37268 28924 38220 28980
rect 38276 28924 40000 28980
rect 39200 28896 40000 28924
rect 29922 28812 29932 28868
rect 29988 28812 32060 28868
rect 32116 28812 32126 28868
rect 8642 28700 8652 28756
rect 8708 28700 9660 28756
rect 9716 28700 9726 28756
rect 12114 28700 12124 28756
rect 12180 28700 15260 28756
rect 15316 28700 15326 28756
rect 15698 28700 15708 28756
rect 15764 28700 18060 28756
rect 18116 28700 18126 28756
rect 27122 28700 27132 28756
rect 27188 28700 30156 28756
rect 30212 28700 30222 28756
rect 37650 28588 37660 28644
rect 37716 28588 38108 28644
rect 38164 28588 38948 28644
rect 13010 28476 13020 28532
rect 13076 28476 15036 28532
rect 15092 28476 15102 28532
rect 16034 28476 16044 28532
rect 16100 28476 19068 28532
rect 19124 28476 19134 28532
rect 26002 28476 26012 28532
rect 26068 28476 28028 28532
rect 28084 28476 28094 28532
rect 28802 28476 28812 28532
rect 28868 28476 31164 28532
rect 31220 28476 31230 28532
rect 33170 28476 33180 28532
rect 33236 28476 35420 28532
rect 35476 28476 35486 28532
rect 32722 28364 32732 28420
rect 32788 28364 35308 28420
rect 35364 28364 35374 28420
rect 38892 28308 38948 28588
rect 39200 28308 40000 28336
rect 29586 28252 29596 28308
rect 29652 28252 31052 28308
rect 31108 28252 31118 28308
rect 38892 28252 40000 28308
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 39200 28224 40000 28252
rect 33394 28140 33404 28196
rect 33460 28140 34412 28196
rect 34468 28140 34478 28196
rect 15362 28028 15372 28084
rect 15428 28028 16268 28084
rect 16324 28028 16334 28084
rect 34738 28028 34748 28084
rect 34804 28028 37884 28084
rect 37940 28028 37950 28084
rect 5506 27916 5516 27972
rect 5572 27916 7980 27972
rect 8036 27916 8046 27972
rect 18274 27916 18284 27972
rect 18340 27916 19628 27972
rect 19684 27916 19694 27972
rect 21074 27916 21084 27972
rect 21140 27916 22316 27972
rect 22372 27916 22382 27972
rect 11778 27804 11788 27860
rect 11844 27804 12572 27860
rect 12628 27804 12638 27860
rect 8306 27692 8316 27748
rect 8372 27692 10668 27748
rect 10724 27692 10734 27748
rect 13234 27692 13244 27748
rect 13300 27692 15820 27748
rect 15876 27692 15886 27748
rect 24210 27692 24220 27748
rect 24276 27692 28476 27748
rect 28532 27692 28542 27748
rect 39200 27636 40000 27664
rect 37650 27580 37660 27636
rect 37716 27580 38220 27636
rect 38276 27580 40000 27636
rect 39200 27552 40000 27580
rect 25778 27468 25788 27524
rect 25844 27468 27020 27524
rect 27076 27468 27086 27524
rect 5864 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6148 27468
rect 15188 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15472 27468
rect 24512 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24796 27468
rect 33836 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34120 27468
rect 9986 27356 9996 27412
rect 10052 27356 12348 27412
rect 12404 27356 12414 27412
rect 12562 27020 12572 27076
rect 12628 27020 14588 27076
rect 14644 27020 14654 27076
rect 29698 27020 29708 27076
rect 29764 27020 32956 27076
rect 33012 27020 33022 27076
rect 34626 27020 34636 27076
rect 34692 27020 36876 27076
rect 36932 27020 36942 27076
rect 39200 26964 40000 26992
rect 6066 26908 6076 26964
rect 6132 26908 6972 26964
rect 7028 26908 7038 26964
rect 9100 26908 11452 26964
rect 11508 26908 11518 26964
rect 11666 26908 11676 26964
rect 11732 26908 13468 26964
rect 13524 26908 13534 26964
rect 27570 26908 27580 26964
rect 27636 26908 29148 26964
rect 29204 26908 29214 26964
rect 38220 26908 40000 26964
rect 9100 26852 9156 26908
rect 38220 26852 38276 26908
rect 39200 26880 40000 26908
rect 9090 26796 9100 26852
rect 9156 26796 9166 26852
rect 31154 26796 31164 26852
rect 31220 26796 33180 26852
rect 33236 26796 33246 26852
rect 38210 26796 38220 26852
rect 38276 26796 38286 26852
rect 30146 26684 30156 26740
rect 30212 26684 34188 26740
rect 34244 26684 34254 26740
rect 10526 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10810 26684
rect 19850 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20134 26684
rect 29174 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29458 26684
rect 38498 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38782 26684
rect 8418 26460 8428 26516
rect 8484 26460 10892 26516
rect 10948 26460 10958 26516
rect 14690 26460 14700 26516
rect 14756 26460 16380 26516
rect 16436 26460 16446 26516
rect 16594 26460 16604 26516
rect 16660 26460 18508 26516
rect 18564 26460 18574 26516
rect 34850 26460 34860 26516
rect 34916 26460 37884 26516
rect 37940 26460 37950 26516
rect 14130 26348 14140 26404
rect 14196 26348 15260 26404
rect 15316 26348 15326 26404
rect 0 26292 800 26320
rect 39200 26292 40000 26320
rect 0 26236 4284 26292
rect 4340 26236 4350 26292
rect 5282 26236 5292 26292
rect 5348 26236 5628 26292
rect 5684 26236 5694 26292
rect 24658 26236 24668 26292
rect 24724 26236 25340 26292
rect 25396 26236 25406 26292
rect 33058 26236 33068 26292
rect 33124 26236 34076 26292
rect 34132 26236 34524 26292
rect 34580 26236 36428 26292
rect 36484 26236 36494 26292
rect 37762 26236 37772 26292
rect 37828 26236 40000 26292
rect 0 26208 800 26236
rect 39200 26208 40000 26236
rect 13682 26124 13692 26180
rect 13748 26124 16268 26180
rect 16324 26124 16334 26180
rect 17826 26124 17836 26180
rect 17892 26124 19404 26180
rect 19460 26124 19470 26180
rect 5864 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6148 25900
rect 15188 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15472 25900
rect 24512 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24796 25900
rect 33836 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34120 25900
rect 16706 25788 16716 25844
rect 16772 25788 18620 25844
rect 18676 25788 18686 25844
rect 39200 25620 40000 25648
rect 3490 25564 3500 25620
rect 3556 25564 4620 25620
rect 4676 25564 4686 25620
rect 21634 25564 21644 25620
rect 21700 25564 22428 25620
rect 22484 25564 22494 25620
rect 23986 25564 23996 25620
rect 24052 25564 25564 25620
rect 25620 25564 25630 25620
rect 37538 25564 37548 25620
rect 37604 25564 40000 25620
rect 39200 25536 40000 25564
rect 8082 25452 8092 25508
rect 8148 25452 9548 25508
rect 9604 25452 9614 25508
rect 29250 25452 29260 25508
rect 29316 25452 33068 25508
rect 33124 25452 33134 25508
rect 1474 25340 1484 25396
rect 1540 25340 2156 25396
rect 2212 25340 2222 25396
rect 6290 25340 6300 25396
rect 6356 25340 10108 25396
rect 10164 25340 10174 25396
rect 20850 25340 20860 25396
rect 20916 25340 23548 25396
rect 23604 25340 23614 25396
rect 35970 25340 35980 25396
rect 36036 25340 36988 25396
rect 37044 25340 37054 25396
rect 5170 25228 5180 25284
rect 5236 25228 5628 25284
rect 5684 25228 8988 25284
rect 9044 25228 9054 25284
rect 18834 25228 18844 25284
rect 18900 25228 20300 25284
rect 20356 25228 21532 25284
rect 21588 25228 21598 25284
rect 33842 25228 33852 25284
rect 33908 25228 34972 25284
rect 35028 25228 35038 25284
rect 11106 25116 11116 25172
rect 11172 25116 11900 25172
rect 11956 25116 11966 25172
rect 10526 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10810 25116
rect 19850 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20134 25116
rect 29174 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29458 25116
rect 38498 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38782 25116
rect 10994 25004 11004 25060
rect 11060 25004 13692 25060
rect 13748 25004 13758 25060
rect 21858 24892 21868 24948
rect 21924 24892 25228 24948
rect 25284 24892 25294 24948
rect 29586 24892 29596 24948
rect 29652 24892 30492 24948
rect 30548 24892 30558 24948
rect 36194 24892 36204 24948
rect 36260 24892 38220 24948
rect 38276 24892 38286 24948
rect 1586 24780 1596 24836
rect 1652 24780 2268 24836
rect 2324 24780 2334 24836
rect 19282 24780 19292 24836
rect 19348 24780 21308 24836
rect 21364 24780 21374 24836
rect 4050 24668 4060 24724
rect 4116 24668 5292 24724
rect 5348 24668 5358 24724
rect 10322 24668 10332 24724
rect 10388 24668 11004 24724
rect 11060 24668 11070 24724
rect 11442 24668 11452 24724
rect 11508 24668 12572 24724
rect 12628 24668 12638 24724
rect 22194 24668 22204 24724
rect 22260 24668 23436 24724
rect 23492 24668 25340 24724
rect 25396 24668 26684 24724
rect 26740 24668 26750 24724
rect 31938 24668 31948 24724
rect 32004 24668 33404 24724
rect 33460 24668 34188 24724
rect 34244 24668 34254 24724
rect 35186 24668 35196 24724
rect 35252 24668 36092 24724
rect 36148 24668 36158 24724
rect 35410 24556 35420 24612
rect 35476 24556 38220 24612
rect 38276 24556 38286 24612
rect 5864 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6148 24332
rect 15188 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15472 24332
rect 24512 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24796 24332
rect 33836 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34120 24332
rect 24770 24108 24780 24164
rect 24836 24108 26572 24164
rect 26628 24108 26638 24164
rect 12450 23996 12460 24052
rect 12516 23996 13468 24052
rect 13524 23996 13534 24052
rect 27122 23996 27132 24052
rect 27188 23996 32956 24052
rect 33012 23996 33022 24052
rect 34178 23996 34188 24052
rect 34244 23996 36988 24052
rect 37044 23996 37212 24052
rect 37268 23996 37278 24052
rect 25554 23884 25564 23940
rect 25620 23884 26236 23940
rect 26292 23884 27580 23940
rect 27636 23884 28252 23940
rect 28308 23884 30380 23940
rect 30436 23884 30446 23940
rect 1922 23772 1932 23828
rect 1988 23772 5740 23828
rect 5796 23772 6300 23828
rect 6356 23772 6366 23828
rect 6626 23772 6636 23828
rect 6692 23772 11452 23828
rect 11508 23772 11518 23828
rect 26450 23772 26460 23828
rect 26516 23772 27244 23828
rect 27300 23772 27310 23828
rect 3714 23660 3724 23716
rect 3780 23660 5852 23716
rect 5908 23660 5918 23716
rect 27010 23660 27020 23716
rect 27076 23660 31164 23716
rect 31220 23660 31230 23716
rect 10526 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10810 23548
rect 19850 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20134 23548
rect 29174 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29458 23548
rect 38498 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38782 23548
rect 3490 23436 3500 23492
rect 3556 23436 5964 23492
rect 6020 23436 6030 23492
rect 7074 23436 7084 23492
rect 7140 23436 7150 23492
rect 12674 23436 12684 23492
rect 12740 23436 16044 23492
rect 16100 23436 16716 23492
rect 16772 23436 17164 23492
rect 17220 23436 17230 23492
rect 7084 23380 7140 23436
rect 4722 23324 4732 23380
rect 4788 23324 7140 23380
rect 24210 23324 24220 23380
rect 24276 23324 28364 23380
rect 28420 23324 28430 23380
rect 36082 23324 36092 23380
rect 36148 23324 36988 23380
rect 37044 23324 37054 23380
rect 19506 23212 19516 23268
rect 19572 23212 20412 23268
rect 20468 23212 20478 23268
rect 4946 23100 4956 23156
rect 5012 23100 6412 23156
rect 6468 23100 6478 23156
rect 14690 23100 14700 23156
rect 14756 23100 15372 23156
rect 15428 23100 15438 23156
rect 21298 23100 21308 23156
rect 21364 23100 21868 23156
rect 21924 23100 21934 23156
rect 33170 23100 33180 23156
rect 33236 23100 34524 23156
rect 34580 23100 34590 23156
rect 10322 22988 10332 23044
rect 10388 22988 12572 23044
rect 12628 22988 12638 23044
rect 14018 22988 14028 23044
rect 14084 22988 17388 23044
rect 17444 22988 17454 23044
rect 28802 22876 28812 22932
rect 28868 22876 33964 22932
rect 34020 22876 34030 22932
rect 25778 22764 25788 22820
rect 25844 22764 30156 22820
rect 30212 22764 30222 22820
rect 5864 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6148 22764
rect 15188 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15472 22764
rect 24512 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24796 22764
rect 33836 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34120 22764
rect 7634 22540 7644 22596
rect 7700 22540 12404 22596
rect 4050 22428 4060 22484
rect 4116 22428 8428 22484
rect 8484 22428 8494 22484
rect 12348 22372 12404 22540
rect 22194 22428 22204 22484
rect 22260 22428 26460 22484
rect 26516 22428 26526 22484
rect 9202 22316 9212 22372
rect 9268 22316 10332 22372
rect 10388 22316 10398 22372
rect 12338 22316 12348 22372
rect 12404 22316 12414 22372
rect 19282 22316 19292 22372
rect 19348 22316 21756 22372
rect 21812 22316 21822 22372
rect 28578 22316 28588 22372
rect 28644 22316 29484 22372
rect 29540 22316 29550 22372
rect 22754 22204 22764 22260
rect 22820 22204 27468 22260
rect 27524 22204 27534 22260
rect 29250 22204 29260 22260
rect 29316 22204 29820 22260
rect 29876 22204 30828 22260
rect 30884 22204 30894 22260
rect 9874 22092 9884 22148
rect 9940 22092 14588 22148
rect 14644 22092 14654 22148
rect 15474 22092 15484 22148
rect 15540 22092 19740 22148
rect 19796 22092 23772 22148
rect 23828 22092 25564 22148
rect 25620 22092 29372 22148
rect 29428 22092 31164 22148
rect 31220 22092 31230 22148
rect 10526 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10810 21980
rect 19850 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20134 21980
rect 29174 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29458 21980
rect 38498 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38782 21980
rect 8530 21756 8540 21812
rect 8596 21756 9660 21812
rect 9716 21756 9726 21812
rect 12674 21756 12684 21812
rect 12740 21756 13692 21812
rect 13748 21756 13758 21812
rect 3042 21644 3052 21700
rect 3108 21644 9100 21700
rect 9156 21644 9166 21700
rect 17826 21644 17836 21700
rect 17892 21644 18508 21700
rect 18564 21644 18574 21700
rect 32050 21644 32060 21700
rect 32116 21644 33068 21700
rect 33124 21644 33134 21700
rect 18508 21588 18564 21644
rect 4162 21532 4172 21588
rect 4228 21532 5404 21588
rect 5460 21532 7756 21588
rect 7812 21532 7822 21588
rect 18508 21532 20636 21588
rect 20692 21532 21308 21588
rect 21364 21532 21812 21588
rect 25330 21532 25340 21588
rect 25396 21532 26908 21588
rect 26964 21532 26974 21588
rect 29586 21532 29596 21588
rect 29652 21532 34636 21588
rect 34692 21532 34702 21588
rect 21756 21476 21812 21532
rect 3938 21420 3948 21476
rect 4004 21420 6076 21476
rect 6132 21420 6142 21476
rect 9986 21420 9996 21476
rect 10052 21420 11564 21476
rect 11620 21420 11630 21476
rect 21746 21420 21756 21476
rect 21812 21420 21822 21476
rect 24658 21420 24668 21476
rect 24724 21420 27580 21476
rect 27636 21420 28476 21476
rect 28532 21420 28542 21476
rect 31714 21420 31724 21476
rect 31780 21420 33404 21476
rect 33460 21420 33470 21476
rect 4050 21308 4060 21364
rect 4116 21308 5964 21364
rect 6020 21308 6030 21364
rect 17938 21196 17948 21252
rect 18004 21196 19404 21252
rect 19460 21196 19470 21252
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 10098 21084 10108 21140
rect 10164 21084 12460 21140
rect 12516 21084 12526 21140
rect 4274 20972 4284 21028
rect 4340 20972 15036 21028
rect 15092 20972 15102 21028
rect 3042 20860 3052 20916
rect 3108 20860 13244 20916
rect 13300 20860 13310 20916
rect 13906 20860 13916 20916
rect 13972 20860 14812 20916
rect 14868 20860 14878 20916
rect 5954 20748 5964 20804
rect 6020 20748 6972 20804
rect 7028 20748 8092 20804
rect 8148 20748 9548 20804
rect 9604 20748 9614 20804
rect 12002 20748 12012 20804
rect 12068 20748 16380 20804
rect 16436 20748 16446 20804
rect 28914 20748 28924 20804
rect 28980 20748 31052 20804
rect 31108 20748 33180 20804
rect 33236 20748 33246 20804
rect 26786 20636 26796 20692
rect 26852 20636 28252 20692
rect 28308 20636 28318 20692
rect 28578 20636 28588 20692
rect 28644 20636 30380 20692
rect 30436 20636 33068 20692
rect 33124 20636 33134 20692
rect 11890 20524 11900 20580
rect 11956 20524 12796 20580
rect 12852 20524 13580 20580
rect 13636 20524 16716 20580
rect 16772 20524 22316 20580
rect 22372 20524 22988 20580
rect 23044 20524 23054 20580
rect 24210 20524 24220 20580
rect 24276 20524 27356 20580
rect 27412 20524 27422 20580
rect 10526 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10810 20412
rect 19850 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20134 20412
rect 29174 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29458 20412
rect 38498 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38782 20412
rect 7522 20188 7532 20244
rect 7588 20188 8764 20244
rect 8820 20188 11564 20244
rect 11620 20188 11630 20244
rect 16370 20188 16380 20244
rect 16436 20188 17612 20244
rect 17668 20188 17678 20244
rect 21522 20188 21532 20244
rect 21588 20188 23268 20244
rect 33282 20188 33292 20244
rect 33348 20188 34972 20244
rect 35028 20188 35038 20244
rect 3602 19964 3612 20020
rect 3668 19964 5964 20020
rect 6020 19964 6030 20020
rect 16146 19964 16156 20020
rect 16212 19964 17276 20020
rect 17332 19964 17342 20020
rect 23212 19908 23268 20188
rect 23426 20132 23436 20188
rect 23492 20132 23502 20188
rect 23436 20076 24220 20132
rect 24276 20076 24286 20132
rect 29810 20076 29820 20132
rect 29876 20076 30604 20132
rect 30660 20076 30670 20132
rect 34850 20076 34860 20132
rect 34916 20076 37436 20132
rect 37492 20076 37502 20132
rect 29138 19964 29148 20020
rect 29204 19964 34412 20020
rect 34468 19964 34478 20020
rect 15026 19852 15036 19908
rect 15092 19852 22092 19908
rect 22148 19852 22158 19908
rect 23202 19852 23212 19908
rect 23268 19852 23278 19908
rect 26898 19852 26908 19908
rect 26964 19852 30940 19908
rect 30996 19852 31006 19908
rect 3042 19740 3052 19796
rect 3108 19740 7756 19796
rect 7812 19740 7822 19796
rect 26002 19740 26012 19796
rect 26068 19740 31948 19796
rect 32004 19740 32014 19796
rect 5864 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6148 19628
rect 15188 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15472 19628
rect 24512 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24796 19628
rect 33836 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34120 19628
rect 10994 19404 11004 19460
rect 11060 19404 13356 19460
rect 13412 19404 13422 19460
rect 28588 19292 29820 19348
rect 29876 19292 30380 19348
rect 30436 19292 30446 19348
rect 28588 19236 28644 19292
rect 22978 19180 22988 19236
rect 23044 19180 27916 19236
rect 27972 19180 28588 19236
rect 28644 19180 28654 19236
rect 29250 19180 29260 19236
rect 29316 19180 32956 19236
rect 33012 19180 33022 19236
rect 33506 19180 33516 19236
rect 33572 19180 35084 19236
rect 35140 19180 35150 19236
rect 11442 19068 11452 19124
rect 11508 19068 12348 19124
rect 12404 19068 12414 19124
rect 2370 18956 2380 19012
rect 2436 18956 5852 19012
rect 5908 18956 5918 19012
rect 11106 18956 11116 19012
rect 11172 18956 11788 19012
rect 11844 18956 11854 19012
rect 14130 18956 14140 19012
rect 14196 18956 17388 19012
rect 17444 18956 17454 19012
rect 26562 18956 26572 19012
rect 26628 18956 27356 19012
rect 27412 18956 27422 19012
rect 27692 18956 32732 19012
rect 32788 18956 32798 19012
rect 27692 18900 27748 18956
rect 26450 18844 26460 18900
rect 26516 18844 27748 18900
rect 10526 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10810 18844
rect 19850 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20134 18844
rect 29174 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29458 18844
rect 38498 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38782 18844
rect 3714 18620 3724 18676
rect 3780 18620 13804 18676
rect 13860 18620 13870 18676
rect 10322 18508 10332 18564
rect 10388 18508 11004 18564
rect 11060 18508 11070 18564
rect 34290 18508 34300 18564
rect 34356 18508 36764 18564
rect 36820 18508 36830 18564
rect 3938 18396 3948 18452
rect 4004 18396 5852 18452
rect 5908 18396 5918 18452
rect 7746 18396 7756 18452
rect 7812 18396 10164 18452
rect 17042 18396 17052 18452
rect 17108 18396 18956 18452
rect 19012 18396 19022 18452
rect 36082 18396 36092 18452
rect 36148 18396 36876 18452
rect 36932 18396 36942 18452
rect 10108 18340 10164 18396
rect 3042 18284 3052 18340
rect 3108 18284 8988 18340
rect 9044 18284 9054 18340
rect 10098 18284 10108 18340
rect 10164 18284 10174 18340
rect 16818 18284 16828 18340
rect 16884 18284 17612 18340
rect 17668 18284 18060 18340
rect 18116 18284 20636 18340
rect 20692 18284 20702 18340
rect 23202 18284 23212 18340
rect 23268 18284 23884 18340
rect 23940 18284 23950 18340
rect 35970 18284 35980 18340
rect 36036 18284 37884 18340
rect 37940 18284 37950 18340
rect 4050 18172 4060 18228
rect 4116 18172 8652 18228
rect 8708 18172 8718 18228
rect 28242 18172 28252 18228
rect 28308 18172 29932 18228
rect 29988 18172 29998 18228
rect 35858 18172 35868 18228
rect 35924 18172 36652 18228
rect 36708 18172 36718 18228
rect 5864 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6148 18060
rect 15188 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15472 18060
rect 24512 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24796 18060
rect 33836 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34120 18060
rect 14802 17836 14812 17892
rect 14868 17836 16940 17892
rect 16996 17836 17006 17892
rect 17938 17836 17948 17892
rect 18004 17836 22876 17892
rect 22932 17836 22942 17892
rect 7970 17612 7980 17668
rect 8036 17612 13916 17668
rect 13972 17612 13982 17668
rect 19394 17612 19404 17668
rect 19460 17612 20188 17668
rect 20244 17612 20254 17668
rect 3042 17500 3052 17556
rect 3108 17500 5516 17556
rect 5572 17500 5582 17556
rect 6962 17388 6972 17444
rect 7028 17388 11788 17444
rect 11844 17388 11854 17444
rect 29810 17388 29820 17444
rect 29876 17388 33068 17444
rect 33124 17388 33134 17444
rect 10526 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10810 17276
rect 19850 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20134 17276
rect 29174 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29458 17276
rect 38498 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38782 17276
rect 21970 17164 21980 17220
rect 22036 17164 23884 17220
rect 23940 17164 24668 17220
rect 24724 17164 25564 17220
rect 25620 17164 27580 17220
rect 27636 17164 27646 17220
rect 12114 17052 12124 17108
rect 12180 17052 14028 17108
rect 14084 17052 14094 17108
rect 15474 17052 15484 17108
rect 15540 17052 16716 17108
rect 16772 17052 16782 17108
rect 22866 17052 22876 17108
rect 22932 17052 30940 17108
rect 30996 17052 31006 17108
rect 33506 17052 33516 17108
rect 33572 17052 34972 17108
rect 35028 17052 35038 17108
rect 2594 16940 2604 16996
rect 2660 16940 3500 16996
rect 3556 16940 3566 16996
rect 10770 16940 10780 16996
rect 10836 16940 11564 16996
rect 11620 16940 11630 16996
rect 24098 16940 24108 16996
rect 24164 16940 31948 16996
rect 32004 16940 32014 16996
rect 32162 16940 32172 16996
rect 32228 16940 34636 16996
rect 34692 16940 34702 16996
rect 39200 16884 40000 16912
rect 2146 16828 2156 16884
rect 2212 16828 5068 16884
rect 5124 16828 5134 16884
rect 5954 16828 5964 16884
rect 6020 16828 9996 16884
rect 10052 16828 10062 16884
rect 11330 16828 11340 16884
rect 11396 16828 13580 16884
rect 13636 16828 13646 16884
rect 20626 16828 20636 16884
rect 20692 16828 21532 16884
rect 21588 16828 22204 16884
rect 22260 16828 22270 16884
rect 26002 16828 26012 16884
rect 26068 16828 26348 16884
rect 26404 16828 26684 16884
rect 26740 16828 26750 16884
rect 29698 16828 29708 16884
rect 29764 16828 30492 16884
rect 30548 16828 30558 16884
rect 32722 16828 32732 16884
rect 32788 16828 34300 16884
rect 34356 16828 34366 16884
rect 34738 16828 34748 16884
rect 34804 16828 36204 16884
rect 36260 16828 36270 16884
rect 37538 16828 37548 16884
rect 37604 16828 40000 16884
rect 39200 16800 40000 16828
rect 3042 16716 3052 16772
rect 3108 16716 6860 16772
rect 6916 16716 6926 16772
rect 7522 16716 7532 16772
rect 7588 16716 10332 16772
rect 10388 16716 12124 16772
rect 12180 16716 12190 16772
rect 12898 16716 12908 16772
rect 12964 16716 23436 16772
rect 23492 16716 23502 16772
rect 2930 16604 2940 16660
rect 2996 16604 5628 16660
rect 5684 16604 5694 16660
rect 29670 16604 29708 16660
rect 29764 16604 29774 16660
rect 5864 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6148 16492
rect 15188 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15472 16492
rect 24512 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24796 16492
rect 33836 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34120 16492
rect 30818 16268 30828 16324
rect 30884 16268 31500 16324
rect 31556 16268 38108 16324
rect 38164 16268 38174 16324
rect 39200 16212 40000 16240
rect 8082 16156 8092 16212
rect 8148 16156 9884 16212
rect 9940 16156 9950 16212
rect 18946 16156 18956 16212
rect 19012 16156 21644 16212
rect 21700 16156 21710 16212
rect 38882 16156 38892 16212
rect 38948 16156 40000 16212
rect 39200 16128 40000 16156
rect 4050 16044 4060 16100
rect 4116 16044 8316 16100
rect 8372 16044 8382 16100
rect 13570 16044 13580 16100
rect 13636 16044 14140 16100
rect 14196 16044 16380 16100
rect 16436 16044 16446 16100
rect 21074 16044 21084 16100
rect 21140 16044 23100 16100
rect 23156 16044 23166 16100
rect 30594 16044 30604 16100
rect 30660 16044 31276 16100
rect 31332 16044 31342 16100
rect 4722 15932 4732 15988
rect 4788 15932 5628 15988
rect 5684 15932 5694 15988
rect 19282 15932 19292 15988
rect 19348 15932 20076 15988
rect 20132 15932 20142 15988
rect 33730 15932 33740 15988
rect 33796 15932 36988 15988
rect 37044 15932 37054 15988
rect 5058 15820 5068 15876
rect 5124 15820 5292 15876
rect 5348 15820 6412 15876
rect 6468 15820 7756 15876
rect 7812 15820 8540 15876
rect 8596 15820 8606 15876
rect 24210 15820 24220 15876
rect 24276 15820 27692 15876
rect 27748 15820 27758 15876
rect 8372 15428 8428 15820
rect 10526 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10810 15708
rect 19850 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20134 15708
rect 29174 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29458 15708
rect 38498 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38782 15708
rect 22754 15484 22764 15540
rect 22820 15484 23660 15540
rect 23716 15484 23726 15540
rect 39200 15456 40000 15568
rect 8372 15372 9100 15428
rect 9156 15372 12796 15428
rect 12852 15372 13580 15428
rect 13636 15372 13646 15428
rect 22642 15372 22652 15428
rect 22708 15372 24108 15428
rect 24164 15372 24174 15428
rect 7074 15260 7084 15316
rect 7140 15260 11452 15316
rect 11508 15260 11518 15316
rect 12114 15260 12124 15316
rect 12180 15260 15708 15316
rect 15764 15260 15774 15316
rect 16034 15260 16044 15316
rect 16100 15260 17836 15316
rect 17892 15260 20412 15316
rect 20468 15260 20478 15316
rect 29026 15260 29036 15316
rect 29092 15260 31724 15316
rect 31780 15260 31790 15316
rect 34626 15260 34636 15316
rect 34692 15260 36428 15316
rect 36484 15260 36494 15316
rect 15372 15204 15428 15260
rect 10098 15148 10108 15204
rect 10164 15148 15148 15204
rect 15204 15148 15214 15204
rect 15362 15148 15372 15204
rect 15428 15148 15438 15204
rect 16370 15148 16380 15204
rect 16436 15148 17500 15204
rect 17556 15148 17566 15204
rect 19506 15148 19516 15204
rect 19572 15148 23772 15204
rect 23828 15148 29372 15204
rect 29428 15148 30604 15204
rect 30660 15148 30670 15204
rect 32918 15148 32956 15204
rect 33012 15148 33022 15204
rect 33506 15148 33516 15204
rect 33572 15148 35980 15204
rect 36036 15148 36046 15204
rect 32274 15036 32284 15092
rect 32340 15036 33292 15092
rect 33348 15036 33358 15092
rect 0 14868 800 14896
rect 5864 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6148 14924
rect 15188 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15472 14924
rect 24512 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24796 14924
rect 33836 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34120 14924
rect 0 14812 1708 14868
rect 1764 14812 1774 14868
rect 17154 14812 17164 14868
rect 17220 14812 17230 14868
rect 0 14784 800 14812
rect 17164 14756 17220 14812
rect 39200 14784 40000 14896
rect 4946 14700 4956 14756
rect 5012 14700 17220 14756
rect 2258 14588 2268 14644
rect 2324 14588 3612 14644
rect 3668 14588 3678 14644
rect 16818 14588 16828 14644
rect 16884 14588 17276 14644
rect 17332 14588 19292 14644
rect 19348 14588 19964 14644
rect 20020 14588 20030 14644
rect 13010 14476 13020 14532
rect 13076 14476 13804 14532
rect 13860 14476 14812 14532
rect 14868 14476 19516 14532
rect 19572 14476 19582 14532
rect 29026 14476 29036 14532
rect 29092 14476 32844 14532
rect 32900 14476 32910 14532
rect 20738 14252 20748 14308
rect 20804 14252 23660 14308
rect 23716 14252 23726 14308
rect 32162 14252 32172 14308
rect 32228 14252 33068 14308
rect 33124 14252 33134 14308
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 39200 14112 40000 14224
rect 26562 14028 26572 14084
rect 26628 14028 27356 14084
rect 27412 14028 27422 14084
rect 31490 14028 31500 14084
rect 31556 14028 36540 14084
rect 36596 14028 36606 14084
rect 21298 13916 21308 13972
rect 21364 13916 22316 13972
rect 22372 13916 22382 13972
rect 32722 13916 32732 13972
rect 32788 13916 33404 13972
rect 33460 13916 33470 13972
rect 31826 13804 31836 13860
rect 31892 13804 33740 13860
rect 33796 13804 33806 13860
rect 32946 13692 32956 13748
rect 33012 13692 34636 13748
rect 34692 13692 34702 13748
rect 33282 13580 33292 13636
rect 33348 13580 33628 13636
rect 33684 13580 33964 13636
rect 34020 13580 37212 13636
rect 37268 13580 37278 13636
rect 1922 13468 1932 13524
rect 1988 13468 5740 13524
rect 5796 13468 5806 13524
rect 23202 13468 23212 13524
rect 23268 13468 25228 13524
rect 25284 13468 25788 13524
rect 25844 13468 25854 13524
rect 26674 13468 26684 13524
rect 26740 13468 31388 13524
rect 31444 13468 31454 13524
rect 34626 13468 34636 13524
rect 34692 13468 35196 13524
rect 35252 13468 35262 13524
rect 39200 13440 40000 13552
rect 26114 13356 26124 13412
rect 26180 13356 28588 13412
rect 28644 13356 28654 13412
rect 5864 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6148 13356
rect 15188 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15472 13356
rect 24512 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24796 13356
rect 33836 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34120 13356
rect 2034 13244 2044 13300
rect 2100 13244 4508 13300
rect 4564 13244 4574 13300
rect 20402 13244 20412 13300
rect 20468 13244 23324 13300
rect 23380 13244 23390 13300
rect 20962 13132 20972 13188
rect 21028 13132 22876 13188
rect 22932 13132 22942 13188
rect 30706 13132 30716 13188
rect 30772 13132 32620 13188
rect 32676 13132 32686 13188
rect 35970 13132 35980 13188
rect 36036 13132 37884 13188
rect 37940 13132 37950 13188
rect 17938 13020 17948 13076
rect 18004 13020 18620 13076
rect 18676 13020 18686 13076
rect 20132 13020 22204 13076
rect 22260 13020 22270 13076
rect 31602 13020 31612 13076
rect 31668 13020 34524 13076
rect 34580 13020 34590 13076
rect 17042 12908 17052 12964
rect 17108 12908 18284 12964
rect 18340 12908 18350 12964
rect 20132 12852 20188 13020
rect 21074 12908 21084 12964
rect 21140 12908 23212 12964
rect 23268 12908 23278 12964
rect 5954 12796 5964 12852
rect 6020 12796 6860 12852
rect 6916 12796 6926 12852
rect 17938 12796 17948 12852
rect 18004 12796 20188 12852
rect 21522 12796 21532 12852
rect 21588 12796 22428 12852
rect 22484 12796 23324 12852
rect 23380 12796 23390 12852
rect 31938 12796 31948 12852
rect 32004 12796 35532 12852
rect 35588 12796 35598 12852
rect 39200 12768 40000 12880
rect 9762 12684 9772 12740
rect 9828 12684 10556 12740
rect 10612 12684 10622 12740
rect 30370 12684 30380 12740
rect 30436 12684 33292 12740
rect 33348 12684 33358 12740
rect 35970 12684 35980 12740
rect 36036 12684 37212 12740
rect 37268 12684 37278 12740
rect 37762 12684 37772 12740
rect 37828 12684 37838 12740
rect 37772 12628 37828 12684
rect 21746 12572 21756 12628
rect 21812 12572 25116 12628
rect 25172 12572 25182 12628
rect 37314 12572 37324 12628
rect 37380 12572 37828 12628
rect 10526 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10810 12572
rect 19850 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20134 12572
rect 29174 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29458 12572
rect 38498 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38782 12572
rect 9538 12460 9548 12516
rect 9604 12460 10332 12516
rect 10388 12460 10398 12516
rect 12450 12348 12460 12404
rect 12516 12348 13916 12404
rect 13972 12348 13982 12404
rect 8306 12236 8316 12292
rect 8372 12236 10108 12292
rect 10164 12236 10174 12292
rect 16370 12236 16380 12292
rect 16436 12236 17724 12292
rect 17780 12236 17790 12292
rect 20132 12236 21532 12292
rect 21588 12236 21598 12292
rect 24546 12236 24556 12292
rect 24612 12236 25564 12292
rect 25620 12236 27580 12292
rect 27636 12236 27646 12292
rect 5618 12124 5628 12180
rect 5684 12124 7308 12180
rect 7364 12124 8092 12180
rect 8148 12124 8158 12180
rect 16930 12124 16940 12180
rect 16996 12124 18844 12180
rect 18900 12124 18910 12180
rect 20132 12068 20188 12236
rect 25778 12124 25788 12180
rect 25844 12124 29036 12180
rect 29092 12124 29102 12180
rect 30146 12124 30156 12180
rect 30212 12124 30940 12180
rect 30996 12124 31006 12180
rect 39200 12096 40000 12208
rect 17938 12012 17948 12068
rect 18004 12012 18732 12068
rect 18788 12012 20188 12068
rect 24882 12012 24892 12068
rect 24948 12012 27244 12068
rect 27300 12012 27310 12068
rect 3378 11900 3388 11956
rect 3444 11900 5964 11956
rect 6020 11900 6030 11956
rect 6850 11788 6860 11844
rect 6916 11788 7868 11844
rect 7924 11788 9884 11844
rect 9940 11788 9950 11844
rect 5864 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6148 11788
rect 15188 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15472 11788
rect 24512 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24796 11788
rect 33836 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34120 11788
rect 1586 11676 1596 11732
rect 1652 11676 2380 11732
rect 2436 11676 2446 11732
rect 8082 11676 8092 11732
rect 8148 11676 10668 11732
rect 10724 11676 10734 11732
rect 11554 11676 11564 11732
rect 11620 11676 12236 11732
rect 12292 11676 12302 11732
rect 26898 11676 26908 11732
rect 26964 11676 30268 11732
rect 30324 11676 30334 11732
rect 15698 11564 15708 11620
rect 15764 11564 16940 11620
rect 16996 11564 17006 11620
rect 19058 11564 19068 11620
rect 19124 11564 19516 11620
rect 19572 11564 19582 11620
rect 22978 11564 22988 11620
rect 23044 11564 26124 11620
rect 26180 11564 26190 11620
rect 26450 11564 26460 11620
rect 26516 11564 26908 11620
rect 27570 11564 27580 11620
rect 27636 11564 29708 11620
rect 29764 11564 29774 11620
rect 32386 11564 32396 11620
rect 32452 11564 34524 11620
rect 34580 11564 34590 11620
rect 20178 11452 20188 11508
rect 20244 11452 22428 11508
rect 22484 11452 22494 11508
rect 26852 11396 26908 11564
rect 39200 11508 40000 11536
rect 38098 11452 38108 11508
rect 38164 11452 40000 11508
rect 39200 11424 40000 11452
rect 26852 11340 36988 11396
rect 37044 11340 37054 11396
rect 5506 11228 5516 11284
rect 5572 11228 7532 11284
rect 7588 11228 7598 11284
rect 9650 11228 9660 11284
rect 9716 11228 12124 11284
rect 12180 11228 12190 11284
rect 19282 11228 19292 11284
rect 19348 11228 19358 11284
rect 19618 11228 19628 11284
rect 19684 11228 23548 11284
rect 23604 11228 23614 11284
rect 34178 11228 34188 11284
rect 34244 11228 34524 11284
rect 34580 11228 34590 11284
rect 19292 11172 19348 11228
rect 2258 11116 2268 11172
rect 2324 11116 6412 11172
rect 6468 11116 6478 11172
rect 10098 11116 10108 11172
rect 10164 11116 11004 11172
rect 11060 11116 11070 11172
rect 12226 11116 12236 11172
rect 12292 11116 12908 11172
rect 12964 11116 12974 11172
rect 18162 11116 18172 11172
rect 18228 11116 20636 11172
rect 20692 11116 20702 11172
rect 26562 11116 26572 11172
rect 26628 11116 29596 11172
rect 29652 11116 29662 11172
rect 31042 11116 31052 11172
rect 31108 11116 34300 11172
rect 34356 11116 34366 11172
rect 35158 11116 35196 11172
rect 35252 11116 35756 11172
rect 35812 11116 35822 11172
rect 10526 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10810 11004
rect 19850 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20134 11004
rect 29174 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29458 11004
rect 38498 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38782 11004
rect 17378 10892 17388 10948
rect 17444 10892 19628 10948
rect 19684 10892 19694 10948
rect 39200 10836 40000 10864
rect 8194 10780 8204 10836
rect 8260 10780 8764 10836
rect 8820 10780 8830 10836
rect 36418 10780 36428 10836
rect 36484 10780 38332 10836
rect 38388 10780 40000 10836
rect 39200 10752 40000 10780
rect 2482 10668 2492 10724
rect 2548 10668 4732 10724
rect 4788 10668 4798 10724
rect 13794 10668 13804 10724
rect 13860 10668 17388 10724
rect 17444 10668 17454 10724
rect 18274 10668 18284 10724
rect 18340 10668 20188 10724
rect 20244 10668 20254 10724
rect 32498 10668 32508 10724
rect 32564 10668 37548 10724
rect 37604 10668 37614 10724
rect 8418 10556 8428 10612
rect 8484 10556 8764 10612
rect 8820 10556 8830 10612
rect 12450 10556 12460 10612
rect 12516 10556 12526 10612
rect 13570 10556 13580 10612
rect 13636 10556 14924 10612
rect 14980 10556 16492 10612
rect 16548 10556 16558 10612
rect 31266 10556 31276 10612
rect 31332 10556 33628 10612
rect 33684 10556 33694 10612
rect 12460 10500 12516 10556
rect 5282 10444 5292 10500
rect 5348 10444 6748 10500
rect 6804 10444 6814 10500
rect 11778 10444 11788 10500
rect 11844 10444 12516 10500
rect 15586 10444 15596 10500
rect 15652 10444 17612 10500
rect 17668 10444 17678 10500
rect 19730 10444 19740 10500
rect 19796 10444 21980 10500
rect 22036 10444 22046 10500
rect 23874 10444 23884 10500
rect 23940 10444 26236 10500
rect 26292 10444 26302 10500
rect 27234 10444 27244 10500
rect 27300 10444 35420 10500
rect 35476 10444 35486 10500
rect 13906 10332 13916 10388
rect 13972 10332 15932 10388
rect 15988 10332 15998 10388
rect 27010 10332 27020 10388
rect 27076 10332 36652 10388
rect 36708 10332 36718 10388
rect 35970 10220 35980 10276
rect 36036 10220 36540 10276
rect 36596 10220 36606 10276
rect 5864 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6148 10220
rect 15188 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15472 10220
rect 24512 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24796 10220
rect 33836 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34120 10220
rect 39200 10164 40000 10192
rect 8978 10108 8988 10164
rect 9044 10108 9660 10164
rect 9716 10108 9726 10164
rect 11106 10108 11116 10164
rect 11172 10108 12460 10164
rect 12516 10108 12526 10164
rect 31602 10108 31612 10164
rect 31668 10108 33292 10164
rect 33348 10108 33358 10164
rect 34188 10108 36988 10164
rect 37044 10108 37054 10164
rect 37772 10108 40000 10164
rect 34188 10052 34244 10108
rect 37772 10052 37828 10108
rect 39200 10080 40000 10108
rect 4722 9996 4732 10052
rect 4788 9996 6524 10052
rect 6580 9996 6590 10052
rect 9202 9996 9212 10052
rect 9268 9996 11900 10052
rect 11956 9996 11966 10052
rect 20290 9996 20300 10052
rect 20356 9996 23548 10052
rect 23604 9996 23614 10052
rect 34066 9996 34076 10052
rect 34132 9996 34244 10052
rect 37762 9996 37772 10052
rect 37828 9996 37838 10052
rect 4946 9884 4956 9940
rect 5012 9884 5404 9940
rect 5460 9884 5470 9940
rect 14018 9884 14028 9940
rect 14084 9884 19292 9940
rect 19348 9884 19358 9940
rect 33842 9884 33852 9940
rect 33908 9884 34748 9940
rect 34804 9884 34814 9940
rect 29586 9772 29596 9828
rect 29652 9772 35756 9828
rect 35812 9772 35822 9828
rect 28242 9660 28252 9716
rect 28308 9660 31948 9716
rect 32004 9660 32014 9716
rect 32284 9660 34748 9716
rect 34804 9660 34814 9716
rect 32284 9604 32340 9660
rect 29698 9548 29708 9604
rect 29764 9548 32340 9604
rect 33394 9548 33404 9604
rect 33460 9548 36988 9604
rect 37044 9548 37054 9604
rect 39200 9492 40000 9520
rect 34934 9436 34972 9492
rect 35028 9436 35038 9492
rect 38892 9436 40000 9492
rect 10526 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10810 9436
rect 19850 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20134 9436
rect 29174 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29458 9436
rect 38498 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38782 9436
rect 11778 9324 11788 9380
rect 11844 9324 14364 9380
rect 14420 9324 14430 9380
rect 38892 9268 38948 9436
rect 39200 9408 40000 9436
rect 31490 9212 31500 9268
rect 31556 9212 32956 9268
rect 33012 9212 33022 9268
rect 37762 9212 37772 9268
rect 37828 9212 38948 9268
rect 31154 9100 31164 9156
rect 31220 9100 33628 9156
rect 33684 9100 33694 9156
rect 11218 8988 11228 9044
rect 11284 8988 15036 9044
rect 15092 8988 15102 9044
rect 27570 8988 27580 9044
rect 27636 8988 34748 9044
rect 34804 8988 34814 9044
rect 3042 8876 3052 8932
rect 3108 8876 5628 8932
rect 5684 8876 7084 8932
rect 7140 8876 7150 8932
rect 26786 8876 26796 8932
rect 26852 8876 28924 8932
rect 28980 8876 28990 8932
rect 32722 8876 32732 8932
rect 32788 8876 35532 8932
rect 35588 8876 35598 8932
rect 39200 8820 40000 8848
rect 30930 8764 30940 8820
rect 30996 8764 40000 8820
rect 39200 8736 40000 8764
rect 5864 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6148 8652
rect 15188 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15472 8652
rect 24512 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24796 8652
rect 33836 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34120 8652
rect 8754 8540 8764 8596
rect 8820 8540 10332 8596
rect 10388 8540 10398 8596
rect 27906 8540 27916 8596
rect 27972 8540 32396 8596
rect 32452 8540 32462 8596
rect 32946 8540 32956 8596
rect 33012 8540 33628 8596
rect 33684 8540 33694 8596
rect 27682 8428 27692 8484
rect 27748 8428 37884 8484
rect 37940 8428 37950 8484
rect 2258 8316 2268 8372
rect 2324 8316 3612 8372
rect 3668 8316 3678 8372
rect 7298 8316 7308 8372
rect 7364 8316 8876 8372
rect 8932 8316 8942 8372
rect 9090 8316 9100 8372
rect 9156 8316 11788 8372
rect 11844 8316 11854 8372
rect 36082 8316 36092 8372
rect 36148 8316 37100 8372
rect 37156 8316 37166 8372
rect 29810 8204 29820 8260
rect 29876 8204 36316 8260
rect 36372 8204 36382 8260
rect 39200 8148 40000 8176
rect 5170 8092 5180 8148
rect 5236 8092 6076 8148
rect 6132 8092 6142 8148
rect 38098 8092 38108 8148
rect 38164 8092 40000 8148
rect 39200 8064 40000 8092
rect 30034 7980 30044 8036
rect 30100 7980 36988 8036
rect 37044 7980 37054 8036
rect 33506 7868 33516 7924
rect 33572 7868 35196 7924
rect 35252 7868 35262 7924
rect 10526 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10810 7868
rect 19850 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20134 7868
rect 29174 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29458 7868
rect 38498 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38782 7868
rect 6626 7644 6636 7700
rect 6692 7644 10668 7700
rect 10724 7644 10734 7700
rect 35074 7532 35084 7588
rect 35140 7532 36652 7588
rect 36708 7532 36718 7588
rect 39200 7476 40000 7504
rect 14690 7420 14700 7476
rect 14756 7420 15708 7476
rect 15764 7420 15774 7476
rect 27346 7420 27356 7476
rect 27412 7420 36988 7476
rect 37044 7420 37054 7476
rect 37762 7420 37772 7476
rect 37828 7420 40000 7476
rect 39200 7392 40000 7420
rect 7746 7308 7756 7364
rect 7812 7308 10556 7364
rect 10612 7308 10622 7364
rect 11666 7308 11676 7364
rect 11732 7308 13356 7364
rect 13412 7308 13422 7364
rect 28690 7308 28700 7364
rect 28756 7308 32844 7364
rect 32900 7308 32910 7364
rect 34934 7308 34972 7364
rect 35028 7308 35038 7364
rect 31826 7196 31836 7252
rect 31892 7196 33068 7252
rect 33124 7196 33134 7252
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 28578 6972 28588 7028
rect 28644 6972 30604 7028
rect 30660 6972 30670 7028
rect 31490 6972 31500 7028
rect 31556 6972 32172 7028
rect 32228 6972 32238 7028
rect 26852 6860 27244 6916
rect 27300 6860 31220 6916
rect 33282 6860 33292 6916
rect 33348 6860 34076 6916
rect 34132 6860 34142 6916
rect 34738 6860 34748 6916
rect 34804 6860 36428 6916
rect 36484 6860 36494 6916
rect 26852 6692 26908 6860
rect 31164 6804 31220 6860
rect 39200 6804 40000 6832
rect 28802 6748 28812 6804
rect 28868 6748 30492 6804
rect 30548 6748 30558 6804
rect 31164 6748 40000 6804
rect 39200 6720 40000 6748
rect 26674 6636 26684 6692
rect 26740 6636 26908 6692
rect 27682 6636 27692 6692
rect 27748 6636 29260 6692
rect 29316 6636 37660 6692
rect 37716 6636 37726 6692
rect 26338 6524 26348 6580
rect 26404 6524 34972 6580
rect 35028 6524 35038 6580
rect 33394 6412 33404 6468
rect 33460 6412 36988 6468
rect 37044 6412 37054 6468
rect 10526 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10810 6300
rect 19850 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20134 6300
rect 29174 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29458 6300
rect 38498 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38782 6300
rect 39200 6132 40000 6160
rect 27682 6076 27692 6132
rect 27748 6076 32956 6132
rect 33012 6076 33022 6132
rect 37538 6076 37548 6132
rect 37604 6076 40000 6132
rect 39200 6048 40000 6076
rect 5282 5964 5292 6020
rect 5348 5964 6860 6020
rect 6916 5964 6926 6020
rect 26562 5964 26572 6020
rect 26628 5964 28028 6020
rect 28084 5964 28094 6020
rect 28354 5964 28364 6020
rect 28420 5964 29596 6020
rect 29652 5964 35868 6020
rect 35924 5964 35934 6020
rect 29698 5852 29708 5908
rect 29764 5852 31948 5908
rect 32004 5852 32014 5908
rect 27682 5740 27692 5796
rect 27748 5740 33852 5796
rect 33908 5740 33918 5796
rect 26450 5628 26460 5684
rect 26516 5628 27468 5684
rect 27524 5628 34244 5684
rect 36306 5628 36316 5684
rect 36372 5628 37436 5684
rect 37492 5628 37502 5684
rect 5864 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6148 5516
rect 15188 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15472 5516
rect 24512 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24796 5516
rect 33836 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34120 5516
rect 34188 5460 34244 5628
rect 39200 5460 40000 5488
rect 27122 5404 27132 5460
rect 27188 5404 33180 5460
rect 33236 5404 33246 5460
rect 34188 5404 40000 5460
rect 39200 5376 40000 5404
rect 26898 5292 26908 5348
rect 26964 5292 29372 5348
rect 29428 5292 29438 5348
rect 30370 5292 30380 5348
rect 30436 5292 36988 5348
rect 37044 5292 37054 5348
rect 31938 5180 31948 5236
rect 32004 5180 34524 5236
rect 34580 5180 34590 5236
rect 32050 5068 32060 5124
rect 32116 5068 35644 5124
rect 35700 5068 35710 5124
rect 30146 4956 30156 5012
rect 30212 4956 37548 5012
rect 37604 4956 37614 5012
rect 26338 4844 26348 4900
rect 26404 4844 28700 4900
rect 28756 4844 28766 4900
rect 29250 4844 29260 4900
rect 29316 4844 30324 4900
rect 30482 4844 30492 4900
rect 30548 4844 38948 4900
rect 30268 4788 30324 4844
rect 38892 4788 38948 4844
rect 39200 4788 40000 4816
rect 30268 4732 32284 4788
rect 32340 4732 32350 4788
rect 38892 4732 40000 4788
rect 10526 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10810 4732
rect 19850 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20134 4732
rect 29174 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29458 4732
rect 38498 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38782 4732
rect 39200 4704 40000 4732
rect 27234 4620 27244 4676
rect 27300 4620 28364 4676
rect 28420 4620 28430 4676
rect 30594 4620 30604 4676
rect 30660 4620 35980 4676
rect 36036 4620 36046 4676
rect 36194 4620 36204 4676
rect 36260 4620 37772 4676
rect 37828 4620 37838 4676
rect 26674 4508 26684 4564
rect 26740 4508 28084 4564
rect 28242 4508 28252 4564
rect 28308 4508 29036 4564
rect 29092 4508 29102 4564
rect 36866 4508 36876 4564
rect 36932 4508 36942 4564
rect 28028 4452 28084 4508
rect 36876 4452 36932 4508
rect 26114 4396 26124 4452
rect 26180 4396 27132 4452
rect 27188 4396 27198 4452
rect 28028 4396 36932 4452
rect 29362 4284 29372 4340
rect 29428 4284 30940 4340
rect 30996 4284 31006 4340
rect 31164 4284 38108 4340
rect 38164 4284 38174 4340
rect 31164 4228 31220 4284
rect 29026 4172 29036 4228
rect 29092 4172 31220 4228
rect 31602 4172 31612 4228
rect 31668 4172 33516 4228
rect 33572 4172 33582 4228
rect 34178 4172 34188 4228
rect 34244 4172 35140 4228
rect 35084 4116 35140 4172
rect 39200 4116 40000 4144
rect 27122 4060 27132 4116
rect 27188 4060 34636 4116
rect 34692 4060 34702 4116
rect 35084 4060 40000 4116
rect 39200 4032 40000 4060
rect 5864 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6148 3948
rect 15188 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15472 3948
rect 24512 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24796 3948
rect 33836 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34120 3948
rect 27682 3724 27692 3780
rect 27748 3724 29708 3780
rect 29764 3724 30940 3780
rect 30996 3724 31006 3780
rect 35186 3724 35196 3780
rect 35252 3724 39676 3780
rect 39732 3724 39742 3780
rect 29586 3612 29596 3668
rect 29652 3612 30492 3668
rect 30548 3612 30558 3668
rect 34962 3612 34972 3668
rect 35028 3612 36428 3668
rect 36484 3612 36494 3668
rect 28018 3500 28028 3556
rect 28084 3500 32172 3556
rect 32228 3500 32238 3556
rect 39200 3444 40000 3472
rect 26114 3388 26124 3444
rect 26180 3388 27580 3444
rect 27636 3388 27646 3444
rect 33030 3388 33068 3444
rect 33124 3388 33134 3444
rect 34738 3388 34748 3444
rect 34804 3388 40000 3444
rect 39200 3360 40000 3388
rect 37314 3276 37324 3332
rect 37380 3276 37884 3332
rect 37940 3276 37950 3332
rect 10526 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10810 3164
rect 19850 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20134 3164
rect 29174 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29458 3164
rect 38498 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38782 3164
rect 39200 2772 40000 2800
rect 35074 2716 35084 2772
rect 35140 2716 40000 2772
rect 39200 2688 40000 2716
rect 39200 2100 40000 2128
rect 35186 2044 35196 2100
rect 35252 2044 40000 2100
rect 39200 2016 40000 2044
rect 39200 1428 40000 1456
rect 37874 1372 37884 1428
rect 37940 1372 40000 1428
rect 39200 1344 40000 1372
rect 33954 1036 33964 1092
rect 34020 1036 34030 1092
rect 33964 756 34020 1036
rect 39200 756 40000 784
rect 33964 700 40000 756
rect 39200 672 40000 700
rect 39200 84 40000 112
rect 37426 28 37436 84
rect 37492 28 40000 84
rect 39200 0 40000 28
<< via3 >>
rect 5874 36820 5930 36876
rect 5978 36820 6034 36876
rect 6082 36820 6138 36876
rect 15198 36820 15254 36876
rect 15302 36820 15358 36876
rect 15406 36820 15462 36876
rect 24522 36820 24578 36876
rect 24626 36820 24682 36876
rect 24730 36820 24786 36876
rect 33846 36820 33902 36876
rect 33950 36820 34006 36876
rect 34054 36820 34110 36876
rect 10536 36036 10592 36092
rect 10640 36036 10696 36092
rect 10744 36036 10800 36092
rect 19860 36036 19916 36092
rect 19964 36036 20020 36092
rect 20068 36036 20124 36092
rect 29184 36036 29240 36092
rect 29288 36036 29344 36092
rect 29392 36036 29448 36092
rect 38508 36036 38564 36092
rect 38612 36036 38668 36092
rect 38716 36036 38772 36092
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 10536 34468 10592 34524
rect 10640 34468 10696 34524
rect 10744 34468 10800 34524
rect 19860 34468 19916 34524
rect 19964 34468 20020 34524
rect 20068 34468 20124 34524
rect 29184 34468 29240 34524
rect 29288 34468 29344 34524
rect 29392 34468 29448 34524
rect 38508 34468 38564 34524
rect 38612 34468 38668 34524
rect 38716 34468 38772 34524
rect 5874 33684 5930 33740
rect 5978 33684 6034 33740
rect 6082 33684 6138 33740
rect 15198 33684 15254 33740
rect 15302 33684 15358 33740
rect 15406 33684 15462 33740
rect 24522 33684 24578 33740
rect 24626 33684 24682 33740
rect 24730 33684 24786 33740
rect 33846 33684 33902 33740
rect 33950 33684 34006 33740
rect 34054 33684 34110 33740
rect 10536 32900 10592 32956
rect 10640 32900 10696 32956
rect 10744 32900 10800 32956
rect 19860 32900 19916 32956
rect 19964 32900 20020 32956
rect 20068 32900 20124 32956
rect 29184 32900 29240 32956
rect 29288 32900 29344 32956
rect 29392 32900 29448 32956
rect 38508 32900 38564 32956
rect 38612 32900 38668 32956
rect 38716 32900 38772 32956
rect 5874 32116 5930 32172
rect 5978 32116 6034 32172
rect 6082 32116 6138 32172
rect 15198 32116 15254 32172
rect 15302 32116 15358 32172
rect 15406 32116 15462 32172
rect 24522 32116 24578 32172
rect 24626 32116 24682 32172
rect 24730 32116 24786 32172
rect 33846 32116 33902 32172
rect 33950 32116 34006 32172
rect 34054 32116 34110 32172
rect 10536 31332 10592 31388
rect 10640 31332 10696 31388
rect 10744 31332 10800 31388
rect 19860 31332 19916 31388
rect 19964 31332 20020 31388
rect 20068 31332 20124 31388
rect 29184 31332 29240 31388
rect 29288 31332 29344 31388
rect 29392 31332 29448 31388
rect 38508 31332 38564 31388
rect 38612 31332 38668 31388
rect 38716 31332 38772 31388
rect 5874 30548 5930 30604
rect 5978 30548 6034 30604
rect 6082 30548 6138 30604
rect 15198 30548 15254 30604
rect 15302 30548 15358 30604
rect 15406 30548 15462 30604
rect 24522 30548 24578 30604
rect 24626 30548 24682 30604
rect 24730 30548 24786 30604
rect 33846 30548 33902 30604
rect 33950 30548 34006 30604
rect 34054 30548 34110 30604
rect 10536 29764 10592 29820
rect 10640 29764 10696 29820
rect 10744 29764 10800 29820
rect 19860 29764 19916 29820
rect 19964 29764 20020 29820
rect 20068 29764 20124 29820
rect 29184 29764 29240 29820
rect 29288 29764 29344 29820
rect 29392 29764 29448 29820
rect 38508 29764 38564 29820
rect 38612 29764 38668 29820
rect 38716 29764 38772 29820
rect 5874 28980 5930 29036
rect 5978 28980 6034 29036
rect 6082 28980 6138 29036
rect 15198 28980 15254 29036
rect 15302 28980 15358 29036
rect 15406 28980 15462 29036
rect 24522 28980 24578 29036
rect 24626 28980 24682 29036
rect 24730 28980 24786 29036
rect 33846 28980 33902 29036
rect 33950 28980 34006 29036
rect 34054 28980 34110 29036
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 5874 27412 5930 27468
rect 5978 27412 6034 27468
rect 6082 27412 6138 27468
rect 15198 27412 15254 27468
rect 15302 27412 15358 27468
rect 15406 27412 15462 27468
rect 24522 27412 24578 27468
rect 24626 27412 24682 27468
rect 24730 27412 24786 27468
rect 33846 27412 33902 27468
rect 33950 27412 34006 27468
rect 34054 27412 34110 27468
rect 10536 26628 10592 26684
rect 10640 26628 10696 26684
rect 10744 26628 10800 26684
rect 19860 26628 19916 26684
rect 19964 26628 20020 26684
rect 20068 26628 20124 26684
rect 29184 26628 29240 26684
rect 29288 26628 29344 26684
rect 29392 26628 29448 26684
rect 38508 26628 38564 26684
rect 38612 26628 38668 26684
rect 38716 26628 38772 26684
rect 5874 25844 5930 25900
rect 5978 25844 6034 25900
rect 6082 25844 6138 25900
rect 15198 25844 15254 25900
rect 15302 25844 15358 25900
rect 15406 25844 15462 25900
rect 24522 25844 24578 25900
rect 24626 25844 24682 25900
rect 24730 25844 24786 25900
rect 33846 25844 33902 25900
rect 33950 25844 34006 25900
rect 34054 25844 34110 25900
rect 10536 25060 10592 25116
rect 10640 25060 10696 25116
rect 10744 25060 10800 25116
rect 19860 25060 19916 25116
rect 19964 25060 20020 25116
rect 20068 25060 20124 25116
rect 29184 25060 29240 25116
rect 29288 25060 29344 25116
rect 29392 25060 29448 25116
rect 38508 25060 38564 25116
rect 38612 25060 38668 25116
rect 38716 25060 38772 25116
rect 5874 24276 5930 24332
rect 5978 24276 6034 24332
rect 6082 24276 6138 24332
rect 15198 24276 15254 24332
rect 15302 24276 15358 24332
rect 15406 24276 15462 24332
rect 24522 24276 24578 24332
rect 24626 24276 24682 24332
rect 24730 24276 24786 24332
rect 33846 24276 33902 24332
rect 33950 24276 34006 24332
rect 34054 24276 34110 24332
rect 10536 23492 10592 23548
rect 10640 23492 10696 23548
rect 10744 23492 10800 23548
rect 19860 23492 19916 23548
rect 19964 23492 20020 23548
rect 20068 23492 20124 23548
rect 29184 23492 29240 23548
rect 29288 23492 29344 23548
rect 29392 23492 29448 23548
rect 38508 23492 38564 23548
rect 38612 23492 38668 23548
rect 38716 23492 38772 23548
rect 5874 22708 5930 22764
rect 5978 22708 6034 22764
rect 6082 22708 6138 22764
rect 15198 22708 15254 22764
rect 15302 22708 15358 22764
rect 15406 22708 15462 22764
rect 24522 22708 24578 22764
rect 24626 22708 24682 22764
rect 24730 22708 24786 22764
rect 33846 22708 33902 22764
rect 33950 22708 34006 22764
rect 34054 22708 34110 22764
rect 10536 21924 10592 21980
rect 10640 21924 10696 21980
rect 10744 21924 10800 21980
rect 19860 21924 19916 21980
rect 19964 21924 20020 21980
rect 20068 21924 20124 21980
rect 29184 21924 29240 21980
rect 29288 21924 29344 21980
rect 29392 21924 29448 21980
rect 38508 21924 38564 21980
rect 38612 21924 38668 21980
rect 38716 21924 38772 21980
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20356 10592 20412
rect 10640 20356 10696 20412
rect 10744 20356 10800 20412
rect 19860 20356 19916 20412
rect 19964 20356 20020 20412
rect 20068 20356 20124 20412
rect 29184 20356 29240 20412
rect 29288 20356 29344 20412
rect 29392 20356 29448 20412
rect 38508 20356 38564 20412
rect 38612 20356 38668 20412
rect 38716 20356 38772 20412
rect 5874 19572 5930 19628
rect 5978 19572 6034 19628
rect 6082 19572 6138 19628
rect 15198 19572 15254 19628
rect 15302 19572 15358 19628
rect 15406 19572 15462 19628
rect 24522 19572 24578 19628
rect 24626 19572 24682 19628
rect 24730 19572 24786 19628
rect 33846 19572 33902 19628
rect 33950 19572 34006 19628
rect 34054 19572 34110 19628
rect 10536 18788 10592 18844
rect 10640 18788 10696 18844
rect 10744 18788 10800 18844
rect 19860 18788 19916 18844
rect 19964 18788 20020 18844
rect 20068 18788 20124 18844
rect 29184 18788 29240 18844
rect 29288 18788 29344 18844
rect 29392 18788 29448 18844
rect 38508 18788 38564 18844
rect 38612 18788 38668 18844
rect 38716 18788 38772 18844
rect 5874 18004 5930 18060
rect 5978 18004 6034 18060
rect 6082 18004 6138 18060
rect 15198 18004 15254 18060
rect 15302 18004 15358 18060
rect 15406 18004 15462 18060
rect 24522 18004 24578 18060
rect 24626 18004 24682 18060
rect 24730 18004 24786 18060
rect 33846 18004 33902 18060
rect 33950 18004 34006 18060
rect 34054 18004 34110 18060
rect 10536 17220 10592 17276
rect 10640 17220 10696 17276
rect 10744 17220 10800 17276
rect 19860 17220 19916 17276
rect 19964 17220 20020 17276
rect 20068 17220 20124 17276
rect 29184 17220 29240 17276
rect 29288 17220 29344 17276
rect 29392 17220 29448 17276
rect 38508 17220 38564 17276
rect 38612 17220 38668 17276
rect 38716 17220 38772 17276
rect 29708 16604 29764 16660
rect 5874 16436 5930 16492
rect 5978 16436 6034 16492
rect 6082 16436 6138 16492
rect 15198 16436 15254 16492
rect 15302 16436 15358 16492
rect 15406 16436 15462 16492
rect 24522 16436 24578 16492
rect 24626 16436 24682 16492
rect 24730 16436 24786 16492
rect 33846 16436 33902 16492
rect 33950 16436 34006 16492
rect 34054 16436 34110 16492
rect 10536 15652 10592 15708
rect 10640 15652 10696 15708
rect 10744 15652 10800 15708
rect 19860 15652 19916 15708
rect 19964 15652 20020 15708
rect 20068 15652 20124 15708
rect 29184 15652 29240 15708
rect 29288 15652 29344 15708
rect 29392 15652 29448 15708
rect 38508 15652 38564 15708
rect 38612 15652 38668 15708
rect 38716 15652 38772 15708
rect 32956 15148 33012 15204
rect 33516 15148 33572 15204
rect 5874 14868 5930 14924
rect 5978 14868 6034 14924
rect 6082 14868 6138 14924
rect 15198 14868 15254 14924
rect 15302 14868 15358 14924
rect 15406 14868 15462 14924
rect 24522 14868 24578 14924
rect 24626 14868 24682 14924
rect 24730 14868 24786 14924
rect 33846 14868 33902 14924
rect 33950 14868 34006 14924
rect 34054 14868 34110 14924
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 5874 13300 5930 13356
rect 5978 13300 6034 13356
rect 6082 13300 6138 13356
rect 15198 13300 15254 13356
rect 15302 13300 15358 13356
rect 15406 13300 15462 13356
rect 24522 13300 24578 13356
rect 24626 13300 24682 13356
rect 24730 13300 24786 13356
rect 33846 13300 33902 13356
rect 33950 13300 34006 13356
rect 34054 13300 34110 13356
rect 10536 12516 10592 12572
rect 10640 12516 10696 12572
rect 10744 12516 10800 12572
rect 19860 12516 19916 12572
rect 19964 12516 20020 12572
rect 20068 12516 20124 12572
rect 29184 12516 29240 12572
rect 29288 12516 29344 12572
rect 29392 12516 29448 12572
rect 38508 12516 38564 12572
rect 38612 12516 38668 12572
rect 38716 12516 38772 12572
rect 5874 11732 5930 11788
rect 5978 11732 6034 11788
rect 6082 11732 6138 11788
rect 15198 11732 15254 11788
rect 15302 11732 15358 11788
rect 15406 11732 15462 11788
rect 24522 11732 24578 11788
rect 24626 11732 24682 11788
rect 24730 11732 24786 11788
rect 33846 11732 33902 11788
rect 33950 11732 34006 11788
rect 34054 11732 34110 11788
rect 35196 11116 35252 11172
rect 10536 10948 10592 11004
rect 10640 10948 10696 11004
rect 10744 10948 10800 11004
rect 19860 10948 19916 11004
rect 19964 10948 20020 11004
rect 20068 10948 20124 11004
rect 29184 10948 29240 11004
rect 29288 10948 29344 11004
rect 29392 10948 29448 11004
rect 38508 10948 38564 11004
rect 38612 10948 38668 11004
rect 38716 10948 38772 11004
rect 5874 10164 5930 10220
rect 5978 10164 6034 10220
rect 6082 10164 6138 10220
rect 15198 10164 15254 10220
rect 15302 10164 15358 10220
rect 15406 10164 15462 10220
rect 24522 10164 24578 10220
rect 24626 10164 24682 10220
rect 24730 10164 24786 10220
rect 33846 10164 33902 10220
rect 33950 10164 34006 10220
rect 34054 10164 34110 10220
rect 29708 9548 29764 9604
rect 34972 9436 35028 9492
rect 10536 9380 10592 9436
rect 10640 9380 10696 9436
rect 10744 9380 10800 9436
rect 19860 9380 19916 9436
rect 19964 9380 20020 9436
rect 20068 9380 20124 9436
rect 29184 9380 29240 9436
rect 29288 9380 29344 9436
rect 29392 9380 29448 9436
rect 38508 9380 38564 9436
rect 38612 9380 38668 9436
rect 38716 9380 38772 9436
rect 5874 8596 5930 8652
rect 5978 8596 6034 8652
rect 6082 8596 6138 8652
rect 15198 8596 15254 8652
rect 15302 8596 15358 8652
rect 15406 8596 15462 8652
rect 24522 8596 24578 8652
rect 24626 8596 24682 8652
rect 24730 8596 24786 8652
rect 33846 8596 33902 8652
rect 33950 8596 34006 8652
rect 34054 8596 34110 8652
rect 33516 7868 33572 7924
rect 10536 7812 10592 7868
rect 10640 7812 10696 7868
rect 10744 7812 10800 7868
rect 19860 7812 19916 7868
rect 19964 7812 20020 7868
rect 20068 7812 20124 7868
rect 29184 7812 29240 7868
rect 29288 7812 29344 7868
rect 29392 7812 29448 7868
rect 38508 7812 38564 7868
rect 38612 7812 38668 7868
rect 38716 7812 38772 7868
rect 34972 7308 35028 7364
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6244 10592 6300
rect 10640 6244 10696 6300
rect 10744 6244 10800 6300
rect 19860 6244 19916 6300
rect 19964 6244 20020 6300
rect 20068 6244 20124 6300
rect 29184 6244 29240 6300
rect 29288 6244 29344 6300
rect 29392 6244 29448 6300
rect 38508 6244 38564 6300
rect 38612 6244 38668 6300
rect 38716 6244 38772 6300
rect 5874 5460 5930 5516
rect 5978 5460 6034 5516
rect 6082 5460 6138 5516
rect 15198 5460 15254 5516
rect 15302 5460 15358 5516
rect 15406 5460 15462 5516
rect 24522 5460 24578 5516
rect 24626 5460 24682 5516
rect 24730 5460 24786 5516
rect 33846 5460 33902 5516
rect 33950 5460 34006 5516
rect 34054 5460 34110 5516
rect 10536 4676 10592 4732
rect 10640 4676 10696 4732
rect 10744 4676 10800 4732
rect 19860 4676 19916 4732
rect 19964 4676 20020 4732
rect 20068 4676 20124 4732
rect 29184 4676 29240 4732
rect 29288 4676 29344 4732
rect 29392 4676 29448 4732
rect 38508 4676 38564 4732
rect 38612 4676 38668 4732
rect 38716 4676 38772 4732
rect 5874 3892 5930 3948
rect 5978 3892 6034 3948
rect 6082 3892 6138 3948
rect 15198 3892 15254 3948
rect 15302 3892 15358 3948
rect 15406 3892 15462 3948
rect 24522 3892 24578 3948
rect 24626 3892 24682 3948
rect 24730 3892 24786 3948
rect 33846 3892 33902 3948
rect 33950 3892 34006 3948
rect 34054 3892 34110 3948
rect 33068 3388 33124 3444
rect 10536 3108 10592 3164
rect 10640 3108 10696 3164
rect 10744 3108 10800 3164
rect 19860 3108 19916 3164
rect 19964 3108 20020 3164
rect 20068 3108 20124 3164
rect 29184 3108 29240 3164
rect 29288 3108 29344 3164
rect 29392 3108 29448 3164
rect 38508 3108 38564 3164
rect 38612 3108 38668 3164
rect 38716 3108 38772 3164
rect 35196 2044 35252 2100
<< metal4 >>
rect 5846 36876 6166 36908
rect 5846 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6166 36876
rect 5846 35308 6166 36820
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33740 6166 35252
rect 5846 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6166 33740
rect 5846 32172 6166 33684
rect 5846 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6166 32172
rect 5846 30604 6166 32116
rect 5846 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6166 30604
rect 5846 29036 6166 30548
rect 5846 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6166 29036
rect 5846 27468 6166 28980
rect 5846 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6166 27468
rect 5846 25900 6166 27412
rect 5846 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6166 25900
rect 5846 24332 6166 25844
rect 5846 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6166 24332
rect 5846 22764 6166 24276
rect 5846 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6166 22764
rect 5846 21196 6166 22708
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19628 6166 21140
rect 5846 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6166 19628
rect 5846 18060 6166 19572
rect 5846 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6166 18060
rect 5846 16492 6166 18004
rect 5846 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6166 16492
rect 5846 14924 6166 16436
rect 5846 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6166 14924
rect 5846 13356 6166 14868
rect 5846 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6166 13356
rect 5846 11788 6166 13300
rect 5846 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6166 11788
rect 5846 10220 6166 11732
rect 5846 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6166 10220
rect 5846 8652 6166 10164
rect 5846 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6166 8652
rect 5846 7084 6166 8596
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5516 6166 7028
rect 5846 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6166 5516
rect 5846 3948 6166 5460
rect 5846 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6166 3948
rect 5846 3076 6166 3892
rect 10508 36092 10828 36908
rect 10508 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10828 36092
rect 10508 34524 10828 36036
rect 10508 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10828 34524
rect 10508 32956 10828 34468
rect 10508 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10828 32956
rect 10508 31388 10828 32900
rect 10508 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10828 31388
rect 10508 29820 10828 31332
rect 10508 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10828 29820
rect 10508 28252 10828 29764
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26684 10828 28196
rect 10508 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10828 26684
rect 10508 25116 10828 26628
rect 10508 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10828 25116
rect 10508 23548 10828 25060
rect 10508 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10828 23548
rect 10508 21980 10828 23492
rect 10508 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10828 21980
rect 10508 20412 10828 21924
rect 10508 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10828 20412
rect 10508 18844 10828 20356
rect 10508 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10828 18844
rect 10508 17276 10828 18788
rect 10508 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10828 17276
rect 10508 15708 10828 17220
rect 10508 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10828 15708
rect 10508 14140 10828 15652
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 10508 12572 10828 14084
rect 10508 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10828 12572
rect 10508 11004 10828 12516
rect 10508 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10828 11004
rect 10508 9436 10828 10948
rect 10508 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10828 9436
rect 10508 7868 10828 9380
rect 10508 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10828 7868
rect 10508 6300 10828 7812
rect 10508 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10828 6300
rect 10508 4732 10828 6244
rect 10508 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10828 4732
rect 10508 3164 10828 4676
rect 10508 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10828 3164
rect 10508 3076 10828 3108
rect 15170 36876 15490 36908
rect 15170 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15490 36876
rect 15170 35308 15490 36820
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33740 15490 35252
rect 15170 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15490 33740
rect 15170 32172 15490 33684
rect 15170 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15490 32172
rect 15170 30604 15490 32116
rect 15170 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15490 30604
rect 15170 29036 15490 30548
rect 15170 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15490 29036
rect 15170 27468 15490 28980
rect 15170 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15490 27468
rect 15170 25900 15490 27412
rect 15170 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15490 25900
rect 15170 24332 15490 25844
rect 15170 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15490 24332
rect 15170 22764 15490 24276
rect 15170 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15490 22764
rect 15170 21196 15490 22708
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19628 15490 21140
rect 15170 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15490 19628
rect 15170 18060 15490 19572
rect 15170 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15490 18060
rect 15170 16492 15490 18004
rect 15170 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15490 16492
rect 15170 14924 15490 16436
rect 15170 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15490 14924
rect 15170 13356 15490 14868
rect 15170 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15490 13356
rect 15170 11788 15490 13300
rect 15170 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15490 11788
rect 15170 10220 15490 11732
rect 15170 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15490 10220
rect 15170 8652 15490 10164
rect 15170 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15490 8652
rect 15170 7084 15490 8596
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5516 15490 7028
rect 15170 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15490 5516
rect 15170 3948 15490 5460
rect 15170 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15490 3948
rect 15170 3076 15490 3892
rect 19832 36092 20152 36908
rect 19832 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20152 36092
rect 19832 34524 20152 36036
rect 19832 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20152 34524
rect 19832 32956 20152 34468
rect 19832 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20152 32956
rect 19832 31388 20152 32900
rect 19832 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20152 31388
rect 19832 29820 20152 31332
rect 19832 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20152 29820
rect 19832 28252 20152 29764
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26684 20152 28196
rect 19832 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20152 26684
rect 19832 25116 20152 26628
rect 19832 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20152 25116
rect 19832 23548 20152 25060
rect 19832 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20152 23548
rect 19832 21980 20152 23492
rect 19832 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20152 21980
rect 19832 20412 20152 21924
rect 19832 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20152 20412
rect 19832 18844 20152 20356
rect 19832 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20152 18844
rect 19832 17276 20152 18788
rect 19832 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20152 17276
rect 19832 15708 20152 17220
rect 19832 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20152 15708
rect 19832 14140 20152 15652
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12572 20152 14084
rect 19832 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20152 12572
rect 19832 11004 20152 12516
rect 19832 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20152 11004
rect 19832 9436 20152 10948
rect 19832 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20152 9436
rect 19832 7868 20152 9380
rect 19832 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20152 7868
rect 19832 6300 20152 7812
rect 19832 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20152 6300
rect 19832 4732 20152 6244
rect 19832 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20152 4732
rect 19832 3164 20152 4676
rect 19832 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20152 3164
rect 19832 3076 20152 3108
rect 24494 36876 24814 36908
rect 24494 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24814 36876
rect 24494 35308 24814 36820
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33740 24814 35252
rect 24494 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24814 33740
rect 24494 32172 24814 33684
rect 24494 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24814 32172
rect 24494 30604 24814 32116
rect 24494 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24814 30604
rect 24494 29036 24814 30548
rect 24494 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24814 29036
rect 24494 27468 24814 28980
rect 24494 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24814 27468
rect 24494 25900 24814 27412
rect 24494 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24814 25900
rect 24494 24332 24814 25844
rect 24494 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24814 24332
rect 24494 22764 24814 24276
rect 24494 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24814 22764
rect 24494 21196 24814 22708
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19628 24814 21140
rect 24494 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24814 19628
rect 24494 18060 24814 19572
rect 24494 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24814 18060
rect 24494 16492 24814 18004
rect 24494 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24814 16492
rect 24494 14924 24814 16436
rect 24494 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24814 14924
rect 24494 13356 24814 14868
rect 24494 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24814 13356
rect 24494 11788 24814 13300
rect 24494 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24814 11788
rect 24494 10220 24814 11732
rect 24494 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24814 10220
rect 24494 8652 24814 10164
rect 24494 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24814 8652
rect 24494 7084 24814 8596
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5516 24814 7028
rect 24494 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24814 5516
rect 24494 3948 24814 5460
rect 24494 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24814 3948
rect 24494 3076 24814 3892
rect 29156 36092 29476 36908
rect 29156 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29476 36092
rect 29156 34524 29476 36036
rect 29156 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29476 34524
rect 29156 32956 29476 34468
rect 29156 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29476 32956
rect 29156 31388 29476 32900
rect 29156 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29476 31388
rect 29156 29820 29476 31332
rect 29156 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29476 29820
rect 29156 28252 29476 29764
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26684 29476 28196
rect 29156 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29476 26684
rect 29156 25116 29476 26628
rect 29156 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29476 25116
rect 29156 23548 29476 25060
rect 29156 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29476 23548
rect 29156 21980 29476 23492
rect 29156 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29476 21980
rect 29156 20412 29476 21924
rect 29156 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29476 20412
rect 29156 18844 29476 20356
rect 29156 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29476 18844
rect 29156 17276 29476 18788
rect 29156 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29476 17276
rect 29156 15708 29476 17220
rect 33818 36876 34138 36908
rect 33818 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34138 36876
rect 33818 35308 34138 36820
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33740 34138 35252
rect 33818 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34138 33740
rect 33818 32172 34138 33684
rect 33818 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34138 32172
rect 33818 30604 34138 32116
rect 33818 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34138 30604
rect 33818 29036 34138 30548
rect 33818 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34138 29036
rect 33818 27468 34138 28980
rect 33818 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34138 27468
rect 33818 25900 34138 27412
rect 33818 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34138 25900
rect 33818 24332 34138 25844
rect 33818 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34138 24332
rect 33818 22764 34138 24276
rect 33818 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34138 22764
rect 33818 21196 34138 22708
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19628 34138 21140
rect 33818 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34138 19628
rect 33818 18060 34138 19572
rect 33818 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34138 18060
rect 29156 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29476 15708
rect 29156 14140 29476 15652
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12572 29476 14084
rect 29156 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29476 12572
rect 29156 11004 29476 12516
rect 29156 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29476 11004
rect 29156 9436 29476 10948
rect 29708 16660 29764 16670
rect 29708 9604 29764 16604
rect 33818 16492 34138 18004
rect 33818 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34138 16492
rect 32956 15204 33012 15214
rect 33516 15204 33572 15214
rect 32956 15092 33124 15148
rect 29708 9538 29764 9548
rect 29156 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29476 9436
rect 29156 7868 29476 9380
rect 29156 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29476 7868
rect 29156 6300 29476 7812
rect 29156 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29476 6300
rect 29156 4732 29476 6244
rect 29156 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29476 4732
rect 29156 3164 29476 4676
rect 33068 3444 33124 15092
rect 33516 7924 33572 15148
rect 33516 7858 33572 7868
rect 33818 14924 34138 16436
rect 33818 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34138 14924
rect 33818 13356 34138 14868
rect 33818 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34138 13356
rect 33818 11788 34138 13300
rect 33818 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34138 11788
rect 33818 10220 34138 11732
rect 38480 36092 38800 36908
rect 38480 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38800 36092
rect 38480 34524 38800 36036
rect 38480 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38800 34524
rect 38480 32956 38800 34468
rect 38480 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38800 32956
rect 38480 31388 38800 32900
rect 38480 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38800 31388
rect 38480 29820 38800 31332
rect 38480 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38800 29820
rect 38480 28252 38800 29764
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26684 38800 28196
rect 38480 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38800 26684
rect 38480 25116 38800 26628
rect 38480 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38800 25116
rect 38480 23548 38800 25060
rect 38480 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38800 23548
rect 38480 21980 38800 23492
rect 38480 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38800 21980
rect 38480 20412 38800 21924
rect 38480 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38800 20412
rect 38480 18844 38800 20356
rect 38480 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38800 18844
rect 38480 17276 38800 18788
rect 38480 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38800 17276
rect 38480 15708 38800 17220
rect 38480 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38800 15708
rect 38480 14140 38800 15652
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 38480 12572 38800 14084
rect 38480 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38800 12572
rect 33818 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34138 10220
rect 33818 8652 34138 10164
rect 35196 11172 35252 11182
rect 33818 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34138 8652
rect 33068 3378 33124 3388
rect 33818 7084 34138 8596
rect 34972 9492 35028 9502
rect 34972 7364 35028 9436
rect 34972 7298 35028 7308
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5516 34138 7028
rect 33818 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34138 5516
rect 33818 3948 34138 5460
rect 33818 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34138 3948
rect 29156 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29476 3164
rect 29156 3076 29476 3108
rect 33818 3076 34138 3892
rect 35196 2100 35252 11116
rect 38480 11004 38800 12516
rect 38480 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38800 11004
rect 38480 9436 38800 10948
rect 38480 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38800 9436
rect 38480 7868 38800 9380
rect 38480 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38800 7868
rect 38480 6300 38800 7812
rect 38480 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38800 6300
rect 38480 4732 38800 6244
rect 38480 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38800 4732
rect 38480 3164 38800 4676
rect 38480 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38800 3164
rect 38480 3076 38800 3108
rect 35196 2034 35252 2044
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31024 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _123_
timestamp 1698431365
transform -1 0 10976 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9632 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _125_
timestamp 1698431365
transform 1 0 9744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _126_
timestamp 1698431365
transform -1 0 8064 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _127_
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _128_
timestamp 1698431365
transform 1 0 1792 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _129_
timestamp 1698431365
transform -1 0 7056 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _130_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _131_
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _132_
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _133_
timestamp 1698431365
transform -1 0 6160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _134_
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _135_
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _136_
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _137_
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _138_
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _139_
timestamp 1698431365
transform -1 0 11200 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _140_
timestamp 1698431365
transform -1 0 10528 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _141_
timestamp 1698431365
transform -1 0 15680 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _142_
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _143_
timestamp 1698431365
transform 1 0 9520 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _144_
timestamp 1698431365
transform -1 0 7728 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _145_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _146_
timestamp 1698431365
transform -1 0 17920 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _147_
timestamp 1698431365
transform -1 0 15344 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _148_
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _149_
timestamp 1698431365
transform 1 0 23072 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _150_
timestamp 1698431365
transform -1 0 22736 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _151_
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _152_
timestamp 1698431365
transform -1 0 18256 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _153_
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _154_
timestamp 1698431365
transform -1 0 20608 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _155_
timestamp 1698431365
transform -1 0 18032 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _156_
timestamp 1698431365
transform -1 0 28336 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _157_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _158_
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _159_
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _160_
timestamp 1698431365
transform -1 0 24752 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _161_
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _162_
timestamp 1698431365
transform -1 0 25760 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _163_
timestamp 1698431365
transform -1 0 24080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _164_
timestamp 1698431365
transform -1 0 22176 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _165_
timestamp 1698431365
transform -1 0 23408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _166_
timestamp 1698431365
transform -1 0 22176 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _167_
timestamp 1698431365
transform -1 0 7728 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _168_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _169_
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _170_
timestamp 1698431365
transform -1 0 6160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _171_
timestamp 1698431365
transform -1 0 6160 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _172_
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _173_
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _174_
timestamp 1698431365
transform 1 0 7392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _175_
timestamp 1698431365
transform 1 0 5600 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _176_
timestamp 1698431365
transform 1 0 1792 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _177_
timestamp 1698431365
transform 1 0 1792 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _178_
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _179_
timestamp 1698431365
transform -1 0 12992 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _180_
timestamp 1698431365
transform -1 0 11312 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _181_
timestamp 1698431365
transform 1 0 13664 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _182_
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _183_
timestamp 1698431365
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _184_
timestamp 1698431365
transform -1 0 14000 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _185_
timestamp 1698431365
transform -1 0 11200 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _186_
timestamp 1698431365
transform -1 0 10640 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _187_
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _188_
timestamp 1698431365
transform -1 0 15120 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _189_
timestamp 1698431365
transform -1 0 22736 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _190_
timestamp 1698431365
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _191_
timestamp 1698431365
transform -1 0 20608 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _192_
timestamp 1698431365
transform 1 0 18704 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _193_
timestamp 1698431365
transform -1 0 18032 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _194_
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _195_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _196_
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _197_
timestamp 1698431365
transform -1 0 17920 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _198_
timestamp 1698431365
transform -1 0 18144 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _199_
timestamp 1698431365
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _200_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _201_
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _202_
timestamp 1698431365
transform -1 0 28560 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _203_
timestamp 1698431365
transform -1 0 27776 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _204_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _205_
timestamp 1698431365
transform -1 0 27888 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _206_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _207_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _208_
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _209_
timestamp 1698431365
transform -1 0 26432 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _210_
timestamp 1698431365
transform -1 0 25760 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _211_
timestamp 1698431365
transform 1 0 30576 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _212_
timestamp 1698431365
transform -1 0 33712 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _213_
timestamp 1698431365
transform 1 0 31584 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _214_
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _215_
timestamp 1698431365
transform -1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _216_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _217_
timestamp 1698431365
transform -1 0 37520 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _218_
timestamp 1698431365
transform -1 0 34496 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _219_
timestamp 1698431365
transform -1 0 32592 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _220_
timestamp 1698431365
transform 1 0 33712 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _221_
timestamp 1698431365
transform -1 0 33600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _222_
timestamp 1698431365
transform 1 0 29456 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _223_
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _224_
timestamp 1698431365
transform -1 0 28784 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _225_
timestamp 1698431365
transform -1 0 33600 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _226_
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _227_
timestamp 1698431365
transform -1 0 37408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _228_
timestamp 1698431365
transform -1 0 33600 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _229_
timestamp 1698431365
transform 1 0 37520 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _230_
timestamp 1698431365
transform 1 0 34832 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _231_
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _232_
timestamp 1698431365
transform -1 0 37520 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _233_
timestamp 1698431365
transform 1 0 31136 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _234_
timestamp 1698431365
transform -1 0 33824 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _235_
timestamp 1698431365
transform -1 0 33600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _236_
timestamp 1698431365
transform -1 0 34720 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _237_
timestamp 1698431365
transform -1 0 34272 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _238_
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _239_
timestamp 1698431365
transform -1 0 37520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _240_
timestamp 1698431365
transform -1 0 37520 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _241_
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _242_
timestamp 1698431365
transform 1 0 37520 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _243_
timestamp 1698431365
transform -1 0 37520 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _244_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _245_
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _246_
timestamp 1698431365
transform -1 0 8512 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _247_
timestamp 1698431365
transform 1 0 3024 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _248_
timestamp 1698431365
transform -1 0 9296 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _249_
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _250_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _251_
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _252_
timestamp 1698431365
transform -1 0 9296 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _253_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _254_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _255_
timestamp 1698431365
transform -1 0 15568 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _256_
timestamp 1698431365
transform 1 0 11088 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _257_
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _258_
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _259_
timestamp 1698431365
transform -1 0 10752 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _260_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _261_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _262_
timestamp 1698431365
transform 1 0 7616 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _263_
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _264_
timestamp 1698431365
transform -1 0 16800 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _265_
timestamp 1698431365
transform 1 0 10976 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _266_
timestamp 1698431365
transform 1 0 19264 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _267_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _268_
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _269_
timestamp 1698431365
transform 1 0 16576 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _270_
timestamp 1698431365
transform 1 0 13216 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _271_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _272_
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _273_
timestamp 1698431365
transform 1 0 13216 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _274_
timestamp 1698431365
transform -1 0 27440 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _275_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _276_
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _277_
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _278_
timestamp 1698431365
transform -1 0 27216 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _279_
timestamp 1698431365
transform 1 0 22176 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _280_
timestamp 1698431365
transform 1 0 20384 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _281_
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _282_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _283_
timestamp 1698431365
transform -1 0 21952 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _284_
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _285_
timestamp 1698431365
transform 1 0 4032 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _286_
timestamp 1698431365
transform 1 0 1904 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _287_
timestamp 1698431365
transform -1 0 5376 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _288_
timestamp 1698431365
transform -1 0 9296 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _289_
timestamp 1698431365
transform 1 0 5264 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _290_
timestamp 1698431365
transform 1 0 4704 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _291_
timestamp 1698431365
transform -1 0 6720 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _292_
timestamp 1698431365
transform -1 0 5376 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _293_
timestamp 1698431365
transform -1 0 5376 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _294_
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _295_
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _296_
timestamp 1698431365
transform 1 0 12320 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _297_
timestamp 1698431365
transform 1 0 11536 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _298_
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _299_
timestamp 1698431365
transform 1 0 8736 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _300_
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _301_
timestamp 1698431365
transform -1 0 9296 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _302_
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _303_
timestamp 1698431365
transform -1 0 12880 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _304_
timestamp 1698431365
transform -1 0 22288 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _305_
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _306_
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _307_
timestamp 1698431365
transform 1 0 14560 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _308_
timestamp 1698431365
transform 1 0 19040 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _309_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _310_
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _311_
timestamp 1698431365
transform -1 0 17136 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _312_
timestamp 1698431365
transform 1 0 13216 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _313_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _314_
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _315_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _316_
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _317_
timestamp 1698431365
transform 1 0 21056 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _318_
timestamp 1698431365
transform -1 0 27216 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _319_
timestamp 1698431365
transform 1 0 21504 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _320_
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _321_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _322_
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _323_
timestamp 1698431365
transform -1 0 24864 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _324_
timestamp 1698431365
transform -1 0 34160 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _325_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _326_
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _327_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _328_
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _329_
timestamp 1698431365
transform 1 0 32816 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _330_
timestamp 1698431365
transform -1 0 36736 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _331_
timestamp 1698431365
transform 1 0 28896 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _332_
timestamp 1698431365
transform 1 0 31024 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _333_
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _334_
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _335_
timestamp 1698431365
transform -1 0 29792 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _336_
timestamp 1698431365
transform -1 0 32816 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _337_
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _338_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _339_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _340_
timestamp 1698431365
transform 1 0 34048 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _341_
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _342_
timestamp 1698431365
transform 1 0 32816 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _343_
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _344_
timestamp 1698431365
transform -1 0 33376 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _345_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _346_
timestamp 1698431365
transform -1 0 34048 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _347_
timestamp 1698431365
transform 1 0 28896 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _348_
timestamp 1698431365
transform 1 0 34160 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _349_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _350_
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _351_
timestamp 1698431365
transform 1 0 32816 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _352_
timestamp 1698431365
transform 1 0 34608 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _353_
timestamp 1698431365
transform -1 0 36736 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32144 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1698431365
transform -1 0 38416 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _382_
timestamp 1698431365
transform 1 0 28224 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _384_
timestamp 1698431365
transform 1 0 21728 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1698431365
transform 1 0 30240 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1698431365
transform 1 0 29568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1698431365
transform 1 0 34160 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _391_
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1698431365
transform 1 0 36064 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _393_
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1698431365
transform -1 0 36064 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _395_
timestamp 1698431365
transform 1 0 28560 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1698431365
transform 1 0 27888 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _400_
timestamp 1698431365
transform -1 0 21056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _402_
timestamp 1698431365
transform 1 0 31472 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _403_
timestamp 1698431365
transform 1 0 26544 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1698431365
transform 1 0 26992 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _406_
timestamp 1698431365
transform 1 0 28112 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1698431365
transform 1 0 21728 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _408_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1698431365
transform 1 0 33488 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1698431365
transform -1 0 30352 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1698431365
transform 1 0 34944 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _412_
timestamp 1698431365
transform 1 0 34272 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1698431365
transform 1 0 34832 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1698431365
transform 1 0 11536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__I
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I
timestamp 1698431365
transform 1 0 30352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698431365
transform 1 0 10640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698431365
transform 1 0 5712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698431365
transform 1 0 11648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698431365
transform 1 0 8624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__CLK
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__CLK
timestamp 1698431365
transform 1 0 15008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__CLK
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__CLK
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__CLK
timestamp 1698431365
transform 1 0 17360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__CLK
timestamp 1698431365
transform 1 0 15904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__CLK
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__CLK
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__CLK
timestamp 1698431365
transform 1 0 16352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__CLK
timestamp 1698431365
transform -1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__CLK
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__CLK
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__CLK
timestamp 1698431365
transform -1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform 1 0 22064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_prog_clk_I
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_prog_clk_I
timestamp 1698431365
transform 1 0 19488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_prog_clk_I
timestamp 1698431365
transform -1 0 15456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_prog_clk_I
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_prog_clk_I
timestamp 1698431365
transform 1 0 22736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_prog_clk_I
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_prog_clk_I
timestamp 1698431365
transform 1 0 25536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_prog_clk_I
timestamp 1698431365
transform -1 0 31472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 37744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 28784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 24304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 35280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 37632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 23632 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 26544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 38416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 37408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 31248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 30912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 26208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 36848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 26208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 38416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 29680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 27216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 29792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 38192 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 18816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 31920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 29344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 20384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 31248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 22960 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 34608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 37296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 29680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 38416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1698431365
transform 1 0 13664 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1698431365
transform 1 0 13888 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1698431365
transform -1 0 31024 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1698431365
transform 1 0 31024 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1698431365
transform -1 0 31024 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1698431365
transform 1 0 31024 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_178 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_210 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_218
timestamp 1698431365
transform 1 0 25760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_251
timestamp 1698431365
transform 1 0 29456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_265
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698431365
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_280
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_297
timestamp 1698431365
transform 1 0 34608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_318
timestamp 1698431365
transform 1 0 36960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 38304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_190
timestamp 1698431365
transform 1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_192
timestamp 1698431365
transform 1 0 22848 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_197
timestamp 1698431365
transform 1 0 23408 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698431365
transform 1 0 24304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_262
timestamp 1698431365
transform 1 0 30688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_266
timestamp 1698431365
transform 1 0 31136 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_292
timestamp 1698431365
transform 1 0 34048 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_306
timestamp 1698431365
transform 1 0 35616 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_209
timestamp 1698431365
transform 1 0 24752 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_251
timestamp 1698431365
transform 1 0 29456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_281
timestamp 1698431365
transform 1 0 32816 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_297
timestamp 1698431365
transform 1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_327
timestamp 1698431365
transform 1 0 37968 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_26
timestamp 1698431365
transform 1 0 4256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_28
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_61
timestamp 1698431365
transform 1 0 8176 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_80
timestamp 1698431365
transform 1 0 10304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_97
timestamp 1698431365
transform 1 0 12208 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_129
timestamp 1698431365
transform 1 0 15792 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_271
timestamp 1698431365
transform 1 0 31696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_288
timestamp 1698431365
transform 1 0 33600 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_299
timestamp 1698431365
transform 1 0 34832 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_41
timestamp 1698431365
transform 1 0 5936 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_58
timestamp 1698431365
transform 1 0 7840 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_74
timestamp 1698431365
transform 1 0 9632 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_98
timestamp 1698431365
transform 1 0 12320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_102
timestamp 1698431365
transform 1 0 12768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_125
timestamp 1698431365
transform 1 0 15344 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_142
timestamp 1698431365
transform 1 0 17248 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_209
timestamp 1698431365
transform 1 0 24752 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_225
timestamp 1698431365
transform 1 0 26544 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_229
timestamp 1698431365
transform 1 0 26992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_269
timestamp 1698431365
transform 1 0 31472 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_273
timestamp 1698431365
transform 1 0 31920 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_306
timestamp 1698431365
transform 1 0 35616 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_327
timestamp 1698431365
transform 1 0 37968 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_36
timestamp 1698431365
transform 1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_40
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_61
timestamp 1698431365
transform 1 0 8176 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_97
timestamp 1698431365
transform 1 0 12208 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_105
timestamp 1698431365
transform 1 0 13104 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_122
timestamp 1698431365
transform 1 0 15008 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_246
timestamp 1698431365
transform 1 0 28896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_250
timestamp 1698431365
transform 1 0 29344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_252
timestamp 1698431365
transform 1 0 29568 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_271
timestamp 1698431365
transform 1 0 31696 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_288
timestamp 1698431365
transform 1 0 33600 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_296
timestamp 1698431365
transform 1 0 34496 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_18
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_55
timestamp 1698431365
transform 1 0 7504 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_87
timestamp 1698431365
transform 1 0 11088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_123
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_127
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_145
timestamp 1698431365
transform 1 0 17584 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_153
timestamp 1698431365
transform 1 0 18480 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_170
timestamp 1698431365
transform 1 0 20384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_188
timestamp 1698431365
transform 1 0 22400 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_236
timestamp 1698431365
transform 1 0 27776 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_251
timestamp 1698431365
transform 1 0 29456 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_258
timestamp 1698431365
transform 1 0 30240 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_262
timestamp 1698431365
transform 1 0 30688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_264
timestamp 1698431365
transform 1 0 30912 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_283
timestamp 1698431365
transform 1 0 33040 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_291
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_293
timestamp 1698431365
transform 1 0 34160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_327
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_10
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_14
timestamp 1698431365
transform 1 0 2912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_49
timestamp 1698431365
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_53
timestamp 1698431365
transform 1 0 7280 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_84
timestamp 1698431365
transform 1 0 10752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_120
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_124
timestamp 1698431365
transform 1 0 15232 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_167
timestamp 1698431365
transform 1 0 20048 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_199
timestamp 1698431365
transform 1 0 23632 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_244
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_261
timestamp 1698431365
transform 1 0 30576 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_327
timestamp 1698431365
transform 1 0 37968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_6
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_23
timestamp 1698431365
transform 1 0 3920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_71
timestamp 1698431365
transform 1 0 9296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_73
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_80
timestamp 1698431365
transform 1 0 10304 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_88
timestamp 1698431365
transform 1 0 11200 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_141
timestamp 1698431365
transform 1 0 17136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_145
timestamp 1698431365
transform 1 0 17584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_149
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_157
timestamp 1698431365
transform 1 0 18928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_202
timestamp 1698431365
transform 1 0 23968 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_218
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_236
timestamp 1698431365
transform 1 0 27776 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_279
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_283
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_287
timestamp 1698431365
transform 1 0 33488 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_327
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_4
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_21
timestamp 1698431365
transform 1 0 3696 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_29
timestamp 1698431365
transform 1 0 4592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_64
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_95
timestamp 1698431365
transform 1 0 11984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_99
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_103
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_148
timestamp 1698431365
transform 1 0 17920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_152
timestamp 1698431365
transform 1 0 18368 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_156
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_174
timestamp 1698431365
transform 1 0 20832 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_182
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_199
timestamp 1698431365
transform 1 0 23632 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_237
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_245
timestamp 1698431365
transform 1 0 28784 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_262
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_316
timestamp 1698431365
transform 1 0 36736 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_327
timestamp 1698431365
transform 1 0 37968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_49
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_94
timestamp 1698431365
transform 1 0 11872 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_127
timestamp 1698431365
transform 1 0 15568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_129
timestamp 1698431365
transform 1 0 15792 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_132
timestamp 1698431365
transform 1 0 16128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_202
timestamp 1698431365
transform 1 0 23968 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_210
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_227
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_257
timestamp 1698431365
transform 1 0 30128 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_298
timestamp 1698431365
transform 1 0 34720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_300
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_74
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_81
timestamp 1698431365
transform 1 0 10416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_85
timestamp 1698431365
transform 1 0 10864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_87
timestamp 1698431365
transform 1 0 11088 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_151
timestamp 1698431365
transform 1 0 18256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_153
timestamp 1698431365
transform 1 0 18480 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_200
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_202
timestamp 1698431365
transform 1 0 23968 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_222
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_247
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_255
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_10
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_51
timestamp 1698431365
transform 1 0 7056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_55
timestamp 1698431365
transform 1 0 7504 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_90
timestamp 1698431365
transform 1 0 11424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_251
timestamp 1698431365
transform 1 0 29456 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_286
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_294
timestamp 1698431365
transform 1 0 34272 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_296
timestamp 1698431365
transform 1 0 34496 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_43
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_62
timestamp 1698431365
transform 1 0 8288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_64
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_67
timestamp 1698431365
transform 1 0 8848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_109
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_160
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_164
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_168
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_323
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_128
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_135
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_149
timestamp 1698431365
transform 1 0 18032 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_184
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_188
timestamp 1698431365
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_190
timestamp 1698431365
transform 1 0 22624 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_265
timestamp 1698431365
transform 1 0 31024 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_316
timestamp 1698431365
transform 1 0 36736 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_324
timestamp 1698431365
transform 1 0 37632 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_328
timestamp 1698431365
transform 1 0 38080 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_43
timestamp 1698431365
transform 1 0 6160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_47
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_186
timestamp 1698431365
transform 1 0 22176 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_194
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_196
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_4
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_61
timestamp 1698431365
transform 1 0 8176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_63
timestamp 1698431365
transform 1 0 8400 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_86
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_121
timestamp 1698431365
transform 1 0 14896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_123
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_161
timestamp 1698431365
transform 1 0 19376 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_169
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_218
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_254
timestamp 1698431365
transform 1 0 29792 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_258
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_326
timestamp 1698431365
transform 1 0 37856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_330
timestamp 1698431365
transform 1 0 38304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_6
timestamp 1698431365
transform 1 0 2016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_179
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_26
timestamp 1698431365
transform 1 0 4256 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_90
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_133
timestamp 1698431365
transform 1 0 16240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_156
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_256
timestamp 1698431365
transform 1 0 30016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_258
timestamp 1698431365
transform 1 0 30240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_275
timestamp 1698431365
transform 1 0 32144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_328
timestamp 1698431365
transform 1 0 38080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_47
timestamp 1698431365
transform 1 0 6608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_49
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_84
timestamp 1698431365
transform 1 0 10752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_141
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_148
timestamp 1698431365
transform 1 0 17920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_156
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_158
timestamp 1698431365
transform 1 0 19040 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_64
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_97
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_105
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_176
timestamp 1698431365
transform 1 0 21056 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_183
timestamp 1698431365
transform 1 0 21840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_187
timestamp 1698431365
transform 1 0 22288 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_191
timestamp 1698431365
transform 1 0 22736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_193
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_258
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_324
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_127
timestamp 1698431365
transform 1 0 15568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_163
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_191
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_195
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_237
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_305
timestamp 1698431365
transform 1 0 35504 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_86
timestamp 1698431365
transform 1 0 10976 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_192
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_200
timestamp 1698431365
transform 1 0 23744 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_288
timestamp 1698431365
transform 1 0 33600 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_295
timestamp 1698431365
transform 1 0 34384 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_162
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_166
timestamp 1698431365
transform 1 0 19936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_218
timestamp 1698431365
transform 1 0 25760 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_222
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_261
timestamp 1698431365
transform 1 0 30576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_122
timestamp 1698431365
transform 1 0 15008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_126
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_156
timestamp 1698431365
transform 1 0 18816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_214
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_265
timestamp 1698431365
transform 1 0 31024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_269
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_316
timestamp 1698431365
transform 1 0 36736 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_324
timestamp 1698431365
transform 1 0 37632 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_328
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_60
timestamp 1698431365
transform 1 0 8064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_68
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_129
timestamp 1698431365
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_165
timestamp 1698431365
transform 1 0 19824 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_191
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_236
timestamp 1698431365
transform 1 0 27776 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_272
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_280
timestamp 1698431365
transform 1 0 32704 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_297
timestamp 1698431365
transform 1 0 34608 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_323
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_4
timestamp 1698431365
transform 1 0 1792 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_21
timestamp 1698431365
transform 1 0 3696 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_29
timestamp 1698431365
transform 1 0 4592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_64
timestamp 1698431365
transform 1 0 8512 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_123
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_149
timestamp 1698431365
transform 1 0 18032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_187
timestamp 1698431365
transform 1 0 22288 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_264
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_268
timestamp 1698431365
transform 1 0 31360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_289
timestamp 1698431365
transform 1 0 33712 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_330
timestamp 1698431365
transform 1 0 38304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_4
timestamp 1698431365
transform 1 0 1792 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_21
timestamp 1698431365
transform 1 0 3696 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_29
timestamp 1698431365
transform 1 0 4592 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_33
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_132
timestamp 1698431365
transform 1 0 16128 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_140
timestamp 1698431365
transform 1 0 17024 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_203
timestamp 1698431365
transform 1 0 24080 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_211
timestamp 1698431365
transform 1 0 24976 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_237
timestamp 1698431365
transform 1 0 27888 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_323
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_327
timestamp 1698431365
transform 1 0 37968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_89
timestamp 1698431365
transform 1 0 11312 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_97
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_316
timestamp 1698431365
transform 1 0 36736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_320
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_49
timestamp 1698431365
transform 1 0 6832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_100
timestamp 1698431365
transform 1 0 12544 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_117
timestamp 1698431365
transform 1 0 14448 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_152
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_154
timestamp 1698431365
transform 1 0 18592 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_161
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_221
timestamp 1698431365
transform 1 0 26096 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_253
timestamp 1698431365
transform 1 0 29680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_257
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_293
timestamp 1698431365
transform 1 0 34160 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_309
timestamp 1698431365
transform 1 0 35952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_327
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_34
timestamp 1698431365
transform 1 0 5152 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_42
timestamp 1698431365
transform 1 0 6048 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_46
timestamp 1698431365
transform 1 0 6496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_48
timestamp 1698431365
transform 1 0 6720 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_65
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_88
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_90
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_137
timestamp 1698431365
transform 1 0 16688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_152
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_169
timestamp 1698431365
transform 1 0 20272 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_258
timestamp 1698431365
transform 1 0 30240 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_270
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_272
timestamp 1698431365
transform 1 0 31808 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_307
timestamp 1698431365
transform 1 0 35728 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_69
timestamp 1698431365
transform 1 0 9072 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_89
timestamp 1698431365
transform 1 0 11312 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_139
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_147
timestamp 1698431365
transform 1 0 17808 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_209
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_225
timestamp 1698431365
transform 1 0 26544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_227
timestamp 1698431365
transform 1 0 26768 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_272
timestamp 1698431365
transform 1 0 31808 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_280
timestamp 1698431365
transform 1 0 32704 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_297
timestamp 1698431365
transform 1 0 34608 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_113
timestamp 1698431365
transform 1 0 14000 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_121
timestamp 1698431365
transform 1 0 14896 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_228
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_257
timestamp 1698431365
transform 1 0 30128 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_273
timestamp 1698431365
transform 1 0 31920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_277
timestamp 1698431365
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_307
timestamp 1698431365
transform 1 0 35728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_317
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_77
timestamp 1698431365
transform 1 0 9968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_79
timestamp 1698431365
transform 1 0 10192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_96
timestamp 1698431365
transform 1 0 12096 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_132
timestamp 1698431365
transform 1 0 16128 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_164
timestamp 1698431365
transform 1 0 19712 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_263
timestamp 1698431365
transform 1 0 30800 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_296
timestamp 1698431365
transform 1 0 34496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_298
timestamp 1698431365
transform 1 0 34720 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_310
timestamp 1698431365
transform 1 0 36064 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_279
timestamp 1698431365
transform 1 0 32592 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_287
timestamp 1698431365
transform 1 0 33488 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_291
timestamp 1698431365
transform 1 0 33936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_322
timestamp 1698431365
transform 1 0 37408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_326
timestamp 1698431365
transform 1 0 37856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_328
timestamp 1698431365
transform 1 0 38080 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_279
timestamp 1698431365
transform 1 0 32592 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_287
timestamp 1698431365
transform 1 0 33488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_289
timestamp 1698431365
transform 1 0 33712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_306
timestamp 1698431365
transform 1 0 35616 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_327
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_322
timestamp 1698431365
transform 1 0 37408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_330
timestamp 1698431365
transform 1 0 38304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_139
timestamp 1698431365
transform 1 0 16912 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_155
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_163
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_167
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_169
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_172
timestamp 1698431365
transform 1 0 20608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_189
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_193
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_199
timestamp 1698431365
transform 1 0 23632 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_211
timestamp 1698431365
transform 1 0 24976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_271
timestamp 1698431365
transform 1 0 31696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_281
timestamp 1698431365
transform 1 0 32816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_327
timestamp 1698431365
transform 1 0 37968 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_152
timestamp 1698431365
transform 1 0 18368 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_162
timestamp 1698431365
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_192
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_241
timestamp 1698431365
transform 1 0 28336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_251
timestamp 1698431365
transform 1 0 29456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_257
timestamp 1698431365
transform 1 0 30128 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_264
timestamp 1698431365
transform 1 0 30912 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_268
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_293
timestamp 1698431365
transform 1 0 34160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_327
timestamp 1698431365
transform 1 0 37968 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_36
timestamp 1698431365
transform 1 0 5376 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_138
timestamp 1698431365
transform 1 0 16800 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_142
timestamp 1698431365
transform 1 0 17248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_199
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_203
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_206
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_214
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_235
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_237
timestamp 1698431365
transform 1 0 27888 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_250
timestamp 1698431365
transform 1 0 29344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_258
timestamp 1698431365
transform 1 0 30240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_265
timestamp 1698431365
transform 1 0 31024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_267
timestamp 1698431365
transform 1 0 31248 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_284
timestamp 1698431365
transform 1 0 33152 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_298
timestamp 1698431365
transform 1 0 34720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_316
timestamp 1698431365
transform 1 0 36736 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_327
timestamp 1698431365
transform 1 0 37968 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35392 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 36400 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 20384 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 32592 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 20832 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform 1 0 17584 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 34608 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform 1 0 9520 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 32704 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform 1 0 6272 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 16128 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 32592 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform 1 0 6384 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 23968 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 24080 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 23968 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform -1 0 12320 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 26768 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 8736 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 20944 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 13216 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 15008 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform -1 0 24752 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 16912 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 38416 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform -1 0 30128 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 11312 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform 1 0 29904 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 28672 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 12096 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform 1 0 15344 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 12208 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 36064 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 8624 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 36064 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform -1 0 28112 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform -1 0 12208 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 19712 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 27216 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform -1 0 27888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform -1 0 37408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold50
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform -1 0 30688 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform -1 0 32144 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 32592 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform 1 0 10416 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 6384 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform -1 0 35952 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform 1 0 2128 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform -1 0 36176 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform -1 0 21056 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform -1 0 29008 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 20048 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform 1 0 10192 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform -1 0 37408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform -1 0 23632 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform 1 0 22064 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold69
timestamp 1698431365
transform 1 0 31024 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold70
timestamp 1698431365
transform -1 0 35728 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold71
timestamp 1698431365
transform 1 0 6048 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold72
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold73
timestamp 1698431365
transform 1 0 32816 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold74
timestamp 1698431365
transform 1 0 6496 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold75
timestamp 1698431365
transform -1 0 30576 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold76
timestamp 1698431365
transform 1 0 15456 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold77
timestamp 1698431365
transform 1 0 25984 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold78
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold79
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold80
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold81
timestamp 1698431365
transform -1 0 31808 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold82
timestamp 1698431365
transform 1 0 33824 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold83
timestamp 1698431365
transform -1 0 21056 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold84
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold85
timestamp 1698431365
transform -1 0 31808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold86
timestamp 1698431365
transform 1 0 1904 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold87
timestamp 1698431365
transform -1 0 16912 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold88
timestamp 1698431365
transform -1 0 17584 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold89
timestamp 1698431365
transform -1 0 33824 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold90
timestamp 1698431365
transform -1 0 35616 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold91
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold92
timestamp 1698431365
transform -1 0 14000 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold93
timestamp 1698431365
transform -1 0 38416 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold94
timestamp 1698431365
transform 1 0 29904 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold95
timestamp 1698431365
transform 1 0 14336 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold96
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold97
timestamp 1698431365
transform -1 0 20272 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold98
timestamp 1698431365
transform 1 0 1904 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold99
timestamp 1698431365
transform -1 0 34608 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold100
timestamp 1698431365
transform -1 0 35728 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold101
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold102
timestamp 1698431365
transform 1 0 1904 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold103
timestamp 1698431365
transform -1 0 13216 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold104
timestamp 1698431365
transform 1 0 6384 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold105
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold106
timestamp 1698431365
transform 1 0 6384 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold107
timestamp 1698431365
transform -1 0 33040 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold108
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold109
timestamp 1698431365
transform -1 0 5264 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 38416 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 29456 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 24304 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 35952 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 37744 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 23632 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 17472 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 27216 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 38416 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 38416 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 38080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 30688 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 31360 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 29568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 27328 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 38416 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 26880 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 28560 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 26544 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 31024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 38416 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 18144 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 29904 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 27440 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 19712 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 31024 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 35280 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 38416 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 27552 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34496 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output39
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output40
timestamp 1698431365
transform -1 0 36624 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41
timestamp 1698431365
transform 1 0 33040 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 33712 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output49 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22512 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output50
timestamp 1698431365
transform 1 0 28336 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output51
timestamp 1698431365
transform -1 0 31024 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698431365
transform 1 0 22512 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform 1 0 29904 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output55
timestamp 1698431365
transform 1 0 25424 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output56
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output57
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform 1 0 27216 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output60
timestamp 1698431365
transform 1 0 36848 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698431365
transform 1 0 33600 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output62
timestamp 1698431365
transform -1 0 27216 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output63
timestamp 1698431365
transform -1 0 20384 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output64
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output65
timestamp 1698431365
transform 1 0 35280 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform 1 0 36848 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 29568 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output69
timestamp 1698431365
transform 1 0 36848 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output70
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output71
timestamp 1698431365
transform 1 0 22288 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__73
timestamp 1698431365
transform -1 0 23408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__74
timestamp 1698431365
transform 1 0 37296 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__75
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__76
timestamp 1698431365
transform -1 0 24864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__77
timestamp 1698431365
transform -1 0 22848 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__78
timestamp 1698431365
transform -1 0 30128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__79
timestamp 1698431365
transform 1 0 36400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__80
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__81
timestamp 1698431365
transform 1 0 35168 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__82
timestamp 1698431365
transform -1 0 30240 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__83
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__84
timestamp 1698431365
transform 1 0 36064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__85
timestamp 1698431365
transform 1 0 33376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__86
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__87
timestamp 1698431365
transform 1 0 33264 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__88
timestamp 1698431365
transform -1 0 35616 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__89
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__90
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__91
timestamp 1698431365
transform 1 0 36624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__92
timestamp 1698431365
transform 1 0 33712 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__93
timestamp 1698431365
transform 1 0 26208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__94
timestamp 1698431365
transform 1 0 33040 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__95
timestamp 1698431365
transform 1 0 31360 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__96
timestamp 1698431365
transform 1 0 34720 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_2__1__97
timestamp 1698431365
transform -1 0 26992 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_95
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_96
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_97
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_98
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_99
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_100
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_101
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_102
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_103
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_104
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_105
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_106
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_107
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_108
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_109
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_110
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_111
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_112
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_113
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_114
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_115
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_116
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_117
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_118
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_119
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_120
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_121
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_123
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_124
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_125
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_126
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_130
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_132
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_135
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_136
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_137
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_140
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_141
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_142
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_143
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_144
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_145
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_146
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_147
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_148
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_152
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_158
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_159
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_162
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_163
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_164
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_165
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_166
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_167
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_168
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_169
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_170
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_171
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_172
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_173
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_174
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_175
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_176
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_177
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_178
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_179
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_180
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_181
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_182
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_183
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_184
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_185
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_186
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_187
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_188
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_189
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_190
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_191
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_192
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_193
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_194
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_195
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_196
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_197
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_198
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_199
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_200
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_201
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_202
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_203
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_204
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_205
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_206
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_207
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_208
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_209
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_210
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_211
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_212
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_213
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_214
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_215
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_216
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_217
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_218
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_219
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_220
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_221
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_222
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_223
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_224
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_225
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_226
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_227
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_228
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_229
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_230
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_231
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_232
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_233
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_234
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_235
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_236
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_237
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_238
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_239
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_240
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_241
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_242
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_243
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_244
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_245
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_246
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_247
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_248
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_249
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_250
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_252
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_253
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_260
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_263
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_264
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_265
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_266
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_267
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_268
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_269
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_270
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_271
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_272
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_273
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_274
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_275
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_276
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_277
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_278
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_279
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_280
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_281
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_282
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_283
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
<< labels >>
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 2 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 3 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 ccff_head
port 6 nsew signal input
flabel metal3 s 39200 16800 40000 16912 0 FreeSans 448 0 0 0 ccff_tail
port 7 nsew signal tristate
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 chanx_left_in[0]
port 8 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 chanx_left_in[10]
port 9 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 chanx_left_in[11]
port 10 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 chanx_left_in[12]
port 11 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chanx_left_in[13]
port 12 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chanx_left_in[14]
port 13 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chanx_left_in[15]
port 14 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 chanx_left_in[16]
port 15 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chanx_left_in[17]
port 16 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chanx_left_in[18]
port 17 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 chanx_left_in[19]
port 18 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chanx_left_in[1]
port 19 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chanx_left_in[2]
port 20 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chanx_left_in[3]
port 21 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 chanx_left_in[4]
port 22 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chanx_left_in[5]
port 23 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chanx_left_in[6]
port 24 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chanx_left_in[7]
port 25 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chanx_left_in[8]
port 26 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chanx_left_in[9]
port 27 nsew signal input
flabel metal2 s 26208 39200 26320 40000 0 FreeSans 448 90 0 0 chanx_left_out[0]
port 28 nsew signal tristate
flabel metal2 s 37632 39200 37744 40000 0 FreeSans 448 90 0 0 chanx_left_out[10]
port 29 nsew signal tristate
flabel metal2 s 36288 39200 36400 40000 0 FreeSans 448 90 0 0 chanx_left_out[11]
port 30 nsew signal tristate
flabel metal2 s 34944 39200 35056 40000 0 FreeSans 448 90 0 0 chanx_left_out[12]
port 31 nsew signal tristate
flabel metal3 s 39200 0 40000 112 0 FreeSans 448 0 0 0 chanx_left_out[13]
port 32 nsew signal tristate
flabel metal3 s 39200 25536 40000 25648 0 FreeSans 448 0 0 0 chanx_left_out[14]
port 33 nsew signal tristate
flabel metal2 s 28896 39200 29008 40000 0 FreeSans 448 90 0 0 chanx_left_out[15]
port 34 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 chanx_left_out[16]
port 35 nsew signal tristate
flabel metal3 s 39200 11424 40000 11536 0 FreeSans 448 0 0 0 chanx_left_out[17]
port 36 nsew signal tristate
flabel metal3 s 39200 39648 40000 39760 0 FreeSans 448 0 0 0 chanx_left_out[18]
port 37 nsew signal tristate
flabel metal2 s 32928 39200 33040 40000 0 FreeSans 448 90 0 0 chanx_left_out[19]
port 38 nsew signal tristate
flabel metal3 s 39200 33600 40000 33712 0 FreeSans 448 0 0 0 chanx_left_out[1]
port 39 nsew signal tristate
flabel metal2 s 31584 39200 31696 40000 0 FreeSans 448 90 0 0 chanx_left_out[2]
port 40 nsew signal tristate
flabel metal3 s 39200 4032 40000 4144 0 FreeSans 448 0 0 0 chanx_left_out[3]
port 41 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 chanx_left_out[4]
port 42 nsew signal tristate
flabel metal2 s 34272 39200 34384 40000 0 FreeSans 448 90 0 0 chanx_left_out[5]
port 43 nsew signal tristate
flabel metal3 s 39200 32928 40000 33040 0 FreeSans 448 0 0 0 chanx_left_out[6]
port 44 nsew signal tristate
flabel metal3 s 39200 3360 40000 3472 0 FreeSans 448 0 0 0 chanx_left_out[7]
port 45 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 chanx_left_out[8]
port 46 nsew signal tristate
flabel metal2 s 33600 39200 33712 40000 0 FreeSans 448 90 0 0 chanx_left_out[9]
port 47 nsew signal tristate
flabel metal3 s 39200 27552 40000 27664 0 FreeSans 448 0 0 0 chany_bottom_in[0]
port 48 nsew signal input
flabel metal2 s 28224 39200 28336 40000 0 FreeSans 448 90 0 0 chany_bottom_in[10]
port 49 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 chany_bottom_in[11]
port 50 nsew signal input
flabel metal2 s 24192 39200 24304 40000 0 FreeSans 448 90 0 0 chany_bottom_in[12]
port 51 nsew signal input
flabel metal3 s 39200 2016 40000 2128 0 FreeSans 448 0 0 0 chany_bottom_in[13]
port 52 nsew signal input
flabel metal2 s 36960 39200 37072 40000 0 FreeSans 448 90 0 0 chany_bottom_in[14]
port 53 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chany_bottom_in[15]
port 54 nsew signal input
flabel metal2 s 23520 39200 23632 40000 0 FreeSans 448 90 0 0 chany_bottom_in[16]
port 55 nsew signal input
flabel metal2 s 18144 39200 18256 40000 0 FreeSans 448 90 0 0 chany_bottom_in[17]
port 56 nsew signal input
flabel metal3 s 39200 5376 40000 5488 0 FreeSans 448 0 0 0 chany_bottom_in[18]
port 57 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 chany_bottom_in[19]
port 58 nsew signal input
flabel metal3 s 39200 26880 40000 26992 0 FreeSans 448 0 0 0 chany_bottom_in[1]
port 59 nsew signal input
flabel metal3 s 39200 28224 40000 28336 0 FreeSans 448 0 0 0 chany_bottom_in[2]
port 60 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chany_bottom_in[3]
port 61 nsew signal input
flabel metal3 s 39200 1344 40000 1456 0 FreeSans 448 0 0 0 chany_bottom_in[4]
port 62 nsew signal input
flabel metal3 s 39200 8736 40000 8848 0 FreeSans 448 0 0 0 chany_bottom_in[5]
port 63 nsew signal input
flabel metal3 s 39200 672 40000 784 0 FreeSans 448 0 0 0 chany_bottom_in[6]
port 64 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 chany_bottom_in[7]
port 65 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 chany_bottom_in[8]
port 66 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 chany_bottom_in[9]
port 67 nsew signal input
flabel metal3 s 39200 34272 40000 34384 0 FreeSans 448 0 0 0 chany_bottom_out[0]
port 68 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 chany_bottom_out[10]
port 69 nsew signal tristate
flabel metal3 s 39200 26208 40000 26320 0 FreeSans 448 0 0 0 chany_bottom_out[11]
port 70 nsew signal tristate
flabel metal2 s 29568 39200 29680 40000 0 FreeSans 448 90 0 0 chany_bottom_out[12]
port 71 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 chany_bottom_out[13]
port 72 nsew signal tristate
flabel metal3 s 39200 9408 40000 9520 0 FreeSans 448 0 0 0 chany_bottom_out[14]
port 73 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 chany_bottom_out[15]
port 74 nsew signal tristate
flabel metal2 s 21504 39200 21616 40000 0 FreeSans 448 90 0 0 chany_bottom_out[16]
port 75 nsew signal tristate
flabel metal2 s 30912 39200 31024 40000 0 FreeSans 448 90 0 0 chany_bottom_out[17]
port 76 nsew signal tristate
flabel metal3 s 39200 38304 40000 38416 0 FreeSans 448 0 0 0 chany_bottom_out[18]
port 77 nsew signal tristate
flabel metal2 s 20832 39200 20944 40000 0 FreeSans 448 90 0 0 chany_bottom_out[19]
port 78 nsew signal tristate
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal2 s 22176 39200 22288 40000 0 FreeSans 448 90 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal3 s 39200 32256 40000 32368 0 FreeSans 448 0 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal2 s 24864 39200 24976 40000 0 FreeSans 448 90 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 39200 2688 40000 2800 0 FreeSans 448 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal3 s 39200 36960 40000 37072 0 FreeSans 448 0 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal3 s 39200 29568 40000 29680 0 FreeSans 448 0 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal3 s 39200 37632 40000 37744 0 FreeSans 448 0 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal3 s 39200 10752 40000 10864 0 FreeSans 448 0 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal3 s 39200 6720 40000 6832 0 FreeSans 448 0 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal2 s 30240 39200 30352 40000 0 FreeSans 448 90 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal3 s 39200 35616 40000 35728 0 FreeSans 448 0 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 18816 39200 18928 40000 0 FreeSans 448 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 chany_top_in[19]
port 98 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 chany_top_in[1]
port 99 nsew signal input
flabel metal2 s 20160 39200 20272 40000 0 FreeSans 448 90 0 0 chany_top_in[2]
port 100 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 chany_top_in[3]
port 101 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 chany_top_in[4]
port 102 nsew signal input
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 chany_top_in[5]
port 103 nsew signal input
flabel metal2 s 22848 39200 22960 40000 0 FreeSans 448 90 0 0 chany_top_in[6]
port 104 nsew signal input
flabel metal2 s 35616 39200 35728 40000 0 FreeSans 448 90 0 0 chany_top_in[7]
port 105 nsew signal input
flabel metal3 s 39200 28896 40000 29008 0 FreeSans 448 0 0 0 chany_top_in[8]
port 106 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 chany_top_in[9]
port 107 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 chany_top_out[0]
port 108 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 chany_top_out[10]
port 109 nsew signal tristate
flabel metal2 s 27552 39200 27664 40000 0 FreeSans 448 90 0 0 chany_top_out[11]
port 110 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 chany_top_out[12]
port 111 nsew signal tristate
flabel metal2 s 26880 39200 26992 40000 0 FreeSans 448 90 0 0 chany_top_out[13]
port 112 nsew signal tristate
flabel metal3 s 39200 8064 40000 8176 0 FreeSans 448 0 0 0 chany_top_out[14]
port 113 nsew signal tristate
flabel metal2 s 32256 39200 32368 40000 0 FreeSans 448 90 0 0 chany_top_out[15]
port 114 nsew signal tristate
flabel metal3 s 39200 31584 40000 31696 0 FreeSans 448 0 0 0 chany_top_out[16]
port 115 nsew signal tristate
flabel metal2 s 25536 39200 25648 40000 0 FreeSans 448 90 0 0 chany_top_out[17]
port 116 nsew signal tristate
flabel metal2 s 19488 39200 19600 40000 0 FreeSans 448 90 0 0 chany_top_out[18]
port 117 nsew signal tristate
flabel metal3 s 39200 10080 40000 10192 0 FreeSans 448 0 0 0 chany_top_out[19]
port 118 nsew signal tristate
flabel metal3 s 39200 36288 40000 36400 0 FreeSans 448 0 0 0 chany_top_out[1]
port 119 nsew signal tristate
flabel metal3 s 39200 34944 40000 35056 0 FreeSans 448 0 0 0 chany_top_out[2]
port 120 nsew signal tristate
flabel metal3 s 39200 38976 40000 39088 0 FreeSans 448 0 0 0 chany_top_out[3]
port 121 nsew signal tristate
flabel metal3 s 39200 30240 40000 30352 0 FreeSans 448 0 0 0 chany_top_out[4]
port 122 nsew signal tristate
flabel metal3 s 39200 4704 40000 4816 0 FreeSans 448 0 0 0 chany_top_out[5]
port 123 nsew signal tristate
flabel metal3 s 39200 6048 40000 6160 0 FreeSans 448 0 0 0 chany_top_out[6]
port 124 nsew signal tristate
flabel metal3 s 39200 7392 40000 7504 0 FreeSans 448 0 0 0 chany_top_out[7]
port 125 nsew signal tristate
flabel metal3 s 39200 30912 40000 31024 0 FreeSans 448 0 0 0 chany_top_out[8]
port 126 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 chany_top_out[9]
port 127 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 128 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 129 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 130 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 131 nsew signal input
flabel metal3 s 39200 16128 40000 16240 0 FreeSans 448 0 0 0 pReset
port 132 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 prog_clk
port 133 nsew signal input
flabel metal3 s 39200 14784 40000 14896 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 134 nsew signal input
flabel metal3 s 39200 15456 40000 15568 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 135 nsew signal input
flabel metal3 s 39200 12768 40000 12880 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 136 nsew signal input
flabel metal3 s 39200 12096 40000 12208 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 137 nsew signal input
flabel metal3 s 39200 13440 40000 13552 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 138 nsew signal input
flabel metal3 s 39200 14112 40000 14224 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 139 nsew signal input
flabel metal4 s 5846 3076 6166 36908 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 15170 3076 15490 36908 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 24494 3076 24814 36908 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 33818 3076 34138 36908 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 10508 3076 10828 36908 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
flabel metal4 s 19832 3076 20152 36908 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
flabel metal4 s 29156 3076 29476 36908 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
flabel metal4 s 38480 3076 38800 36908 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
rlabel metal1 19992 36848 19992 36848 0 vdd
rlabel via1 20072 36064 20072 36064 0 vss
rlabel metal2 10024 10528 10024 10528 0 _000_
rlabel metal2 10136 12152 10136 12152 0 _001_
rlabel metal2 5544 11032 5544 11032 0 _002_
rlabel metal2 6216 9632 6216 9632 0 _003_
rlabel metal2 2296 11984 2296 11984 0 _004_
rlabel metal2 4760 8848 4760 8848 0 _005_
rlabel metal2 5880 15512 5880 15512 0 _006_
rlabel metal2 2072 13776 2072 13776 0 _007_
rlabel metal2 6216 17192 6216 17192 0 _008_
rlabel metal3 5208 15960 5208 15960 0 _009_
rlabel metal2 16296 17920 16296 17920 0 _010_
rlabel metal2 12376 18872 12376 18872 0 _011_
rlabel metal3 13104 17080 13104 17080 0 _012_
rlabel metal2 12488 15232 12488 15232 0 _013_
rlabel metal2 10920 17080 10920 17080 0 _014_
rlabel metal2 7784 18704 7784 18704 0 _015_
rlabel metal3 12656 15176 12656 15176 0 _016_
rlabel metal2 12376 12656 12376 12656 0 _017_
rlabel metal2 9800 11760 9800 11760 0 _018_
rlabel metal2 7560 15848 7560 15848 0 _019_
rlabel metal3 15624 10696 15624 10696 0 _020_
rlabel metal2 14168 9464 14168 9464 0 _021_
rlabel metal2 22232 12600 22232 12600 0 _022_
rlabel metal2 23464 12656 23464 12656 0 _023_
rlabel metal3 21196 13048 21196 13048 0 _024_
rlabel metal2 19544 11424 19544 11424 0 _025_
rlabel metal2 16408 12320 16408 12320 0 _026_
rlabel metal2 16296 14000 16296 14000 0 _027_
rlabel metal2 19320 15904 19320 15904 0 _028_
rlabel metal2 16408 14560 16408 14560 0 _029_
rlabel metal2 24360 15512 24360 15512 0 _030_
rlabel metal2 28056 14168 28056 14168 0 _031_
rlabel metal2 26040 12488 26040 12488 0 _032_
rlabel metal2 24248 13104 24248 13104 0 _033_
rlabel metal3 25984 15848 25984 15848 0 _034_
rlabel metal2 25256 17192 25256 17192 0 _035_
rlabel metal2 23576 17696 23576 17696 0 _036_
rlabel metal2 21784 18144 21784 18144 0 _037_
rlabel metal2 22904 18088 22904 18088 0 _038_
rlabel metal2 18984 15848 18984 15848 0 _039_
rlabel metal3 9128 21784 9128 21784 0 _040_
rlabel metal2 7112 21616 7112 21616 0 _041_
rlabel metal2 4984 18592 4984 18592 0 _042_
rlabel metal2 2408 17248 2408 17248 0 _043_
rlabel metal3 5040 21448 5040 21448 0 _044_
rlabel metal2 8344 19264 8344 19264 0 _045_
rlabel metal2 7896 24080 7896 24080 0 _046_
rlabel metal2 3752 23520 3752 23520 0 _047_
rlabel metal2 2352 24024 2352 24024 0 _048_
rlabel metal2 2296 22008 2296 22008 0 _049_
rlabel metal3 11312 21112 11312 21112 0 _050_
rlabel metal2 10920 22568 10920 22568 0 _051_
rlabel metal2 14168 25984 14168 25984 0 _052_
rlabel metal3 15568 26488 15568 26488 0 _053_
rlabel metal3 12992 24024 12992 24024 0 _054_
rlabel metal3 12600 26936 12600 26936 0 _055_
rlabel metal2 8344 27104 8344 27104 0 _056_
rlabel metal2 10136 25088 10136 25088 0 _057_
rlabel metal2 14280 22848 14280 22848 0 _058_
rlabel metal2 14616 21504 14616 21504 0 _059_
rlabel metal2 21336 24416 21336 24416 0 _060_
rlabel metal2 20216 24640 20216 24640 0 _061_
rlabel metal2 18984 25312 18984 25312 0 _062_
rlabel metal2 17528 25816 17528 25816 0 _063_
rlabel metal2 21840 21672 21840 21672 0 _064_
rlabel metal2 20440 21224 20440 21224 0 _065_
rlabel metal2 18760 21056 18760 21056 0 _066_
rlabel metal2 17416 19040 17416 19040 0 _067_
rlabel metal3 17024 20216 17024 20216 0 _068_
rlabel metal2 14056 22400 14056 22400 0 _069_
rlabel metal3 30072 24920 30072 24920 0 _070_
rlabel metal2 28280 22736 28280 22736 0 _071_
rlabel metal2 26488 23744 26488 23744 0 _072_
rlabel metal2 28392 22904 28392 22904 0 _073_
rlabel metal2 27384 20608 27384 20608 0 _074_
rlabel metal2 24584 21952 24584 21952 0 _075_
rlabel metal2 29400 27552 29400 27552 0 _076_
rlabel metal2 27720 25984 27720 25984 0 _077_
rlabel metal2 25928 25256 25928 25256 0 _078_
rlabel metal2 25256 24864 25256 24864 0 _079_
rlabel metal2 33208 25816 33208 25816 0 _080_
rlabel metal2 32088 25032 32088 25032 0 _081_
rlabel metal2 37744 21784 37744 21784 0 _082_
rlabel metal2 37016 22904 37016 22904 0 _083_
rlabel metal2 37408 24024 37408 24024 0 _084_
rlabel metal2 36008 25312 36008 25312 0 _085_
rlabel metal2 33992 25144 33992 25144 0 _086_
rlabel metal2 31864 27104 31864 27104 0 _087_
rlabel metal2 34216 21000 34216 21000 0 _088_
rlabel metal2 32088 21728 32088 21728 0 _089_
rlabel metal2 28504 16688 28504 16688 0 _090_
rlabel metal3 27552 20664 27552 20664 0 _091_
rlabel metal2 33096 17192 33096 17192 0 _092_
rlabel metal2 28560 15624 28560 15624 0 _093_
rlabel metal2 36120 18536 36120 18536 0 _094_
rlabel metal2 32200 19432 32200 19432 0 _095_
rlabel metal2 37240 17528 37240 17528 0 _096_
rlabel metal2 35112 20356 35112 20356 0 _097_
rlabel metal2 36008 17864 36008 17864 0 _098_
rlabel metal2 36792 20188 36792 20188 0 _099_
rlabel metal2 33320 12488 33320 12488 0 _100_
rlabel metal2 33096 14056 33096 14056 0 _101_
rlabel metal2 34328 11312 34328 11312 0 _102_
rlabel metal3 32816 13832 32816 13832 0 _103_
rlabel metal3 37576 12600 37576 12600 0 _104_
rlabel metal2 35896 11760 35896 11760 0 _105_
rlabel metal2 37016 13384 37016 13384 0 _106_
rlabel metal2 37912 12768 37912 12768 0 _107_
rlabel metal2 37800 14896 37800 14896 0 _108_
rlabel metal2 33768 15736 33768 15736 0 _109_
rlabel metal2 7560 20440 7560 20440 0 _110_
rlabel metal2 5824 16072 5824 16072 0 _111_
rlabel metal2 7560 16464 7560 16464 0 _112_
rlabel metal2 21560 12544 21560 12544 0 _113_
rlabel metal2 27608 17584 27608 17584 0 _114_
rlabel metal2 1960 23128 1960 23128 0 _115_
rlabel metal2 11032 26208 11032 26208 0 _116_
rlabel metal2 20328 24584 20328 24584 0 _117_
rlabel metal2 27608 21112 27608 21112 0 _118_
rlabel metal2 31752 19880 31752 19880 0 _119_
rlabel metal3 29512 20664 29512 20664 0 _120_
rlabel metal2 33320 14392 33320 14392 0 _121_
rlabel metal2 1736 15400 1736 15400 0 ccff_head
rlabel metal2 37576 17304 37576 17304 0 ccff_tail
rlabel metal3 37464 3752 37464 3752 0 chanx_left_out[16]
rlabel metal3 38682 11480 38682 11480 0 chanx_left_out[17]
rlabel metal3 35448 35112 35448 35112 0 chanx_left_out[18]
rlabel metal2 33656 36232 33656 36232 0 chanx_left_out[19]
rlabel metal2 38248 27720 38248 27720 0 chany_bottom_in[0]
rlabel metal2 28728 36344 28728 36344 0 chany_bottom_in[10]
rlabel metal2 24248 37114 24248 37114 0 chany_bottom_in[12]
rlabel metal2 35784 11200 35784 11200 0 chany_bottom_in[13]
rlabel metal2 37688 32984 37688 32984 0 chany_bottom_in[14]
rlabel metal2 23688 35784 23688 35784 0 chany_bottom_in[16]
rlabel metal2 17976 36456 17976 36456 0 chany_bottom_in[17]
rlabel metal2 26488 5712 26488 5712 0 chany_bottom_in[18]
rlabel metal2 38248 26600 38248 26600 0 chany_bottom_in[1]
rlabel metal3 38528 28616 38528 28616 0 chany_bottom_in[2]
rlabel metal3 38570 1400 38570 1400 0 chany_bottom_in[4]
rlabel metal2 30968 8904 30968 8904 0 chany_bottom_in[5]
rlabel metal3 33992 896 33992 896 0 chany_bottom_in[6]
rlabel metal2 21560 2086 21560 2086 0 chany_bottom_in[8]
rlabel metal2 28952 2058 28952 2058 0 chany_bottom_in[9]
rlabel metal3 32592 4200 32592 4200 0 chany_bottom_out[10]
rlabel metal2 37800 26600 37800 26600 0 chany_bottom_out[11]
rlabel metal2 33656 854 33656 854 0 chany_bottom_out[13]
rlabel metal2 37800 8792 37800 8792 0 chany_bottom_out[14]
rlabel metal2 38416 4872 38416 4872 0 chany_bottom_out[15]
rlabel metal2 30968 37954 30968 37954 0 chany_bottom_out[17]
rlabel metal2 37800 37520 37800 37520 0 chany_bottom_out[18]
rlabel metal2 21336 37184 21336 37184 0 chany_bottom_out[19]
rlabel metal2 28280 2058 28280 2058 0 chany_bottom_out[1]
rlabel metal2 37016 2058 37016 2058 0 chany_bottom_out[2]
rlabel metal2 23128 36904 23128 36904 0 chany_bottom_out[3]
rlabel metal3 30072 3640 30072 3640 0 chany_bottom_out[5]
rlabel metal3 33880 5096 33880 5096 0 chany_bottom_out[6]
rlabel metal2 26152 36624 26152 36624 0 chany_bottom_out[7]
rlabel metal2 37688 36008 37688 36008 0 chany_bottom_out[9]
rlabel metal2 27608 3472 27608 3472 0 chany_top_in[0]
rlabel metal2 38248 29848 38248 29848 0 chany_top_in[10]
rlabel metal2 38248 35560 38248 35560 0 chany_top_in[11]
rlabel metal2 32984 1246 32984 1246 0 chany_top_in[12]
rlabel metal3 38794 10808 38794 10808 0 chany_top_in[13]
rlabel metal2 36344 2058 36344 2058 0 chany_top_in[14]
rlabel metal2 26712 6328 26712 6328 0 chany_top_in[15]
rlabel metal3 30016 36456 30016 36456 0 chany_top_in[16]
rlabel metal2 38192 31080 38192 31080 0 chany_top_in[17]
rlabel metal2 18648 36456 18648 36456 0 chany_top_in[18]
rlabel metal2 34328 1246 34328 1246 0 chany_top_in[19]
rlabel metal2 29288 7000 29288 7000 0 chany_top_in[1]
rlabel metal2 19824 35784 19824 35784 0 chany_top_in[2]
rlabel metal2 30296 2058 30296 2058 0 chany_top_in[4]
rlabel metal2 38360 854 38360 854 0 chany_top_in[5]
rlabel metal2 23016 35784 23016 35784 0 chany_top_in[6]
rlabel metal3 35392 35784 35392 35784 0 chany_top_in[7]
rlabel metal2 38248 29176 38248 29176 0 chany_top_in[8]
rlabel metal2 29736 3696 29736 3696 0 chany_top_in[9]
rlabel metal3 35728 3640 35728 3640 0 chany_top_out[10]
rlabel metal2 28840 36624 28840 36624 0 chany_top_out[11]
rlabel metal2 27832 35784 27832 35784 0 chany_top_out[13]
rlabel metal2 38136 7840 38136 7840 0 chany_top_out[14]
rlabel metal3 33376 36568 33376 36568 0 chany_top_out[15]
rlabel metal2 26040 36456 26040 36456 0 chany_top_out[17]
rlabel metal2 19544 37898 19544 37898 0 chany_top_out[18]
rlabel metal3 37800 10080 37800 10080 0 chany_top_out[19]
rlabel metal2 36456 35952 36456 35952 0 chany_top_out[1]
rlabel metal2 37800 35224 37800 35224 0 chany_top_out[2]
rlabel metal2 37576 36232 37576 36232 0 chany_top_out[3]
rlabel metal2 30520 4704 30520 4704 0 chany_top_out[5]
rlabel metal2 37576 8288 37576 8288 0 chany_top_out[6]
rlabel metal2 37800 7056 37800 7056 0 chany_top_out[7]
rlabel metal2 22232 1526 22232 1526 0 chany_top_out[9]
rlabel metal2 23464 20776 23464 20776 0 clknet_0_prog_clk
rlabel metal2 1848 7924 1848 7924 0 clknet_3_0__leaf_prog_clk
rlabel metal2 20664 17976 20664 17976 0 clknet_3_1__leaf_prog_clk
rlabel metal2 5656 25760 5656 25760 0 clknet_3_2__leaf_prog_clk
rlabel via2 12600 27048 12600 27048 0 clknet_3_3__leaf_prog_clk
rlabel metal2 21112 13328 21112 13328 0 clknet_3_4__leaf_prog_clk
rlabel metal2 34328 16408 34328 16408 0 clknet_3_5__leaf_prog_clk
rlabel metal2 26936 21896 26936 21896 0 clknet_3_6__leaf_prog_clk
rlabel metal3 30016 20776 30016 20776 0 clknet_3_7__leaf_prog_clk
rlabel metal2 23464 16520 23464 16520 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 3080 16352 3080 16352 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal2 11480 15568 11480 15568 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 13048 16268 13048 16268 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 14616 15512 14616 15512 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 7000 17192 7000 17192 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal3 17192 14784 17192 14784 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal3 5656 8120 5656 8120 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal3 4312 17528 4312 17528 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal2 3080 21952 3080 21952 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal2 11480 22400 11480 22400 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal2 8120 26208 8120 26208 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 1568 21784 1568 21784 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal3 1960 24808 1960 24808 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal2 2968 23576 2968 23576 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal2 8456 25704 8456 25704 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal2 5544 26824 5544 26824 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 9128 26656 9128 26656 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal2 12488 28392 12488 28392 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal2 13104 25704 13104 25704 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal2 15288 28000 15288 28000 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal3 17584 28504 17584 28504 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal2 18312 27608 18312 27608 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal2 19768 25256 19768 25256 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal3 22232 25368 22232 25368 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal2 18536 25704 18536 25704 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal2 9128 24584 9128 24584 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal2 15064 25144 15064 25144 0 mem_bottom_track_33.DFFR_5_.Q
rlabel metal2 3080 18424 3080 18424 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal2 5656 22120 5656 22120 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal2 2408 10696 2408 10696 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal2 2968 13944 2968 13944 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal2 3080 19432 3080 19432 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal2 3080 20776 3080 20776 0 mem_left_track_1.DFFR_0_.Q
rlabel metal2 14728 16912 14728 16912 0 mem_left_track_1.DFFR_1_.Q
rlabel metal3 12208 19432 12208 19432 0 mem_left_track_1.DFFR_2_.Q
rlabel metal2 19544 22120 19544 22120 0 mem_left_track_1.DFFR_3_.Q
rlabel metal2 20664 19432 20664 19432 0 mem_left_track_1.DFFR_4_.Q
rlabel metal2 22792 22008 22792 22008 0 mem_left_track_1.DFFR_5_.Q
rlabel metal2 34776 22232 34776 22232 0 mem_left_track_11.DFFR_0_.D
rlabel metal2 31976 19936 31976 19936 0 mem_left_track_11.DFFR_0_.Q
rlabel metal3 29120 18200 29120 18200 0 mem_left_track_11.DFFR_1_.Q
rlabel metal2 33208 8456 33208 8456 0 mem_left_track_13.DFFR_0_.Q
rlabel metal2 26600 10416 26600 10416 0 mem_left_track_13.DFFR_1_.Q
rlabel metal2 30576 7560 30576 7560 0 mem_left_track_15.DFFR_0_.Q
rlabel metal2 30296 8568 30296 8568 0 mem_left_track_15.DFFR_1_.Q
rlabel metal2 26600 8260 26600 8260 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 27720 8008 27720 8008 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 31696 4984 31696 4984 0 mem_left_track_19.DFFR_0_.Q
rlabel metal2 32536 9408 32536 9408 0 mem_left_track_19.DFFR_1_.Q
rlabel metal3 31024 9576 31024 9576 0 mem_left_track_21.DFFR_0_.Q
rlabel metal3 30408 15288 30408 15288 0 mem_left_track_21.DFFR_1_.Q
rlabel metal2 26432 13720 26432 13720 0 mem_left_track_23.DFFR_0_.Q
rlabel metal2 35784 18200 35784 18200 0 mem_left_track_23.DFFR_1_.Q
rlabel metal2 36624 17640 36624 17640 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 37912 16632 37912 16632 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 37240 19768 37240 19768 0 mem_left_track_27.DFFR_0_.Q
rlabel metal2 36344 17416 36344 17416 0 mem_left_track_27.DFFR_1_.Q
rlabel metal4 32984 15148 32984 15148 0 mem_left_track_29.DFFR_0_.Q
rlabel metal2 25256 21140 25256 21140 0 mem_left_track_3.DFFR_0_.Q
rlabel metal2 23464 20356 23464 20356 0 mem_left_track_3.DFFR_1_.Q
rlabel metal2 24808 23744 24808 23744 0 mem_left_track_3.DFFR_2_.Q
rlabel metal3 29120 23688 29120 23688 0 mem_left_track_3.DFFR_3_.Q
rlabel metal2 28840 22344 28840 22344 0 mem_left_track_3.DFFR_4_.Q
rlabel metal2 30184 25816 30184 25816 0 mem_left_track_3.DFFR_5_.Q
rlabel metal2 32760 27048 32760 27048 0 mem_left_track_5.DFFR_0_.Q
rlabel metal2 30408 27720 30408 27720 0 mem_left_track_5.DFFR_1_.Q
rlabel metal3 21728 27944 21728 27944 0 mem_left_track_5.DFFR_2_.Q
rlabel metal2 26040 27888 26040 27888 0 mem_left_track_5.DFFR_3_.Q
rlabel metal2 28840 27496 28840 27496 0 mem_left_track_5.DFFR_4_.Q
rlabel metal2 30072 27944 30072 27944 0 mem_left_track_5.DFFR_5_.Q
rlabel metal3 33376 33208 33376 33208 0 mem_left_track_7.DFFR_0_.Q
rlabel metal2 33040 26488 33040 26488 0 mem_left_track_7.DFFR_1_.Q
rlabel metal2 36792 33320 36792 33320 0 mem_left_track_7.DFFR_2_.Q
rlabel metal3 37240 24920 37240 24920 0 mem_left_track_7.DFFR_3_.Q
rlabel metal2 36792 23352 36792 23352 0 mem_left_track_7.DFFR_4_.Q
rlabel metal2 38248 23184 38248 23184 0 mem_left_track_7.DFFR_5_.Q
rlabel metal2 32648 20748 32648 20748 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 6888 9016 6888 9016 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 5432 12488 5432 12488 0 mem_top_track_0.DFFR_1_.Q
rlabel metal3 6104 5992 6104 5992 0 mem_top_track_0.DFFR_2_.Q
rlabel metal2 5656 5992 5656 5992 0 mem_top_track_0.DFFR_3_.Q
rlabel metal2 6664 6944 6664 6944 0 mem_top_track_0.DFFR_4_.Q
rlabel metal3 3640 10696 3640 10696 0 mem_top_track_0.DFFR_5_.Q
rlabel metal2 11816 7168 11816 7168 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 14392 8456 14392 8456 0 mem_top_track_0.DFFR_7_.Q
rlabel metal2 10416 10696 10416 10696 0 mem_top_track_16.DFFR_0_.D
rlabel metal2 17192 8260 17192 8260 0 mem_top_track_16.DFFR_0_.Q
rlabel metal2 15736 10640 15736 10640 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 23576 9856 23576 9856 0 mem_top_track_16.DFFR_2_.Q
rlabel metal2 19768 8260 19768 8260 0 mem_top_track_16.DFFR_3_.Q
rlabel metal2 22960 10696 22960 10696 0 mem_top_track_16.DFFR_4_.Q
rlabel metal2 26152 11424 26152 11424 0 mem_top_track_16.DFFR_5_.Q
rlabel metal2 24920 12768 24920 12768 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 30408 11200 30408 11200 0 mem_top_track_24.DFFR_1_.Q
rlabel metal2 29960 9688 29960 9688 0 mem_top_track_24.DFFR_2_.Q
rlabel metal2 20720 9688 20720 9688 0 mem_top_track_24.DFFR_3_.Q
rlabel metal2 19432 9688 19432 9688 0 mem_top_track_24.DFFR_4_.Q
rlabel metal2 19656 13552 19656 13552 0 mem_top_track_24.DFFR_5_.Q
rlabel metal2 18312 11032 18312 11032 0 mem_top_track_32.DFFR_0_.Q
rlabel metal2 17864 17192 17864 17192 0 mem_top_track_32.DFFR_1_.Q
rlabel metal3 23408 15400 23408 15400 0 mem_top_track_32.DFFR_2_.Q
rlabel metal3 28056 16968 28056 16968 0 mem_top_track_32.DFFR_3_.Q
rlabel metal2 26152 15400 26152 15400 0 mem_top_track_32.DFFR_4_.Q
rlabel metal2 15736 7000 15736 7000 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 12040 8456 12040 8456 0 mem_top_track_8.DFFR_1_.Q
rlabel metal2 11928 8792 11928 8792 0 mem_top_track_8.DFFR_2_.Q
rlabel metal2 12488 9128 12488 9128 0 mem_top_track_8.DFFR_3_.Q
rlabel metal2 12824 9912 12824 9912 0 mem_top_track_8.DFFR_4_.Q
rlabel metal2 2128 15848 2128 15848 0 net1
rlabel metal3 36400 26488 36400 26488 0 net10
rlabel metal2 18760 8372 18760 8372 0 net100
rlabel metal2 29904 14504 29904 14504 0 net101
rlabel metal2 14952 16968 14952 16968 0 net102
rlabel metal2 19432 14056 19432 14056 0 net103
rlabel metal2 4088 16128 4088 16128 0 net104
rlabel metal2 19208 17584 19208 17584 0 net105
rlabel metal2 29736 26264 29736 26264 0 net106
rlabel metal2 11144 25648 11144 25648 0 net107
rlabel metal2 29624 27272 29624 27272 0 net108
rlabel metal2 7672 23296 7672 23296 0 net109
rlabel metal2 37912 28952 37912 28952 0 net11
rlabel metal2 12264 28448 12264 28448 0 net110
rlabel metal2 4256 15288 4256 15288 0 net111
rlabel metal2 26936 19152 26936 19152 0 net112
rlabel metal2 8008 17192 8008 17192 0 net113
rlabel metal2 20216 12208 20216 12208 0 net114
rlabel metal2 21672 25144 21672 25144 0 net115
rlabel metal2 21336 14616 21336 14616 0 net116
rlabel metal2 6104 13608 6104 13608 0 net117
rlabel metal2 21784 13160 21784 13160 0 net118
rlabel metal2 4760 22456 4760 22456 0 net119
rlabel metal2 37576 4200 37576 4200 0 net12
rlabel metal2 19600 19320 19600 19320 0 net120
rlabel metal2 11816 14448 11816 14448 0 net121
rlabel metal2 11704 8176 11704 8176 0 net122
rlabel metal2 21112 16464 21112 16464 0 net123
rlabel metal2 12152 26320 12152 26320 0 net124
rlabel metal2 4816 16184 4816 16184 0 net125
rlabel metal3 35560 18536 35560 18536 0 net126
rlabel metal2 28504 28504 28504 28504 0 net127
rlabel metal2 8680 27104 8680 27104 0 net128
rlabel metal2 31416 6944 31416 6944 0 net129
rlabel metal3 32424 9128 32424 9128 0 net13
rlabel metal2 27048 28112 27048 28112 0 net130
rlabel metal2 9464 28504 9464 28504 0 net131
rlabel metal2 16968 10640 16968 10640 0 net132
rlabel metal2 11480 10808 11480 10808 0 net133
rlabel metal2 14056 11816 14056 11816 0 net134
rlabel metal2 8680 9968 8680 9968 0 net135
rlabel metal3 34328 19208 34328 19208 0 net136
rlabel metal2 6104 26600 6104 26600 0 net137
rlabel metal2 33432 26824 33432 26824 0 net138
rlabel metal2 22232 22400 22232 22400 0 net139
rlabel metal2 33096 6608 33096 6608 0 net14
rlabel metal2 8456 21616 8456 21616 0 net140
rlabel metal2 8120 12936 8120 12936 0 net141
rlabel metal2 3976 18088 3976 18088 0 net142
rlabel metal2 15512 27048 15512 27048 0 net143
rlabel metal2 24024 24752 24024 24752 0 net144
rlabel metal2 23912 11704 23912 11704 0 net145
rlabel metal3 35672 24696 35672 24696 0 net146
rlabel metal2 10136 13328 10136 13328 0 net147
rlabel metal2 27608 10752 27608 10752 0 net148
rlabel metal2 25704 12992 25704 12992 0 net149
rlabel metal2 22120 5824 22120 5824 0 net15
rlabel metal2 29736 18032 29736 18032 0 net150
rlabel metal2 3808 20888 3808 20888 0 net151
rlabel metal2 22904 17360 22904 17360 0 net152
rlabel metal3 14224 20776 14224 20776 0 net153
rlabel metal2 3752 7392 3752 7392 0 net154
rlabel metal2 33544 28224 33544 28224 0 net155
rlabel metal2 2632 16912 2632 16912 0 net156
rlabel metal3 33096 13048 33096 13048 0 net157
rlabel metal3 18704 21224 18704 21224 0 net158
rlabel metal2 26600 15064 26600 15064 0 net159
rlabel metal3 28672 4536 28672 4536 0 net16
rlabel metal2 16744 16184 16744 16184 0 net160
rlabel metal3 12152 10472 12152 10472 0 net161
rlabel metal2 35504 21560 35504 21560 0 net162
rlabel metal2 33656 24192 33656 24192 0 net163
rlabel metal2 19768 11312 19768 11312 0 net164
rlabel metal2 23016 27384 23016 27384 0 net165
rlabel metal2 32368 5208 32368 5208 0 net166
rlabel metal2 34384 27720 34384 27720 0 net167
rlabel metal2 7672 8680 7672 8680 0 net168
rlabel metal2 4088 24360 4088 24360 0 net169
rlabel metal2 27832 4200 27832 4200 0 net17
rlabel metal2 34328 6160 34328 6160 0 net170
rlabel metal2 9912 16912 9912 16912 0 net171
rlabel metal2 26824 11704 26824 11704 0 net172
rlabel metal2 16856 7588 16856 7588 0 net173
rlabel metal3 26992 18984 26992 18984 0 net174
rlabel metal3 5040 21336 5040 21336 0 net175
rlabel metal2 27608 8680 27608 8680 0 net176
rlabel metal2 4088 18256 4088 18256 0 net177
rlabel metal2 27160 28280 27160 28280 0 net178
rlabel metal2 35952 26264 35952 26264 0 net179
rlabel metal2 37912 30464 37912 30464 0 net18
rlabel metal2 17864 25816 17864 25816 0 net180
rlabel metal2 15960 17696 15960 17696 0 net181
rlabel metal2 25816 22176 25816 22176 0 net182
rlabel metal2 3416 11200 3416 11200 0 net183
rlabel metal2 13048 27384 13048 27384 0 net184
rlabel metal2 15960 9352 15960 9352 0 net185
rlabel metal2 32536 6776 32536 6776 0 net186
rlabel metal2 33936 18424 33936 18424 0 net187
rlabel metal3 22400 20216 22400 20216 0 net188
rlabel metal2 10024 26432 10024 26432 0 net189
rlabel metal3 37912 31528 37912 31528 0 net19
rlabel metal3 35504 16856 35504 16856 0 net190
rlabel metal2 31584 7336 31584 7336 0 net191
rlabel metal2 16072 25592 16072 25592 0 net192
rlabel metal2 8568 17640 8568 17640 0 net193
rlabel metal2 16744 24864 16744 24864 0 net194
rlabel metal2 3528 24024 3528 24024 0 net195
rlabel metal2 27160 24360 27160 24360 0 net196
rlabel metal2 34664 24024 34664 24024 0 net197
rlabel metal3 34776 15176 34776 15176 0 net198
rlabel metal3 4088 25592 4088 25592 0 net199
rlabel metal3 36344 28056 36344 28056 0 net2
rlabel metal2 27384 4760 27384 4760 0 net20
rlabel metal3 10808 21448 10808 21448 0 net200
rlabel metal2 8008 6776 8008 6776 0 net201
rlabel metal2 2296 14168 2296 14168 0 net202
rlabel metal2 7896 7840 7896 7840 0 net203
rlabel metal2 26712 14896 26712 14896 0 net204
rlabel metal3 30800 7336 30800 7336 0 net205
rlabel metal2 2296 7896 2296 7896 0 net206
rlabel metal3 33096 8232 33096 8232 0 net21
rlabel metal2 26544 4312 26544 4312 0 net22
rlabel metal2 28392 4536 28392 4536 0 net23
rlabel metal2 30520 35952 30520 35952 0 net24
rlabel metal2 37912 31248 37912 31248 0 net25
rlabel metal3 20272 35784 20272 35784 0 net26
rlabel metal2 26936 4424 26936 4424 0 net27
rlabel metal2 27944 7560 27944 7560 0 net28
rlabel metal2 21224 35840 21224 35840 0 net29
rlabel metal2 28952 36120 28952 36120 0 net3
rlabel metal2 28840 6328 28840 6328 0 net30
rlabel metal2 29512 7112 29512 7112 0 net31
rlabel metal3 24416 34888 24416 34888 0 net32
rlabel metal2 32424 35336 32424 35336 0 net33
rlabel metal2 37912 29736 37912 29736 0 net34
rlabel metal3 30128 3528 30128 3528 0 net35
rlabel metal2 30856 16184 30856 16184 0 net36
rlabel metal2 38304 17640 38304 17640 0 net37
rlabel metal2 27160 3752 27160 3752 0 net38
rlabel metal2 26376 5432 26376 5432 0 net39
rlabel metal3 25760 34776 25760 34776 0 net4
rlabel metal3 37128 33208 37128 33208 0 net40
rlabel metal2 32648 35224 32648 35224 0 net41
rlabel metal2 32592 3416 32592 3416 0 net42
rlabel metal2 37016 26880 37016 26880 0 net43
rlabel metal2 27720 5376 27720 5376 0 net44
rlabel metal3 33544 8008 33544 8008 0 net45
rlabel metal3 28056 4480 28056 4480 0 net46
rlabel metal2 30744 36064 30744 36064 0 net47
rlabel metal2 36568 33432 36568 33432 0 net48
rlabel metal2 22232 36176 22232 36176 0 net49
rlabel metal2 26824 5936 26824 5936 0 net5
rlabel metal2 28616 4200 28616 4200 0 net50
rlabel metal2 31192 5096 31192 5096 0 net51
rlabel metal2 21560 36064 21560 36064 0 net52
rlabel metal2 30072 3808 30072 3808 0 net53
rlabel metal2 35560 9240 35560 9240 0 net54
rlabel metal2 25704 35616 25704 35616 0 net55
rlabel metal2 37016 35168 37016 35168 0 net56
rlabel metal2 36008 4088 36008 4088 0 net57
rlabel metal2 27944 36232 27944 36232 0 net58
rlabel metal2 27048 35224 27048 35224 0 net59
rlabel metal2 31640 33432 31640 33432 0 net6
rlabel metal2 27048 5376 27048 5376 0 net60
rlabel metal3 32872 35896 32872 35896 0 net61
rlabel metal2 26376 35224 26376 35224 0 net62
rlabel metal2 20552 36176 20552 36176 0 net63
rlabel metal2 33432 8624 33432 8624 0 net64
rlabel metal2 35336 35224 35336 35224 0 net65
rlabel metal2 34776 34832 34776 34832 0 net66
rlabel metal3 36288 33320 36288 33320 0 net67
rlabel metal2 29848 5376 29848 5376 0 net68
rlabel metal2 33992 9632 33992 9632 0 net69
rlabel metal2 26152 35336 26152 35336 0 net7
rlabel metal2 33432 6272 33432 6272 0 net70
rlabel metal2 22456 5768 22456 5768 0 net71
rlabel metal2 37128 30856 37128 30856 0 net72
rlabel metal2 22904 1470 22904 1470 0 net73
rlabel metal2 37632 29624 37632 29624 0 net74
rlabel metal2 37576 30184 37576 30184 0 net75
rlabel metal2 24248 2030 24248 2030 0 net76
rlabel metal2 22568 36400 22568 36400 0 net77
rlabel metal2 29736 35896 29736 35896 0 net78
rlabel metal3 37170 2744 37170 2744 0 net79
rlabel metal2 20776 35952 20776 35952 0 net8
rlabel metal2 36456 31304 36456 31304 0 net80
rlabel metal2 35336 32648 35336 32648 0 net81
rlabel metal2 29960 36512 29960 36512 0 net82
rlabel metal2 37576 25984 37576 25984 0 net83
rlabel metal3 38346 56 38346 56 0 net84
rlabel metal2 33656 34440 33656 34440 0 net85
rlabel metal3 35112 34216 35112 34216 0 net86
rlabel metal3 35728 34776 35728 34776 0 net87
rlabel metal3 34776 36344 34776 36344 0 net88
rlabel metal3 31304 4760 31304 4760 0 net89
rlabel metal3 30352 6104 30352 6104 0 net9
rlabel metal2 36400 9576 36400 9576 0 net90
rlabel metal3 37912 32760 37912 32760 0 net91
rlabel metal2 33992 34944 33992 34944 0 net92
rlabel metal2 26712 2520 26712 2520 0 net93
rlabel metal2 33320 8008 33320 8008 0 net94
rlabel metal2 31640 37786 31640 37786 0 net95
rlabel metal2 35000 33208 35000 33208 0 net96
rlabel metal2 26712 37072 26712 37072 0 net97
rlabel metal2 32200 17304 32200 17304 0 net98
rlabel metal3 34272 17080 34272 17080 0 net99
rlabel metal2 38360 20356 38360 20356 0 pReset
rlabel metal3 2534 26264 2534 26264 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
