VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 170.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 114.240 170.000 114.800 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 166.000 44.240 170.000 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.080 4.000 10.640 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 166.000 124.880 170.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 137.760 170.000 138.320 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 166.000 47.600 170.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 166.000 3.920 170.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 157.920 170.000 158.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 3.360 170.000 3.920 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 166.000 40.880 170.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 127.680 170.000 128.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 166.000 94.640 170.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 166.000 141.680 170.000 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 166.000 64.400 170.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 166.000 77.840 170.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 154.560 170.000 155.120 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 166.000 81.200 170.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 141.120 170.000 141.680 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 166.000 128.240 170.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 166.000 10.640 170.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.440 4.000 14.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 36.960 170.000 37.520 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 20.160 170.000 20.720 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 166.000 34.160 170.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 166.000 134.960 170.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 166.000 50.960 170.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 134.400 170.000 134.960 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 166.000 84.560 170.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 30.240 170.000 30.800 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 166.000 27.440 170.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 26.880 170.000 27.440 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 166.000 30.800 170.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 23.520 170.000 24.080 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 166.000 17.360 170.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 166.000 138.320 170.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 166.000 61.040 170.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 166.000 14.000 170.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 10.080 170.000 10.640 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 166.000 20.720 170.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 166.000 131.600 170.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 166.000 54.320 170.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 131.040 170.000 131.600 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 166.000 91.280 170.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 33.600 170.000 34.160 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 6.720 170.000 7.280 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 16.800 170.000 17.360 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 166.000 24.080 170.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 166.000 57.680 170.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 166.000 145.040 170.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 166.000 74.480 170.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 151.200 170.000 151.760 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 147.840 170.000 148.400 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 166.000 71.120 170.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 166.000 87.920 170.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 166.000 37.520 170.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 144.480 170.000 145.040 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 13.440 170.000 14.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 166.000 7.280 170.000 ;
    END
  END chany_top_out[9]
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 166.000 67.760 170.000 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END prog_clk
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
  PIN top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 40.320 170.000 40.880 ;
    END
  END top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
  PIN top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 0.000 170.000 0.560 ;
    END
  END top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 25.450 15.380 27.050 153.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.510 15.380 66.110 153.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.570 15.380 105.170 153.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 142.630 15.380 144.230 153.180 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 44.980 15.380 46.580 153.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 84.040 15.380 85.640 153.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 123.100 15.380 124.700 153.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.160 15.380 163.760 153.180 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 163.760 153.850 ;
      LAYER Metal2 ;
        RECT 0.700 165.700 3.060 166.000 ;
        RECT 4.220 165.700 6.420 166.000 ;
        RECT 7.580 165.700 9.780 166.000 ;
        RECT 10.940 165.700 13.140 166.000 ;
        RECT 14.300 165.700 16.500 166.000 ;
        RECT 17.660 165.700 19.860 166.000 ;
        RECT 21.020 165.700 23.220 166.000 ;
        RECT 24.380 165.700 26.580 166.000 ;
        RECT 27.740 165.700 29.940 166.000 ;
        RECT 31.100 165.700 33.300 166.000 ;
        RECT 34.460 165.700 36.660 166.000 ;
        RECT 37.820 165.700 40.020 166.000 ;
        RECT 41.180 165.700 43.380 166.000 ;
        RECT 44.540 165.700 46.740 166.000 ;
        RECT 47.900 165.700 50.100 166.000 ;
        RECT 51.260 165.700 53.460 166.000 ;
        RECT 54.620 165.700 56.820 166.000 ;
        RECT 57.980 165.700 60.180 166.000 ;
        RECT 61.340 165.700 63.540 166.000 ;
        RECT 64.700 165.700 66.900 166.000 ;
        RECT 68.060 165.700 70.260 166.000 ;
        RECT 71.420 165.700 73.620 166.000 ;
        RECT 74.780 165.700 76.980 166.000 ;
        RECT 78.140 165.700 80.340 166.000 ;
        RECT 81.500 165.700 83.700 166.000 ;
        RECT 84.860 165.700 87.060 166.000 ;
        RECT 88.220 165.700 90.420 166.000 ;
        RECT 91.580 165.700 93.780 166.000 ;
        RECT 94.940 165.700 124.020 166.000 ;
        RECT 125.180 165.700 127.380 166.000 ;
        RECT 128.540 165.700 130.740 166.000 ;
        RECT 131.900 165.700 134.100 166.000 ;
        RECT 135.260 165.700 137.460 166.000 ;
        RECT 138.620 165.700 140.820 166.000 ;
        RECT 141.980 165.700 144.180 166.000 ;
        RECT 145.340 165.700 163.620 166.000 ;
        RECT 0.700 4.300 163.620 165.700 ;
        RECT 0.860 3.450 3.060 4.300 ;
        RECT 4.220 3.450 6.420 4.300 ;
        RECT 7.580 3.450 9.780 4.300 ;
        RECT 10.940 3.450 13.140 4.300 ;
        RECT 14.300 3.450 16.500 4.300 ;
        RECT 17.660 3.450 19.860 4.300 ;
        RECT 21.020 3.450 23.220 4.300 ;
        RECT 24.380 3.450 26.580 4.300 ;
        RECT 27.740 3.450 29.940 4.300 ;
        RECT 31.100 3.450 33.300 4.300 ;
        RECT 34.460 3.450 36.660 4.300 ;
        RECT 37.820 3.450 40.020 4.300 ;
        RECT 41.180 3.450 43.380 4.300 ;
        RECT 44.540 3.450 46.740 4.300 ;
        RECT 47.900 3.450 50.100 4.300 ;
        RECT 51.260 3.450 53.460 4.300 ;
        RECT 54.620 3.450 56.820 4.300 ;
        RECT 57.980 3.450 60.180 4.300 ;
        RECT 61.340 3.450 63.540 4.300 ;
        RECT 64.700 3.450 66.900 4.300 ;
        RECT 68.060 3.450 70.260 4.300 ;
        RECT 71.420 3.450 73.620 4.300 ;
        RECT 74.780 3.450 76.980 4.300 ;
        RECT 78.140 3.450 80.340 4.300 ;
        RECT 81.500 3.450 83.700 4.300 ;
        RECT 84.860 3.450 87.060 4.300 ;
        RECT 88.220 3.450 90.420 4.300 ;
        RECT 91.580 3.450 93.780 4.300 ;
        RECT 94.940 3.450 97.140 4.300 ;
        RECT 98.300 3.450 100.500 4.300 ;
        RECT 101.660 3.450 103.860 4.300 ;
        RECT 105.020 3.450 107.220 4.300 ;
        RECT 108.380 3.450 110.580 4.300 ;
        RECT 111.740 3.450 113.940 4.300 ;
        RECT 115.100 3.450 117.300 4.300 ;
        RECT 118.460 3.450 120.660 4.300 ;
        RECT 121.820 3.450 124.020 4.300 ;
        RECT 125.180 3.450 127.380 4.300 ;
        RECT 128.540 3.450 130.740 4.300 ;
        RECT 131.900 3.450 134.100 4.300 ;
        RECT 135.260 3.450 137.460 4.300 ;
        RECT 138.620 3.450 140.820 4.300 ;
        RECT 141.980 3.450 144.180 4.300 ;
        RECT 145.340 3.450 147.540 4.300 ;
        RECT 148.700 3.450 150.900 4.300 ;
        RECT 152.060 3.450 154.260 4.300 ;
        RECT 155.420 3.450 157.620 4.300 ;
        RECT 158.780 3.450 160.980 4.300 ;
        RECT 162.140 3.450 163.620 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 167.700 166.000 168.420 ;
        RECT 0.650 165.500 166.000 167.700 ;
        RECT 4.300 164.340 166.000 165.500 ;
        RECT 0.650 162.140 166.000 164.340 ;
        RECT 4.300 160.980 166.000 162.140 ;
        RECT 0.650 158.780 166.000 160.980 ;
        RECT 4.300 157.620 165.700 158.780 ;
        RECT 0.650 155.420 166.000 157.620 ;
        RECT 4.300 154.260 165.700 155.420 ;
        RECT 0.650 152.060 166.000 154.260 ;
        RECT 4.300 150.900 165.700 152.060 ;
        RECT 0.650 148.700 166.000 150.900 ;
        RECT 4.300 147.540 165.700 148.700 ;
        RECT 0.650 145.340 166.000 147.540 ;
        RECT 4.300 144.180 165.700 145.340 ;
        RECT 0.650 141.980 166.000 144.180 ;
        RECT 4.300 140.820 165.700 141.980 ;
        RECT 0.650 138.620 166.000 140.820 ;
        RECT 4.300 137.460 165.700 138.620 ;
        RECT 0.650 135.260 166.000 137.460 ;
        RECT 4.300 134.100 165.700 135.260 ;
        RECT 0.650 131.900 166.000 134.100 ;
        RECT 4.300 130.740 165.700 131.900 ;
        RECT 0.650 128.540 166.000 130.740 ;
        RECT 4.300 127.380 165.700 128.540 ;
        RECT 0.650 125.180 166.000 127.380 ;
        RECT 4.300 124.020 166.000 125.180 ;
        RECT 0.650 121.820 166.000 124.020 ;
        RECT 4.300 120.660 166.000 121.820 ;
        RECT 0.650 118.460 166.000 120.660 ;
        RECT 4.300 117.300 166.000 118.460 ;
        RECT 0.650 115.100 166.000 117.300 ;
        RECT 4.300 113.940 165.700 115.100 ;
        RECT 0.650 111.740 166.000 113.940 ;
        RECT 4.300 110.580 166.000 111.740 ;
        RECT 0.650 108.380 166.000 110.580 ;
        RECT 4.300 107.220 166.000 108.380 ;
        RECT 0.650 105.020 166.000 107.220 ;
        RECT 4.300 103.860 166.000 105.020 ;
        RECT 0.650 101.660 166.000 103.860 ;
        RECT 4.300 100.500 166.000 101.660 ;
        RECT 0.650 98.300 166.000 100.500 ;
        RECT 4.300 97.140 166.000 98.300 ;
        RECT 0.650 41.180 166.000 97.140 ;
        RECT 0.650 40.020 165.700 41.180 ;
        RECT 0.650 37.820 166.000 40.020 ;
        RECT 0.650 36.660 165.700 37.820 ;
        RECT 0.650 34.460 166.000 36.660 ;
        RECT 4.300 33.300 165.700 34.460 ;
        RECT 0.650 31.100 166.000 33.300 ;
        RECT 4.300 29.940 165.700 31.100 ;
        RECT 0.650 27.740 166.000 29.940 ;
        RECT 4.300 26.580 165.700 27.740 ;
        RECT 0.650 24.380 166.000 26.580 ;
        RECT 4.300 23.220 165.700 24.380 ;
        RECT 0.650 21.020 166.000 23.220 ;
        RECT 4.300 19.860 165.700 21.020 ;
        RECT 0.650 17.660 166.000 19.860 ;
        RECT 4.300 16.500 165.700 17.660 ;
        RECT 0.650 14.300 166.000 16.500 ;
        RECT 4.300 13.140 165.700 14.300 ;
        RECT 0.650 10.940 166.000 13.140 ;
        RECT 4.300 9.780 165.700 10.940 ;
        RECT 0.650 7.580 166.000 9.780 ;
        RECT 0.650 6.420 165.700 7.580 ;
        RECT 0.650 4.220 166.000 6.420 ;
        RECT 0.650 3.500 165.700 4.220 ;
      LAYER Metal4 ;
        RECT 9.660 18.010 25.060 145.510 ;
  END
END sb_0__1_
END LIBRARY

