// This is the unpowered netlist.
module sb_1__1_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    ccff_head,
    ccff_tail,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input ccff_head;
 output ccff_tail;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input [19:0] chanx_left_in;
 output [19:0] chanx_left_out;
 input [19:0] chanx_right_in;
 output [19:0] chanx_right_out;
 input [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;
 input [19:0] chany_top_in;
 output [19:0] chany_top_out;

 wire net143;
 wire net140;
 wire net139;
 wire net142;
 wire net141;
 wire net138;
 wire net135;
 wire net134;
 wire net137;
 wire net136;
 wire net133;
 wire net130;
 wire net129;
 wire net132;
 wire net131;
 wire net128;
 wire net125;
 wire net124;
 wire net127;
 wire net126;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire clknet_0_prog_clk;
 wire clknet_4_0_0_prog_clk;
 wire clknet_4_10_0_prog_clk;
 wire clknet_4_11_0_prog_clk;
 wire clknet_4_12_0_prog_clk;
 wire clknet_4_13_0_prog_clk;
 wire clknet_4_14_0_prog_clk;
 wire clknet_4_15_0_prog_clk;
 wire clknet_4_1_0_prog_clk;
 wire clknet_4_2_0_prog_clk;
 wire clknet_4_3_0_prog_clk;
 wire clknet_4_4_0_prog_clk;
 wire clknet_4_5_0_prog_clk;
 wire clknet_4_6_0_prog_clk;
 wire clknet_4_7_0_prog_clk;
 wire clknet_4_8_0_prog_clk;
 wire clknet_4_9_0_prog_clk;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_1.DFFR_2_.Q ;
 wire \mem_bottom_track_1.DFFR_3_.Q ;
 wire \mem_bottom_track_1.DFFR_4_.Q ;
 wire \mem_bottom_track_1.DFFR_5_.Q ;
 wire \mem_bottom_track_1.DFFR_6_.Q ;
 wire \mem_bottom_track_1.DFFR_7_.Q ;
 wire \mem_bottom_track_17.DFFR_0_.D ;
 wire \mem_bottom_track_17.DFFR_0_.Q ;
 wire \mem_bottom_track_17.DFFR_1_.Q ;
 wire \mem_bottom_track_17.DFFR_2_.Q ;
 wire \mem_bottom_track_17.DFFR_3_.Q ;
 wire \mem_bottom_track_17.DFFR_4_.Q ;
 wire \mem_bottom_track_17.DFFR_5_.Q ;
 wire \mem_bottom_track_17.DFFR_6_.Q ;
 wire \mem_bottom_track_17.DFFR_7_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_2_.Q ;
 wire \mem_bottom_track_25.DFFR_3_.Q ;
 wire \mem_bottom_track_25.DFFR_4_.Q ;
 wire \mem_bottom_track_25.DFFR_5_.Q ;
 wire \mem_bottom_track_25.DFFR_6_.Q ;
 wire \mem_bottom_track_25.DFFR_7_.Q ;
 wire \mem_bottom_track_33.DFFR_0_.Q ;
 wire \mem_bottom_track_33.DFFR_1_.Q ;
 wire \mem_bottom_track_33.DFFR_2_.Q ;
 wire \mem_bottom_track_33.DFFR_3_.Q ;
 wire \mem_bottom_track_33.DFFR_4_.Q ;
 wire \mem_bottom_track_33.DFFR_5_.Q ;
 wire \mem_bottom_track_33.DFFR_6_.Q ;
 wire \mem_bottom_track_33.DFFR_7_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_bottom_track_9.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_2_.Q ;
 wire \mem_bottom_track_9.DFFR_3_.Q ;
 wire \mem_bottom_track_9.DFFR_4_.Q ;
 wire \mem_bottom_track_9.DFFR_5_.Q ;
 wire \mem_bottom_track_9.DFFR_6_.Q ;
 wire \mem_left_track_1.DFFR_0_.Q ;
 wire \mem_left_track_1.DFFR_1_.Q ;
 wire \mem_left_track_1.DFFR_2_.Q ;
 wire \mem_left_track_1.DFFR_3_.Q ;
 wire \mem_left_track_1.DFFR_4_.Q ;
 wire \mem_left_track_1.DFFR_5_.Q ;
 wire \mem_left_track_1.DFFR_6_.Q ;
 wire \mem_left_track_1.DFFR_7_.Q ;
 wire \mem_left_track_17.DFFR_0_.D ;
 wire \mem_left_track_17.DFFR_0_.Q ;
 wire \mem_left_track_17.DFFR_1_.Q ;
 wire \mem_left_track_17.DFFR_2_.Q ;
 wire \mem_left_track_17.DFFR_3_.Q ;
 wire \mem_left_track_17.DFFR_4_.Q ;
 wire \mem_left_track_17.DFFR_5_.Q ;
 wire \mem_left_track_17.DFFR_6_.Q ;
 wire \mem_left_track_17.DFFR_7_.Q ;
 wire \mem_left_track_25.DFFR_0_.Q ;
 wire \mem_left_track_25.DFFR_1_.Q ;
 wire \mem_left_track_25.DFFR_2_.Q ;
 wire \mem_left_track_25.DFFR_3_.Q ;
 wire \mem_left_track_25.DFFR_4_.Q ;
 wire \mem_left_track_25.DFFR_5_.Q ;
 wire \mem_left_track_25.DFFR_6_.Q ;
 wire \mem_left_track_25.DFFR_7_.Q ;
 wire \mem_left_track_33.DFFR_0_.Q ;
 wire \mem_left_track_33.DFFR_1_.Q ;
 wire \mem_left_track_33.DFFR_2_.Q ;
 wire \mem_left_track_33.DFFR_3_.Q ;
 wire \mem_left_track_33.DFFR_4_.Q ;
 wire \mem_left_track_33.DFFR_5_.Q ;
 wire \mem_left_track_33.DFFR_6_.Q ;
 wire \mem_left_track_9.DFFR_0_.Q ;
 wire \mem_left_track_9.DFFR_1_.Q ;
 wire \mem_left_track_9.DFFR_2_.Q ;
 wire \mem_left_track_9.DFFR_3_.Q ;
 wire \mem_left_track_9.DFFR_4_.Q ;
 wire \mem_left_track_9.DFFR_5_.Q ;
 wire \mem_left_track_9.DFFR_6_.Q ;
 wire \mem_right_track_0.DFFR_0_.D ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_0.DFFR_2_.Q ;
 wire \mem_right_track_0.DFFR_3_.Q ;
 wire \mem_right_track_0.DFFR_4_.Q ;
 wire \mem_right_track_0.DFFR_5_.Q ;
 wire \mem_right_track_0.DFFR_6_.Q ;
 wire \mem_right_track_0.DFFR_7_.Q ;
 wire \mem_right_track_16.DFFR_0_.D ;
 wire \mem_right_track_16.DFFR_0_.Q ;
 wire \mem_right_track_16.DFFR_1_.Q ;
 wire \mem_right_track_16.DFFR_2_.Q ;
 wire \mem_right_track_16.DFFR_3_.Q ;
 wire \mem_right_track_16.DFFR_4_.Q ;
 wire \mem_right_track_16.DFFR_5_.Q ;
 wire \mem_right_track_16.DFFR_6_.Q ;
 wire \mem_right_track_16.DFFR_7_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_2_.Q ;
 wire \mem_right_track_24.DFFR_3_.Q ;
 wire \mem_right_track_24.DFFR_4_.Q ;
 wire \mem_right_track_24.DFFR_5_.Q ;
 wire \mem_right_track_24.DFFR_6_.Q ;
 wire \mem_right_track_24.DFFR_7_.Q ;
 wire \mem_right_track_32.DFFR_0_.Q ;
 wire \mem_right_track_32.DFFR_1_.Q ;
 wire \mem_right_track_32.DFFR_2_.Q ;
 wire \mem_right_track_32.DFFR_3_.Q ;
 wire \mem_right_track_32.DFFR_4_.Q ;
 wire \mem_right_track_32.DFFR_5_.Q ;
 wire \mem_right_track_32.DFFR_6_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire \mem_right_track_8.DFFR_1_.Q ;
 wire \mem_right_track_8.DFFR_2_.Q ;
 wire \mem_right_track_8.DFFR_3_.Q ;
 wire \mem_right_track_8.DFFR_4_.Q ;
 wire \mem_right_track_8.DFFR_5_.Q ;
 wire \mem_right_track_8.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_0.DFFR_2_.Q ;
 wire \mem_top_track_0.DFFR_3_.Q ;
 wire \mem_top_track_0.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_5_.Q ;
 wire \mem_top_track_0.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_7_.Q ;
 wire \mem_top_track_16.DFFR_0_.D ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_2_.Q ;
 wire \mem_top_track_16.DFFR_3_.Q ;
 wire \mem_top_track_16.DFFR_4_.Q ;
 wire \mem_top_track_16.DFFR_5_.Q ;
 wire \mem_top_track_16.DFFR_6_.Q ;
 wire \mem_top_track_16.DFFR_7_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_2_.Q ;
 wire \mem_top_track_24.DFFR_3_.Q ;
 wire \mem_top_track_24.DFFR_4_.Q ;
 wire \mem_top_track_24.DFFR_5_.Q ;
 wire \mem_top_track_24.DFFR_6_.Q ;
 wire \mem_top_track_24.DFFR_7_.Q ;
 wire \mem_top_track_32.DFFR_0_.Q ;
 wire \mem_top_track_32.DFFR_1_.Q ;
 wire \mem_top_track_32.DFFR_2_.Q ;
 wire \mem_top_track_32.DFFR_3_.Q ;
 wire \mem_top_track_32.DFFR_4_.Q ;
 wire \mem_top_track_32.DFFR_5_.Q ;
 wire \mem_top_track_32.DFFR_6_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire \mem_top_track_8.DFFR_1_.Q ;
 wire \mem_top_track_8.DFFR_2_.Q ;
 wire \mem_top_track_8.DFFR_3_.Q ;
 wire \mem_top_track_8.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_5_.Q ;
 wire \mem_top_track_8.DFFR_6_.Q ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net13;
 wire net14;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__I (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__191__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__213__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__I (.I(_166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__I (.I(_161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__I (.I(_177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__D (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__CLK (.I(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__CLK (.I(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__D (.I(\mem_left_track_17.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__CLK (.I(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__577__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(chanx_left_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(chanx_left_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(chanx_left_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(chanx_left_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(chanx_left_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(chanx_left_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(chanx_left_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(chanx_right_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(chanx_right_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(chanx_right_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(chanx_right_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(chanx_right_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(chanx_right_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(chanx_right_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(chanx_right_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(chanx_right_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(chanx_right_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(chanx_right_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(chanx_right_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(chanx_right_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(chanx_left_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(chanx_right_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(chanx_right_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(chany_bottom_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(chany_bottom_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(chany_bottom_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(chany_bottom_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(chany_bottom_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(chany_bottom_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(chany_bottom_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(chany_bottom_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(chanx_left_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(chany_bottom_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(chany_bottom_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(chany_bottom_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(chany_bottom_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(chany_bottom_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(chany_bottom_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(chany_bottom_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(chany_top_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(chany_top_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(chany_top_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(chanx_left_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(chany_top_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(chany_top_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(chany_top_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(chany_top_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(chany_top_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(chany_top_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(chany_top_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(chany_top_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(chany_top_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(chany_top_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(chanx_left_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(chany_top_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(chany_top_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(chanx_left_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(chanx_left_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(chanx_left_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(chanx_left_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_165 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _178_ (.I(net62),
    .Z(_160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _179_ (.I(_160_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _180_ (.I(_161_),
    .Z(_162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _181_ (.I(_162_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _182_ (.I(_162_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _183_ (.I(_162_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _184_ (.I(_162_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _185_ (.I(_162_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _186_ (.I(_162_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _187_ (.I(_162_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _188_ (.I(_162_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _189_ (.I(_162_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _190_ (.I(_162_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _191_ (.I(_161_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _192_ (.I(_163_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _193_ (.I(_163_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _194_ (.I(_163_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _195_ (.I(_163_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _196_ (.I(_163_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _197_ (.I(_163_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _198_ (.I(_163_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _199_ (.I(_163_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _200_ (.I(_163_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _201_ (.I(_163_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _202_ (.I(_161_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _203_ (.I(_164_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _204_ (.I(_164_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _205_ (.I(_164_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _206_ (.I(_164_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _207_ (.I(_164_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _208_ (.I(_164_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _209_ (.I(_164_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _210_ (.I(_164_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _211_ (.I(_164_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _212_ (.I(_164_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _213_ (.I(_161_),
    .Z(_165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _214_ (.I(_165_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _215_ (.I(_165_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _216_ (.I(_165_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _217_ (.I(_165_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _218_ (.I(_165_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _219_ (.I(_165_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _220_ (.I(_165_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _221_ (.I(_165_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _222_ (.I(_165_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _223_ (.I(_165_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _224_ (.I(_161_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _225_ (.I(_166_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _226_ (.I(_166_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _227_ (.I(_166_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _228_ (.I(_166_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _229_ (.I(_166_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _230_ (.I(_166_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _231_ (.I(_166_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _232_ (.I(_166_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _233_ (.I(_166_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _234_ (.I(_166_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _235_ (.I(_161_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _236_ (.I(_167_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _237_ (.I(_167_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _238_ (.I(_167_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _239_ (.I(_167_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _240_ (.I(_167_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _241_ (.I(_167_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _242_ (.I(_167_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _243_ (.I(_167_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _244_ (.I(_167_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _245_ (.I(_167_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _246_ (.I(_161_),
    .Z(_168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _247_ (.I(_168_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _248_ (.I(_168_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _249_ (.I(_168_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _250_ (.I(_168_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _251_ (.I(_168_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _252_ (.I(_168_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _253_ (.I(_168_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _254_ (.I(_168_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _255_ (.I(_168_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _256_ (.I(_168_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _257_ (.I(_161_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _258_ (.I(_169_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _259_ (.I(_169_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _260_ (.I(_169_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _261_ (.I(_169_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _262_ (.I(_169_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _263_ (.I(_169_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _264_ (.I(_169_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _265_ (.I(_169_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _266_ (.I(_169_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _267_ (.I(_169_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _268_ (.I(_161_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _269_ (.I(_170_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _270_ (.I(_170_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _271_ (.I(_170_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _272_ (.I(_170_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _273_ (.I(_170_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _274_ (.I(_170_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _275_ (.I(_170_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _276_ (.I(_170_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _277_ (.I(_170_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _278_ (.I(_170_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _279_ (.I(_161_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _280_ (.I(_171_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _281_ (.I(_171_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _282_ (.I(_171_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _283_ (.I(_171_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _284_ (.I(_171_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _285_ (.I(_171_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _286_ (.I(_171_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _287_ (.I(_171_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _288_ (.I(_171_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _289_ (.I(_171_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _290_ (.I(_160_),
    .Z(_172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _291_ (.I(_172_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _292_ (.I(_172_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _293_ (.I(_172_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _294_ (.I(_172_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _295_ (.I(_172_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _296_ (.I(_172_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _297_ (.I(_172_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _298_ (.I(_172_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _299_ (.I(_172_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _300_ (.I(_172_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _301_ (.I(_160_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _302_ (.I(_173_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _303_ (.I(_173_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _304_ (.I(_173_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _305_ (.I(_173_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _306_ (.I(_173_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _307_ (.I(_173_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _308_ (.I(_173_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _309_ (.I(_173_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _310_ (.I(_173_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _311_ (.I(_173_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _312_ (.I(_160_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _313_ (.I(_174_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _314_ (.I(_174_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _315_ (.I(_174_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _316_ (.I(_174_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _317_ (.I(_174_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _318_ (.I(_174_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _319_ (.I(_174_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _320_ (.I(_174_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _321_ (.I(_174_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _322_ (.I(_174_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _323_ (.I(_160_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _324_ (.I(_175_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _325_ (.I(_175_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _326_ (.I(_175_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _327_ (.I(_175_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _328_ (.I(_175_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _329_ (.I(_175_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _330_ (.I(_175_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _331_ (.I(_175_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _332_ (.I(_175_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _333_ (.I(_175_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _334_ (.I(_160_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _335_ (.I(_176_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _336_ (.I(_176_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _337_ (.I(_176_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _338_ (.I(_176_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _339_ (.I(_176_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _340_ (.I(_176_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _341_ (.I(_176_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _342_ (.I(_176_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _343_ (.I(_176_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _344_ (.I(_176_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _345_ (.I(_160_),
    .Z(_177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _346_ (.I(_177_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _347_ (.I(_177_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _348_ (.I(_177_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _349_ (.I(_177_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _350_ (.I(_177_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _351_ (.I(_177_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _352_ (.I(_177_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _353_ (.I(_177_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _354_ (.I(_177_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _355_ (.I(_177_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _356_ (.D(net192),
    .RN(_000_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _357_ (.D(net268),
    .RN(_001_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _358_ (.D(net193),
    .RN(_002_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _359_ (.D(net275),
    .RN(_003_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _360_ (.D(net191),
    .RN(_004_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _361_ (.D(net255),
    .RN(_005_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _362_ (.D(net300),
    .RN(_006_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _363_ (.D(net1),
    .RN(_007_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _364_ (.D(net215),
    .RN(_008_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _365_ (.D(net224),
    .RN(_009_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _366_ (.D(net293),
    .RN(_010_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _367_ (.D(net279),
    .RN(_011_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _368_ (.D(net296),
    .RN(_012_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _369_ (.D(net299),
    .RN(_013_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _370_ (.D(net234),
    .RN(_014_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _371_ (.D(net298),
    .RN(_015_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _372_ (.D(net245),
    .RN(_016_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _373_ (.D(net232),
    .RN(_017_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _374_ (.D(net233),
    .RN(_018_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _375_ (.D(net178),
    .RN(_019_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _376_ (.D(net277),
    .RN(_020_),
    .CLK(clknet_4_3_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _377_ (.D(net195),
    .RN(_021_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _378_ (.D(net147),
    .RN(_022_),
    .CLK(clknet_4_1_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _379_ (.D(net276),
    .RN(_023_),
    .CLK(clknet_4_3_0_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _380_ (.D(net251),
    .RN(_024_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _381_ (.D(net206),
    .RN(_025_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _382_ (.D(net267),
    .RN(_026_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _383_ (.D(net212),
    .RN(_027_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _384_ (.D(net264),
    .RN(_028_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _385_ (.D(net202),
    .RN(_029_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _386_ (.D(net253),
    .RN(_030_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _387_ (.D(net177),
    .RN(_031_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _388_ (.D(net244),
    .RN(_032_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _389_ (.D(net153),
    .RN(_033_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _390_ (.D(net283),
    .RN(_034_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _391_ (.D(net252),
    .RN(_035_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _392_ (.D(net288),
    .RN(_036_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _393_ (.D(net289),
    .RN(_037_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _394_ (.D(net157),
    .RN(_038_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _395_ (.D(net301),
    .RN(_039_),
    .CLK(clknet_4_4_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _396_ (.D(net259),
    .RN(_040_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _397_ (.D(net146),
    .RN(_041_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _398_ (.D(net240),
    .RN(_042_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _399_ (.D(net238),
    .RN(_043_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _400_ (.D(net287),
    .RN(_044_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _401_ (.D(net261),
    .RN(_045_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _402_ (.D(net281),
    .RN(_046_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _403_ (.D(net220),
    .RN(_047_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _404_ (.D(net198),
    .RN(_048_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _405_ (.D(net179),
    .RN(_049_),
    .CLK(clknet_4_5_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _406_ (.D(net164),
    .RN(_050_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _407_ (.D(net272),
    .RN(_051_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _408_ (.D(net170),
    .RN(_052_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _409_ (.D(net171),
    .RN(_053_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _410_ (.D(net204),
    .RN(_054_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _411_ (.D(net216),
    .RN(_055_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _412_ (.D(net169),
    .RN(_056_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _413_ (.D(net174),
    .RN(_057_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _414_ (.D(net282),
    .RN(_058_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _415_ (.D(net260),
    .RN(_059_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _416_ (.D(net188),
    .RN(_060_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _417_ (.D(net219),
    .RN(_061_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _418_ (.D(net228),
    .RN(_062_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _419_ (.D(net256),
    .RN(_063_),
    .CLK(clknet_4_7_0_prog_clk),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _420_ (.D(net218),
    .RN(_064_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _421_ (.D(net151),
    .RN(_065_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _422_ (.D(net285),
    .RN(_066_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _423_ (.D(net148),
    .RN(_067_),
    .CLK(clknet_4_0_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _424_ (.D(net150),
    .RN(_068_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _425_ (.D(net295),
    .RN(_069_),
    .CLK(clknet_4_3_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _426_ (.D(net181),
    .RN(_070_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _427_ (.D(net246),
    .RN(_071_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _428_ (.D(net199),
    .RN(_072_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _429_ (.D(net250),
    .RN(_073_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _430_ (.D(net182),
    .RN(_074_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _431_ (.D(net225),
    .RN(_075_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _432_ (.D(net167),
    .RN(_076_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _433_ (.D(net165),
    .RN(_077_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _434_ (.D(net284),
    .RN(_078_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _435_ (.D(net209),
    .RN(_079_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _436_ (.D(net269),
    .RN(_080_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _437_ (.D(net221),
    .RN(_081_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _438_ (.D(net200),
    .RN(_082_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _439_ (.D(net162),
    .RN(_083_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _440_ (.D(net266),
    .RN(_084_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _441_ (.D(net213),
    .RN(_085_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _442_ (.D(net231),
    .RN(_086_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _443_ (.D(net210),
    .RN(_087_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _444_ (.D(net160),
    .RN(_088_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _445_ (.D(net294),
    .RN(_089_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _446_ (.D(net196),
    .RN(_090_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _447_ (.D(net243),
    .RN(_091_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _448_ (.D(net222),
    .RN(_092_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _449_ (.D(net205),
    .RN(_093_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _450_ (.D(net258),
    .RN(_094_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _451_ (.D(net197),
    .RN(_095_),
    .CLK(clknet_4_10_0_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _452_ (.D(net223),
    .RN(_096_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _453_ (.D(net203),
    .RN(_097_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _454_ (.D(net183),
    .RN(_098_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _455_ (.D(net173),
    .RN(_099_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _456_ (.D(net271),
    .RN(_100_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _457_ (.D(net227),
    .RN(_101_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _458_ (.D(net263),
    .RN(_102_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _459_ (.D(net175),
    .RN(_103_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _460_ (.D(net254),
    .RN(_104_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _461_ (.D(net149),
    .RN(_105_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _462_ (.D(net190),
    .RN(_106_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _463_ (.D(net280),
    .RN(_107_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _464_ (.D(net155),
    .RN(_108_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _465_ (.D(net297),
    .RN(_109_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _466_ (.D(net184),
    .RN(_110_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _467_ (.D(net186),
    .RN(_111_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _468_ (.D(net292),
    .RN(_112_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _469_ (.D(net286),
    .RN(_113_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _470_ (.D(net194),
    .RN(_114_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _471_ (.D(net235),
    .RN(_115_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _472_ (.D(net291),
    .RN(_116_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _473_ (.D(net262),
    .RN(_117_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _474_ (.D(net248),
    .RN(_118_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _475_ (.D(net214),
    .RN(_119_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_17.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _476_ (.D(net208),
    .RN(_120_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _477_ (.D(net145),
    .RN(_121_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _478_ (.D(net156),
    .RN(_122_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _479_ (.D(net189),
    .RN(_123_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _480_ (.D(net257),
    .RN(_124_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _481_ (.D(net237),
    .RN(_125_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _482_ (.D(net242),
    .RN(_126_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _483_ (.D(\mem_left_track_17.DFFR_7_.Q ),
    .RN(_127_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_left_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _484_ (.D(net226),
    .RN(_128_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _485_ (.D(net159),
    .RN(_129_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _486_ (.D(net211),
    .RN(_130_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _487_ (.D(net176),
    .RN(_131_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _488_ (.D(net163),
    .RN(_132_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _489_ (.D(net187),
    .RN(_133_),
    .CLK(clknet_4_3_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _490_ (.D(net249),
    .RN(_134_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _491_ (.D(net185),
    .RN(_135_),
    .CLK(clknet_4_6_0_prog_clk),
    .Q(\mem_top_track_32.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _492_ (.D(net161),
    .RN(_136_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _493_ (.D(net154),
    .RN(_137_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _494_ (.D(net273),
    .RN(_138_),
    .CLK(clknet_4_3_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _495_ (.D(net265),
    .RN(_139_),
    .CLK(clknet_4_2_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _496_ (.D(net158),
    .RN(_140_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _497_ (.D(net168),
    .RN(_141_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _498_ (.D(net239),
    .RN(_142_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _499_ (.D(net172),
    .RN(_143_),
    .CLK(clknet_4_12_0_prog_clk),
    .Q(\mem_right_track_32.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _500_ (.D(net166),
    .RN(_144_),
    .CLK(clknet_4_8_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _501_ (.D(net241),
    .RN(_145_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _502_ (.D(net247),
    .RN(_146_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _503_ (.D(net217),
    .RN(_147_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _504_ (.D(net230),
    .RN(_148_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _505_ (.D(net290),
    .RN(_149_),
    .CLK(clknet_4_9_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _506_ (.D(net207),
    .RN(_150_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _507_ (.D(net180),
    .RN(_151_),
    .CLK(clknet_4_11_0_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _508_ (.D(net152),
    .RN(_152_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _509_ (.D(net229),
    .RN(_153_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _510_ (.D(net201),
    .RN(_154_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _511_ (.D(net236),
    .RN(_155_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _512_ (.D(net270),
    .RN(_156_),
    .CLK(clknet_4_14_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _513_ (.D(net278),
    .RN(_157_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _514_ (.D(net144),
    .RN(_158_),
    .CLK(clknet_4_15_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _515_ (.D(net274),
    .RN(_159_),
    .CLK(clknet_4_13_0_prog_clk),
    .Q(\mem_left_track_33.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _536_ (.I(net24),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _537_ (.I(net23),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _538_ (.I(net22),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _539_ (.I(net21),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _540_ (.I(net20),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _541_ (.I(net19),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _542_ (.I(net18),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _543_ (.I(net31),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _544_ (.I(net30),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _545_ (.I(net29),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _546_ (.I(net28),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _547_ (.I(net27),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _548_ (.I(net26),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _549_ (.I(net25),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _550_ (.I(net17),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _551_ (.I(net9),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _552_ (.I(net8),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _553_ (.I(net7),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _554_ (.I(net6),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _555_ (.I(net5),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _556_ (.I(net4),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _557_ (.I(net3),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _558_ (.I(net16),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _559_ (.I(net15),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _560_ (.I(net14),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _561_ (.I(net13),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _562_ (.I(net12),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _563_ (.I(net11),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _564_ (.I(net10),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _565_ (.I(net2),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _566_ (.I(net54),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _567_ (.I(net53),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _568_ (.I(net52),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _569_ (.I(net51),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _570_ (.I(net50),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _571_ (.I(net49),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _572_ (.I(net48),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _573_ (.I(net61),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _574_ (.I(net60),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _575_ (.I(net59),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _576_ (.I(net58),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _577_ (.I(net57),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _578_ (.I(net56),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _579_ (.I(net55),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _580_ (.I(net47),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _581_ (.I(net39),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _582_ (.I(net38),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _583_ (.I(net37),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _584_ (.I(net36),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _585_ (.I(net35),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _586_ (.I(net34),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _587_ (.I(net33),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _588_ (.I(net46),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _589_ (.I(net45),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _590_ (.I(net44),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _591_ (.I(net43),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _592_ (.I(net42),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _593_ (.I(net41),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _594_ (.I(net40),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _595_ (.I(net32),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_0_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_10_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_11_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_12_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_13_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_14_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_15_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_1_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_2_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_3_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_4_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_5_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_6_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_7_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_8_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_4_9_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\mem_left_track_33.DFFR_0_.Q ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\mem_right_track_0.DFFR_5_.Q ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(\mem_bottom_track_25.DFFR_3_.Q ),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(\mem_right_track_0.DFFR_6_.Q ),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(\mem_top_track_16.DFFR_6_.Q ),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(\mem_bottom_track_1.DFFR_0_.D ),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(\mem_bottom_track_33.DFFR_4_.Q ),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(\mem_left_track_17.DFFR_0_.Q ),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(\mem_top_track_32.DFFR_0_.Q ),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(\mem_bottom_track_9.DFFR_5_.Q ),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold108 (.I(\mem_top_track_24.DFFR_6_.Q ),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(\mem_right_track_0.DFFR_3_.Q ),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\mem_right_track_32.DFFR_5_.Q ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold110 (.I(\mem_top_track_24.DFFR_0_.Q ),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold111 (.I(\mem_left_track_9.DFFR_6_.Q ),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold112 (.I(\mem_top_track_0.DFFR_1_.Q ),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold113 (.I(\mem_right_track_16.DFFR_7_.Q ),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold114 (.I(\mem_left_track_25.DFFR_2_.Q ),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold115 (.I(\mem_bottom_track_25.DFFR_0_.Q ),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold116 (.I(\mem_right_track_8.DFFR_6_.Q ),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold117 (.I(\mem_right_track_24.DFFR_3_.Q ),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold118 (.I(\mem_right_track_8.DFFR_1_.Q ),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold119 (.I(\mem_left_track_17.DFFR_1_.Q ),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\mem_left_track_9.DFFR_2_.Q ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold120 (.I(\mem_left_track_1.DFFR_0_.Q ),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold121 (.I(\mem_top_track_24.DFFR_2_.Q ),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold122 (.I(\mem_right_track_32.DFFR_3_.Q ),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold123 (.I(\mem_bottom_track_17.DFFR_2_.Q ),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold124 (.I(\mem_top_track_24.DFFR_4_.Q ),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold125 (.I(\mem_top_track_0.DFFR_5_.Q ),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold126 (.I(\mem_bottom_track_17.DFFR_6_.Q ),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold127 (.I(\mem_left_track_33.DFFR_2_.Q ),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold128 (.I(\mem_left_track_1.DFFR_2_.Q ),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold129 (.I(\mem_right_track_16.DFFR_3_.Q ),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\mem_left_track_25.DFFR_4_.Q ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold130 (.I(\mem_right_track_32.DFFR_4_.Q ),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold131 (.I(\mem_left_track_25.DFFR_7_.Q ),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold132 (.I(\mem_top_track_0.DFFR_3_.Q ),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold133 (.I(\mem_top_track_16.DFFR_0_.D ),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold134 (.I(\mem_top_track_16.DFFR_2_.Q ),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold135 (.I(\mem_left_track_33.DFFR_1_.Q ),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold136 (.I(\mem_top_track_8.DFFR_3_.Q ),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold137 (.I(\mem_left_track_9.DFFR_3_.Q ),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold138 (.I(\mem_right_track_8.DFFR_0_.Q ),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold139 (.I(\mem_right_track_24.DFFR_4_.Q ),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\mem_right_track_0.DFFR_0_.Q ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold140 (.I(\mem_right_track_0.DFFR_4_.Q ),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold141 (.I(\mem_bottom_track_9.DFFR_0_.Q ),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold142 (.I(\mem_bottom_track_1.DFFR_4_.Q ),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold143 (.I(\mem_left_track_17.DFFR_5_.Q ),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold144 (.I(\mem_right_track_8.DFFR_2_.Q ),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold145 (.I(\mem_right_track_0.DFFR_2_.Q ),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold146 (.I(\mem_right_track_0.DFFR_1_.Q ),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold147 (.I(\mem_bottom_track_33.DFFR_1_.Q ),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold148 (.I(\mem_left_track_17.DFFR_2_.Q ),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold149 (.I(\mem_left_track_17.DFFR_6_.Q ),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\mem_right_track_32.DFFR_2_.Q ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold150 (.I(\mem_top_track_8.DFFR_4_.Q ),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold151 (.I(\mem_bottom_track_25.DFFR_5_.Q ),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold152 (.I(\mem_bottom_track_1.DFFR_1_.Q ),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold153 (.I(\mem_top_track_8.DFFR_2_.Q ),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold154 (.I(\mem_left_track_9.DFFR_1_.Q ),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold155 (.I(\mem_top_track_0.DFFR_7_.Q ),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold156 (.I(\mem_top_track_8.DFFR_1_.Q ),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold157 (.I(\mem_top_track_0.DFFR_0_.Q ),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold158 (.I(\mem_right_track_0.DFFR_0_.D ),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\mem_top_track_32.DFFR_5_.Q ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\mem_bottom_track_25.DFFR_6_.Q ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\mem_right_track_32.DFFR_6_.Q ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\mem_bottom_track_17.DFFR_3_.Q ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\mem_left_track_25.DFFR_5_.Q ),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\mem_top_track_32.DFFR_2_.Q ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\mem_right_track_16.DFFR_4_.Q ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\mem_bottom_track_9.DFFR_1_.Q ),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\mem_bottom_track_33.DFFR_6_.Q ),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\mem_bottom_track_9.DFFR_2_.Q ),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\mem_right_track_32.DFFR_1_.Q ),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\mem_right_track_24.DFFR_6_.Q ),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\mem_right_track_16.DFFR_2_.Q ),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\mem_right_track_16.DFFR_1_.Q ),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\mem_right_track_24.DFFR_7_.Q ),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\mem_right_track_8.DFFR_5_.Q ),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\mem_left_track_1.DFFR_3_.Q ),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\mem_right_track_24.DFFR_5_.Q ),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\mem_bottom_track_33.DFFR_7_.Q ),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\mem_top_track_32.DFFR_3_.Q ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\mem_top_track_16.DFFR_7_.Q ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\mem_top_track_16.DFFR_3_.Q ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\mem_right_track_16.DFFR_5_.Q ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\mem_bottom_track_25.DFFR_7_.Q ),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\mem_bottom_track_1.DFFR_0_.Q ),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\mem_bottom_track_9.DFFR_4_.Q ),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\mem_top_track_16.DFFR_0_.Q ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\mem_left_track_1.DFFR_4_.Q ),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\mem_left_track_9.DFFR_0_.Q ),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\mem_top_track_24.DFFR_7_.Q ),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\mem_left_track_1.DFFR_7_.Q ),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\mem_top_track_32.DFFR_1_.Q ),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\mem_right_track_24.DFFR_2_.Q ),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\mem_left_track_25.DFFR_3_.Q ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\mem_left_track_9.DFFR_4_.Q ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(\mem_top_track_0.DFFR_2_.Q ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\mem_top_track_0.DFFR_6_.Q ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\mem_bottom_track_1.DFFR_3_.Q ),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(\mem_top_track_0.DFFR_4_.Q ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\mem_left_track_17.DFFR_4_.Q ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(\mem_top_track_16.DFFR_1_.Q ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\mem_bottom_track_25.DFFR_4_.Q ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(\mem_bottom_track_17.DFFR_7_.Q ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\mem_right_track_16.DFFR_6_.Q ),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(\mem_bottom_track_9.DFFR_6_.Q ),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\mem_bottom_track_17.DFFR_4_.Q ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(\mem_left_track_33.DFFR_4_.Q ),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\mem_top_track_24.DFFR_1_.Q ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\mem_left_track_9.DFFR_5_.Q ),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(\mem_left_track_1.DFFR_5_.Q ),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\mem_right_track_16.DFFR_0_.Q ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(\mem_bottom_track_25.DFFR_1_.Q ),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\mem_top_track_24.DFFR_5_.Q ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(\mem_bottom_track_33.DFFR_0_.Q ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\mem_left_track_25.DFFR_6_.Q ),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(\mem_bottom_track_1.DFFR_7_.Q ),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\mem_bottom_track_17.DFFR_0_.D ),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(\mem_top_track_32.DFFR_4_.Q ),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\mem_top_track_24.DFFR_3_.Q ),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\mem_bottom_track_1.DFFR_2_.Q ),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(\mem_bottom_track_17.DFFR_1_.Q ),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\mem_left_track_17.DFFR_0_.D ),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(\mem_top_track_8.DFFR_6_.Q ),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\mem_right_track_16.DFFR_0_.D ),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(\mem_bottom_track_33.DFFR_3_.Q ),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\mem_bottom_track_1.DFFR_6_.Q ),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(\mem_right_track_24.DFFR_1_.Q ),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\mem_right_track_0.DFFR_7_.Q ),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(\mem_bottom_track_17.DFFR_5_.Q ),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\mem_bottom_track_25.DFFR_2_.Q ),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\mem_bottom_track_1.DFFR_5_.Q ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(\mem_left_track_1.DFFR_6_.Q ),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\mem_top_track_8.DFFR_5_.Q ),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(\mem_bottom_track_9.DFFR_3_.Q ),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\mem_top_track_32.DFFR_6_.Q ),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(\mem_left_track_1.DFFR_1_.Q ),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\mem_right_track_24.DFFR_0_.Q ),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(\mem_left_track_33.DFFR_5_.Q ),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\mem_bottom_track_33.DFFR_2_.Q ),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(\mem_bottom_track_17.DFFR_0_.Q ),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\mem_top_track_16.DFFR_5_.Q ),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\mem_left_track_33.DFFR_6_.Q ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(\mem_top_track_16.DFFR_4_.Q ),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\mem_top_track_8.DFFR_0_.Q ),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(\mem_left_track_17.DFFR_3_.Q ),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\mem_left_track_33.DFFR_3_.Q ),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(\mem_left_track_25.DFFR_1_.Q ),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(\mem_right_track_8.DFFR_3_.Q ),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(\mem_right_track_32.DFFR_0_.Q ),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(\mem_right_track_8.DFFR_4_.Q ),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(\mem_bottom_track_33.DFFR_5_.Q ),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(\mem_left_track_25.DFFR_0_.Q ),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(chanx_left_in[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(chanx_left_in[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(chanx_left_in[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(chanx_left_in[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(chanx_left_in[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(chanx_left_in[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(chanx_left_in[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(chanx_right_in[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(chanx_right_in[10]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(chanx_right_in[12]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(chanx_left_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(chanx_right_in[13]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(chanx_right_in[14]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(chanx_right_in[16]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(chanx_right_in[17]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(chanx_right_in[18]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(chanx_right_in[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(chanx_right_in[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(chanx_right_in[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(chanx_right_in[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(chanx_right_in[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(chanx_left_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(chanx_right_in[8]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(chanx_right_in[9]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(chany_bottom_in[0]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(chany_bottom_in[10]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(chany_bottom_in[12]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(chany_bottom_in[13]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(chany_bottom_in[14]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(chany_bottom_in[16]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(chany_bottom_in[17]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(chany_bottom_in[18]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(chanx_left_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(chany_bottom_in[1]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(chany_bottom_in[2]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(chany_bottom_in[4]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(chany_bottom_in[5]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(chany_bottom_in[6]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(chany_bottom_in[8]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(chany_bottom_in[9]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(chany_top_in[0]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(chany_top_in[10]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(chany_top_in[12]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(chanx_left_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(chany_top_in[13]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(chany_top_in[14]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(chany_top_in[16]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(chany_top_in[17]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(chany_top_in[18]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(chany_top_in[1]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(chany_top_in[2]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(chany_top_in[4]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(chany_top_in[5]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(chany_top_in[6]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(chanx_left_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(chany_top_in[8]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(chany_top_in[9]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input62 (.I(pReset),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(chanx_left_in[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(chanx_left_in[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(chanx_left_in[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output100 (.I(net100),
    .Z(chany_bottom_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output101 (.I(net101),
    .Z(chany_bottom_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output102 (.I(net102),
    .Z(chany_bottom_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output103 (.I(net103),
    .Z(chany_bottom_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output104 (.I(net104),
    .Z(chany_bottom_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output105 (.I(net105),
    .Z(chany_bottom_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output106 (.I(net106),
    .Z(chany_bottom_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output107 (.I(net107),
    .Z(chany_bottom_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output108 (.I(net108),
    .Z(chany_bottom_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output109 (.I(net109),
    .Z(chany_top_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output110 (.I(net110),
    .Z(chany_top_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output111 (.I(net111),
    .Z(chany_top_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output112 (.I(net112),
    .Z(chany_top_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output113 (.I(net113),
    .Z(chany_top_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output114 (.I(net114),
    .Z(chany_top_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output115 (.I(net115),
    .Z(chany_top_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output116 (.I(net116),
    .Z(chany_top_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output117 (.I(net117),
    .Z(chany_top_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output118 (.I(net118),
    .Z(chany_top_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output119 (.I(net119),
    .Z(chany_top_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output120 (.I(net120),
    .Z(chany_top_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output121 (.I(net121),
    .Z(chany_top_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output122 (.I(net122),
    .Z(chany_top_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output123 (.I(net123),
    .Z(chany_top_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output63 (.I(net63),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output64 (.I(net64),
    .Z(chanx_left_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output65 (.I(net65),
    .Z(chanx_left_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output66 (.I(net66),
    .Z(chanx_left_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output67 (.I(net67),
    .Z(chanx_left_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(chanx_left_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output69 (.I(net69),
    .Z(chanx_left_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output70 (.I(net70),
    .Z(chanx_left_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output71 (.I(net71),
    .Z(chanx_left_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(chanx_left_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output73 (.I(net73),
    .Z(chanx_left_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output74 (.I(net74),
    .Z(chanx_left_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output75 (.I(net75),
    .Z(chanx_left_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output76 (.I(net76),
    .Z(chanx_left_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output77 (.I(net77),
    .Z(chanx_left_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output78 (.I(net78),
    .Z(chanx_left_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output79 (.I(net79),
    .Z(chanx_right_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output80 (.I(net80),
    .Z(chanx_right_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output81 (.I(net81),
    .Z(chanx_right_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output82 (.I(net82),
    .Z(chanx_right_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output83 (.I(net83),
    .Z(chanx_right_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output84 (.I(net84),
    .Z(chanx_right_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output85 (.I(net85),
    .Z(chanx_right_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output86 (.I(net86),
    .Z(chanx_right_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output87 (.I(net87),
    .Z(chanx_right_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output88 (.I(net88),
    .Z(chanx_right_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output89 (.I(net89),
    .Z(chanx_right_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output90 (.I(net90),
    .Z(chanx_right_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output91 (.I(net91),
    .Z(chanx_right_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output92 (.I(net92),
    .Z(chanx_right_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output93 (.I(net93),
    .Z(chanx_right_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output94 (.I(net94),
    .Z(chany_bottom_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output95 (.I(net95),
    .Z(chany_bottom_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output96 (.I(net96),
    .Z(chany_bottom_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output97 (.I(net97),
    .Z(chany_bottom_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output98 (.I(net98),
    .Z(chany_bottom_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output99 (.I(net99),
    .Z(chany_bottom_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__1__143 (.ZN(net143));
 assign chanx_left_out[0] = net143;
 assign chanx_left_out[12] = net140;
 assign chanx_left_out[16] = net139;
 assign chanx_left_out[4] = net142;
 assign chanx_left_out[8] = net141;
 assign chanx_right_out[0] = net138;
 assign chanx_right_out[12] = net135;
 assign chanx_right_out[16] = net134;
 assign chanx_right_out[4] = net137;
 assign chanx_right_out[8] = net136;
 assign chany_bottom_out[0] = net133;
 assign chany_bottom_out[12] = net130;
 assign chany_bottom_out[16] = net129;
 assign chany_bottom_out[4] = net132;
 assign chany_bottom_out[8] = net131;
 assign chany_top_out[0] = net128;
 assign chany_top_out[12] = net125;
 assign chany_top_out[16] = net124;
 assign chany_top_out[4] = net127;
 assign chany_top_out[8] = net126;
endmodule

