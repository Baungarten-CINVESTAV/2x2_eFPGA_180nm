magic
tech gf180mcuD
magscale 1 5
timestamp 1702148884
<< obsm1 >>
rect 672 1538 33320 32174
<< metal2 >>
rect 28224 33600 28280 34000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 20160 0 20216 400
rect 20496 0 20552 400
rect 21840 0 21896 400
rect 22176 0 22232 400
rect 24192 0 24248 400
rect 27216 0 27272 400
<< obsm2 >>
rect 854 33570 28194 33600
rect 28310 33570 33138 33600
rect 854 430 33138 33570
rect 854 400 978 430
rect 1094 400 1314 430
rect 1430 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2322 430
rect 2438 400 2658 430
rect 2774 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 4002 430
rect 4118 400 4338 430
rect 4454 400 4674 430
rect 4790 400 5010 430
rect 5126 400 20130 430
rect 20246 400 20466 430
rect 20582 400 21810 430
rect 21926 400 22146 430
rect 22262 400 24162 430
rect 24278 400 27186 430
rect 27302 400 33138 430
<< metal3 >>
rect 33600 31248 34000 31304
rect 0 23856 400 23912
rect 0 18144 400 18200
rect 33600 15456 34000 15512
rect 0 12432 400 12488
<< obsm3 >>
rect 400 31334 33600 32158
rect 400 31218 33570 31334
rect 400 23942 33600 31218
rect 430 23826 33600 23942
rect 400 18230 33600 23826
rect 430 18114 33600 18230
rect 400 15542 33600 18114
rect 400 15426 33570 15542
rect 400 12518 33600 15426
rect 430 12402 33600 12518
rect 400 1554 33600 12402
<< metal4 >>
rect 2224 1538 2384 32174
rect 9904 1538 10064 32174
rect 17584 1538 17744 32174
rect 25264 1538 25424 32174
rect 32944 1538 33104 32174
<< obsm4 >>
rect 20678 9865 25234 20151
rect 25454 9865 27034 20151
<< labels >>
rlabel metal2 s 0 0 56 400 6 bottom_width_0_height_0_subtile_0__pin_I_10_
port 1 nsew signal input
rlabel metal2 s 336 0 392 400 6 bottom_width_0_height_0_subtile_0__pin_I_2_
port 2 nsew signal input
rlabel metal2 s 672 0 728 400 6 bottom_width_0_height_0_subtile_0__pin_I_6_
port 3 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 bottom_width_0_height_0_subtile_0__pin_O_2_
port 4 nsew signal output
rlabel metal2 s 24192 0 24248 400 6 bottom_width_0_height_0_subtile_0__pin_O_6_
port 5 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 ccff_head
port 6 nsew signal input
rlabel metal3 s 33600 15456 34000 15512 6 ccff_tail
port 7 nsew signal output
rlabel metal2 s 1008 0 1064 400 6 clk
port 8 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 left_width_0_height_0_subtile_0__pin_I_11_
port 9 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 left_width_0_height_0_subtile_0__pin_I_3_
port 10 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 left_width_0_height_0_subtile_0__pin_I_7_
port 11 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 left_width_0_height_0_subtile_0__pin_O_3_
port 12 nsew signal output
rlabel metal3 s 33600 31248 34000 31304 6 left_width_0_height_0_subtile_0__pin_O_7_
port 13 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 pReset
port 14 nsew signal input
rlabel metal3 s 0 23856 400 23912 6 prog_clk
port 15 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 reset
port 16 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 right_width_0_height_0_subtile_0__pin_I_1_
port 17 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 right_width_0_height_0_subtile_0__pin_I_5_
port 18 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 right_width_0_height_0_subtile_0__pin_I_9_
port 19 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 right_width_0_height_0_subtile_0__pin_O_1_
port 20 nsew signal output
rlabel metal2 s 21840 0 21896 400 6 right_width_0_height_0_subtile_0__pin_O_5_
port 21 nsew signal output
rlabel metal2 s 3696 0 3752 400 6 set
port 22 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 top_width_0_height_0_subtile_0__pin_I_0_
port 23 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 top_width_0_height_0_subtile_0__pin_I_4_
port 24 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 top_width_0_height_0_subtile_0__pin_I_8_
port 25 nsew signal input
rlabel metal2 s 28224 33600 28280 34000 6 top_width_0_height_0_subtile_0__pin_O_0_
port 26 nsew signal output
rlabel metal2 s 22176 0 22232 400 6 top_width_0_height_0_subtile_0__pin_O_4_
port 27 nsew signal output
rlabel metal2 s 5040 0 5096 400 6 top_width_0_height_0_subtile_0__pin_clk_0_
port 28 nsew signal input
rlabel metal4 s 2224 1538 2384 32174 6 vdd
port 29 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 32174 6 vdd
port 29 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 32174 6 vdd
port 29 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 32174 6 vss
port 30 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 32174 6 vss
port 30 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 34000 34000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1489778
string GDS_FILE /home/baungarten/Desktop/2x2_FPGA_180nmD/openlane/grid_clb/runs/23_12_09_13_07/results/signoff/grid_clb.magic.gds
string GDS_START 99142
<< end >>

