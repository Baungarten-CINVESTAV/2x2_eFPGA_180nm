// This is the unpowered netlist.
module grid_clb (bottom_width_0_height_0_subtile_0__pin_I_10_,
    bottom_width_0_height_0_subtile_0__pin_I_2_,
    bottom_width_0_height_0_subtile_0__pin_I_6_,
    bottom_width_0_height_0_subtile_0__pin_O_2_,
    bottom_width_0_height_0_subtile_0__pin_O_6_,
    ccff_head,
    ccff_tail,
    clk,
    left_width_0_height_0_subtile_0__pin_I_11_,
    left_width_0_height_0_subtile_0__pin_I_3_,
    left_width_0_height_0_subtile_0__pin_I_7_,
    left_width_0_height_0_subtile_0__pin_O_3_,
    left_width_0_height_0_subtile_0__pin_O_7_,
    pReset,
    prog_clk,
    reset,
    right_width_0_height_0_subtile_0__pin_I_1_,
    right_width_0_height_0_subtile_0__pin_I_5_,
    right_width_0_height_0_subtile_0__pin_I_9_,
    right_width_0_height_0_subtile_0__pin_O_1_,
    right_width_0_height_0_subtile_0__pin_O_5_,
    set,
    top_width_0_height_0_subtile_0__pin_I_0_,
    top_width_0_height_0_subtile_0__pin_I_4_,
    top_width_0_height_0_subtile_0__pin_I_8_,
    top_width_0_height_0_subtile_0__pin_O_0_,
    top_width_0_height_0_subtile_0__pin_O_4_,
    top_width_0_height_0_subtile_0__pin_clk_0_);
 input bottom_width_0_height_0_subtile_0__pin_I_10_;
 input bottom_width_0_height_0_subtile_0__pin_I_2_;
 input bottom_width_0_height_0_subtile_0__pin_I_6_;
 output bottom_width_0_height_0_subtile_0__pin_O_2_;
 output bottom_width_0_height_0_subtile_0__pin_O_6_;
 input ccff_head;
 output ccff_tail;
 input clk;
 input left_width_0_height_0_subtile_0__pin_I_11_;
 input left_width_0_height_0_subtile_0__pin_I_3_;
 input left_width_0_height_0_subtile_0__pin_I_7_;
 output left_width_0_height_0_subtile_0__pin_O_3_;
 output left_width_0_height_0_subtile_0__pin_O_7_;
 input pReset;
 input prog_clk;
 input reset;
 input right_width_0_height_0_subtile_0__pin_I_1_;
 input right_width_0_height_0_subtile_0__pin_I_5_;
 input right_width_0_height_0_subtile_0__pin_I_9_;
 output right_width_0_height_0_subtile_0__pin_O_1_;
 output right_width_0_height_0_subtile_0__pin_O_5_;
 input set;
 input top_width_0_height_0_subtile_0__pin_I_0_;
 input top_width_0_height_0_subtile_0__pin_I_4_;
 input top_width_0_height_0_subtile_0__pin_I_8_;
 output top_width_0_height_0_subtile_0__pin_O_0_;
 output top_width_0_height_0_subtile_0__pin_O_4_;
 input top_width_0_height_0_subtile_0__pin_clk_0_;

 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire clknet_0_prog_clk;
 wire clknet_1_0__leaf_prog_clk;
 wire clknet_1_1__leaf_prog_clk;
 wire clknet_leaf_0_prog_clk;
 wire clknet_leaf_10_prog_clk;
 wire clknet_leaf_11_prog_clk;
 wire clknet_leaf_12_prog_clk;
 wire clknet_leaf_13_prog_clk;
 wire clknet_leaf_14_prog_clk;
 wire clknet_leaf_15_prog_clk;
 wire clknet_leaf_16_prog_clk;
 wire clknet_leaf_17_prog_clk;
 wire clknet_leaf_18_prog_clk;
 wire clknet_leaf_19_prog_clk;
 wire clknet_leaf_1_prog_clk;
 wire clknet_leaf_20_prog_clk;
 wire clknet_leaf_21_prog_clk;
 wire clknet_leaf_22_prog_clk;
 wire clknet_leaf_2_prog_clk;
 wire clknet_leaf_3_prog_clk;
 wire clknet_leaf_4_prog_clk;
 wire clknet_leaf_5_prog_clk;
 wire clknet_leaf_6_prog_clk;
 wire clknet_leaf_7_prog_clk;
 wire clknet_leaf_8_prog_clk;
 wire clknet_leaf_9_prog_clk;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_8_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_9_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_4_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_5_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_6_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_7_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_8_.Q ;
 wire net1;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__I (.I(_274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__I (.I(_276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__380__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__I (.I(_279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__I (.I(_272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__I (.I(_291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__I (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__552__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__563__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__I (.I(_265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__591__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__592__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__593__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__595__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__596__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__597__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__598__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__607__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__608__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__610__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__611__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__612__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__613__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__614__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__617__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__619__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__620__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__621__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__622__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__627__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__628__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__628__D (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__631__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__634__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__638__D (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__639__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__641__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__642__D (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__643__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__645__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__647__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__648__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__649__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__650__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__651__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__652__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__653__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__654__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__655__CLK (.I(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__657__CLK (.I(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__659__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__660__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__661__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__662__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__663__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__664__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__665__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__666__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__667__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__676__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__677__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__680__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__681__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__682__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__683__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__684__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__685__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__687__CLK (.I(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__728__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__729__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__730__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__731__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__732__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__733__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__CLK (.I(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__735__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__D (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__738__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__744__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__745__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__747__CLK (.I(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__748__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__751__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__765__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__766__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__768__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__769__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__770__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__771__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__772__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__773__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__774__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__775__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__776__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__777__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__778__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__779__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__780__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__782__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__783__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__784__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__785__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__786__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__787__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__788__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__789__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__790__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__791__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__792__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__793__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__794__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__795__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__797__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__798__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__800__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__803__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__804__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__805__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__809__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__810__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__813__CLK (.I(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__814__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__815__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__816__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__818__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__819__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__820__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__821__CLK (.I(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__822__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__823__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__825__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__826__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__827__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__829__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__830__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__831__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__835__CLK (.I(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__839__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__841__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__842__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__843__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__844__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__845__CLK (.I(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__847__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__848__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__849__CLK (.I(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__850__CLK (.I(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__850__D (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__851__CLK (.I(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_prog_clk_I (.I(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_prog_clk_I (.I(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold229_I (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold261_I (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _294_ (.I(_270_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _295_ (.I(_270_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _296_ (.I(_270_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _297_ (.I(_270_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _298_ (.I(_270_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _299_ (.I(_270_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _300_ (.I(_270_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _301_ (.I(_270_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _302_ (.I(_265_),
    .Z(_271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _303_ (.I(_271_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _304_ (.I(_271_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _305_ (.I(_271_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _306_ (.I(_271_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _307_ (.I(_271_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _308_ (.I(_271_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _309_ (.I(_271_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _310_ (.I(_271_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _311_ (.I(_271_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _312_ (.I(_271_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _313_ (.I(_264_),
    .Z(_272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _314_ (.I(_272_),
    .Z(_273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _315_ (.I(_273_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _316_ (.I(_273_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _317_ (.I(_273_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _318_ (.I(_273_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _319_ (.I(_273_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _320_ (.I(_273_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _321_ (.I(_273_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _322_ (.I(_273_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _323_ (.I(_273_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _324_ (.I(_273_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _325_ (.I(_272_),
    .Z(_274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _326_ (.I(_274_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _327_ (.I(_274_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _328_ (.I(_274_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _329_ (.I(_274_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _330_ (.I(_274_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _331_ (.I(_274_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _332_ (.I(_274_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _333_ (.I(_274_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _334_ (.I(_274_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _335_ (.I(_274_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _336_ (.I(_272_),
    .Z(_275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _337_ (.I(_275_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _338_ (.I(_275_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _339_ (.I(_275_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _340_ (.I(_275_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _341_ (.I(_275_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _342_ (.I(_275_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _343_ (.I(_275_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _344_ (.I(_275_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _345_ (.I(_275_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _346_ (.I(_275_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _347_ (.I(_272_),
    .Z(_276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _348_ (.I(_276_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _349_ (.I(_276_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _350_ (.I(_276_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _351_ (.I(_276_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _352_ (.I(_276_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _353_ (.I(_276_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _354_ (.I(_276_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _355_ (.I(_276_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _356_ (.I(_276_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _357_ (.I(_276_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _358_ (.I(_272_),
    .Z(_277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _359_ (.I(_277_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _360_ (.I(_277_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _361_ (.I(_277_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _362_ (.I(_277_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _363_ (.I(_277_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _364_ (.I(_277_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _365_ (.I(_277_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _366_ (.I(_277_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _367_ (.I(_277_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _368_ (.I(_277_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _369_ (.I(_272_),
    .Z(_278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _370_ (.I(_278_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _371_ (.I(_278_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _372_ (.I(_278_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _373_ (.I(_278_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _374_ (.I(_278_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _375_ (.I(_278_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _376_ (.I(_278_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _377_ (.I(_278_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _378_ (.I(_278_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _379_ (.I(_278_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _380_ (.I(_272_),
    .Z(_279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _381_ (.I(_279_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _382_ (.I(_279_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _383_ (.I(_279_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _384_ (.I(_279_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _385_ (.I(_279_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _386_ (.I(_279_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _387_ (.I(_279_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _388_ (.I(_279_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _389_ (.I(_279_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _390_ (.I(_279_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _391_ (.I(_272_),
    .Z(_280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _392_ (.I(_280_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _393_ (.I(_280_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _394_ (.I(_280_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _395_ (.I(_280_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _396_ (.I(_280_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _397_ (.I(_280_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _398_ (.I(_280_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _399_ (.I(_280_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _400_ (.I(_280_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _401_ (.I(_280_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _402_ (.I(_272_),
    .Z(_281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _403_ (.I(_281_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _404_ (.I(_281_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _405_ (.I(_281_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _406_ (.I(_281_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _407_ (.I(_281_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _408_ (.I(_281_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _409_ (.I(_281_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _410_ (.I(_281_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _411_ (.I(_281_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _412_ (.I(_281_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _413_ (.I(_272_),
    .Z(_282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _414_ (.I(_282_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _415_ (.I(_282_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _416_ (.I(_282_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _417_ (.I(_282_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _418_ (.I(_282_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _419_ (.I(_282_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _420_ (.I(_282_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _421_ (.I(_282_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _422_ (.I(_282_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _423_ (.I(_282_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _424_ (.I(_264_),
    .Z(_283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _425_ (.I(_283_),
    .Z(_284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _426_ (.I(_284_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _427_ (.I(_284_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _428_ (.I(_284_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _429_ (.I(_284_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _430_ (.I(_284_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _431_ (.I(_284_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _432_ (.I(_284_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _433_ (.I(_284_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _434_ (.I(_284_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _435_ (.I(_284_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _436_ (.I(_283_),
    .Z(_285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _437_ (.I(_285_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _438_ (.I(_285_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _439_ (.I(_285_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _440_ (.I(_285_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _441_ (.I(_285_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _442_ (.I(_285_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _443_ (.I(_285_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _444_ (.I(_285_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _445_ (.I(_285_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _446_ (.I(_285_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _447_ (.I(_283_),
    .Z(_286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _448_ (.I(_286_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _449_ (.I(_286_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _450_ (.I(_286_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _451_ (.I(_286_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _452_ (.I(_286_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _453_ (.I(_286_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _454_ (.I(_286_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _455_ (.I(_286_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _456_ (.I(_286_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _457_ (.I(_286_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _458_ (.I(_283_),
    .Z(_287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _459_ (.I(_287_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _460_ (.I(_287_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _461_ (.I(_287_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _462_ (.I(_287_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _463_ (.I(_287_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _464_ (.I(_287_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _465_ (.I(_287_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _466_ (.I(_287_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _467_ (.I(_287_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _468_ (.I(_287_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _469_ (.I(_283_),
    .Z(_288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _470_ (.I(_288_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _471_ (.I(_288_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _472_ (.I(_288_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _473_ (.I(_288_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _474_ (.I(_288_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _475_ (.I(_288_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _476_ (.I(_288_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _477_ (.I(_288_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _478_ (.I(_288_),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _479_ (.I(_288_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _480_ (.I(_283_),
    .Z(_289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _481_ (.I(_289_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _482_ (.I(_289_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _483_ (.I(_289_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _484_ (.I(_289_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _485_ (.I(_289_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _486_ (.I(_289_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _487_ (.I(_289_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _488_ (.I(_289_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _489_ (.I(_289_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _490_ (.I(_289_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _491_ (.I(_283_),
    .Z(_290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _492_ (.I(_290_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _493_ (.I(_290_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _494_ (.I(_290_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _495_ (.I(_290_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _496_ (.I(_290_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _497_ (.I(_290_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _498_ (.I(_290_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _499_ (.I(_290_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _500_ (.I(_290_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _501_ (.I(_290_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _502_ (.I(_283_),
    .Z(_291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _503_ (.I(_291_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _504_ (.I(_291_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _505_ (.I(_291_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _506_ (.I(_291_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _507_ (.I(_291_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _508_ (.I(_291_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _509_ (.I(_291_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _510_ (.I(_291_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _511_ (.I(_291_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _512_ (.I(_291_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _513_ (.I(_283_),
    .Z(_292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _514_ (.I(_292_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _515_ (.I(_292_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _516_ (.I(_292_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _517_ (.I(_292_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _518_ (.I(_292_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _519_ (.I(_292_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _520_ (.I(_292_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _521_ (.I(_292_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _522_ (.I(_292_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _523_ (.I(_292_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _524_ (.I(_283_),
    .Z(_293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _525_ (.I(_293_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _526_ (.I(_293_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _527_ (.I(_293_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _528_ (.I(_293_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _529_ (.I(_293_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _530_ (.I(_293_),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _531_ (.I(_293_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _532_ (.I(_293_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _533_ (.I(_293_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _534_ (.I(_293_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _535_ (.I(_265_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _536_ (.I(_265_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _537_ (.I(_265_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _538_ (.I(_265_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _539_ (.I(net2),
    .Z(_264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _540_ (.I(_264_),
    .Z(_265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _541_ (.I(_265_),
    .Z(_266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _542_ (.I(_266_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _543_ (.I(_266_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _544_ (.I(_266_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _545_ (.I(_266_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _546_ (.I(_266_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _547_ (.I(_266_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _548_ (.I(_266_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _549_ (.I(_266_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _550_ (.I(_266_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _551_ (.I(_266_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _552_ (.I(_265_),
    .Z(_267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _553_ (.I(_267_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _554_ (.I(_267_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _555_ (.I(_267_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _556_ (.I(_267_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _557_ (.I(_267_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _558_ (.I(_267_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _559_ (.I(_267_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _560_ (.I(_267_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _561_ (.I(_267_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _562_ (.I(_267_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _563_ (.I(_265_),
    .Z(_268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _564_ (.I(_268_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _565_ (.I(_268_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _566_ (.I(_268_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _567_ (.I(_268_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _568_ (.I(_268_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _569_ (.I(_268_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _570_ (.I(_268_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _571_ (.I(_268_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _572_ (.I(_268_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _573_ (.I(_268_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _574_ (.I(_265_),
    .Z(_269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _575_ (.I(_269_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _576_ (.I(_269_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _577_ (.I(_269_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _578_ (.I(_269_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _579_ (.I(_269_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _580_ (.I(_269_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _581_ (.I(_269_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _582_ (.I(_269_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _583_ (.I(_269_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _584_ (.I(_269_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _585_ (.I(_265_),
    .Z(_270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _586_ (.I(_270_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _587_ (.I(_270_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _588_ (.D(net235),
    .RN(_000_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _589_ (.D(net250),
    .RN(_001_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _590_ (.D(net42),
    .RN(_002_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _591_ (.D(net207),
    .RN(_003_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _592_ (.D(net78),
    .RN(_004_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _593_ (.D(net59),
    .RN(_005_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _594_ (.D(net85),
    .RN(_006_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _595_ (.D(net177),
    .RN(_007_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _596_ (.D(net135),
    .RN(_008_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _597_ (.D(net153),
    .RN(_009_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _598_ (.D(net121),
    .RN(_010_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _599_ (.D(net56),
    .RN(_011_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _600_ (.D(net148),
    .RN(_012_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _601_ (.D(net166),
    .RN(_013_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _602_ (.D(net129),
    .RN(_014_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _603_ (.D(net203),
    .RN(_015_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _604_ (.D(net156),
    .RN(_016_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _605_ (.D(net239),
    .RN(_017_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _606_ (.D(net241),
    .RN(_018_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _607_ (.D(net69),
    .RN(_019_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _608_ (.D(net35),
    .RN(_020_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _609_ (.D(net84),
    .RN(_021_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _610_ (.D(net72),
    .RN(_022_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _611_ (.D(net221),
    .RN(_023_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _612_ (.D(net115),
    .RN(_024_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _613_ (.D(net172),
    .RN(_025_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _614_ (.D(net259),
    .RN(_026_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _615_ (.D(net66),
    .RN(_027_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _616_ (.D(net169),
    .RN(_028_),
    .CLK(clknet_leaf_15_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _617_ (.D(net79),
    .RN(_029_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _618_ (.D(net193),
    .RN(_030_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _619_ (.D(net51),
    .RN(_031_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _620_ (.D(net159),
    .RN(_032_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _621_ (.D(net191),
    .RN(_033_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _622_ (.D(net141),
    .RN(_034_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _623_ (.D(net95),
    .RN(_035_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _624_ (.D(net81),
    .RN(_036_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _625_ (.D(net171),
    .RN(_037_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _626_ (.D(net64),
    .RN(_038_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _627_ (.D(net62),
    .RN(_039_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _628_ (.D(net274),
    .RN(_040_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _629_ (.D(net15),
    .RN(_041_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _630_ (.D(net76),
    .RN(_042_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _631_ (.D(net87),
    .RN(_043_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _632_ (.D(net154),
    .RN(_044_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _633_ (.D(net17),
    .RN(_045_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _634_ (.D(net103),
    .RN(_046_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _635_ (.D(net12),
    .RN(_047_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _636_ (.D(net236),
    .RN(_048_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _637_ (.D(net238),
    .RN(_049_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _638_ (.D(net271),
    .RN(_050_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _639_ (.D(net25),
    .RN(_051_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _640_ (.D(net212),
    .RN(_052_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _641_ (.D(net30),
    .RN(_053_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _642_ (.D(net249),
    .RN(_054_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _643_ (.D(net27),
    .RN(_055_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _644_ (.D(net102),
    .RN(_056_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _645_ (.D(net28),
    .RN(_057_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _646_ (.D(net198),
    .RN(_058_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _647_ (.D(net140),
    .RN(_059_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _648_ (.D(net110),
    .RN(_060_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _649_ (.D(net65),
    .RN(_061_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _650_ (.D(net86),
    .RN(_062_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _651_ (.D(net126),
    .RN(_063_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _652_ (.D(net165),
    .RN(_064_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _653_ (.D(net63),
    .RN(_065_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _654_ (.D(net83),
    .RN(_066_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _655_ (.D(net33),
    .RN(_067_),
    .CLK(clknet_leaf_13_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _656_ (.D(net94),
    .RN(_068_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _657_ (.D(net70),
    .RN(_069_),
    .CLK(clknet_leaf_14_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _658_ (.D(net151),
    .RN(_070_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _659_ (.D(net40),
    .RN(_071_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _660_ (.D(net118),
    .RN(_072_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _661_ (.D(net112),
    .RN(_073_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _662_ (.D(net107),
    .RN(_074_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _663_ (.D(net125),
    .RN(_075_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _664_ (.D(net138),
    .RN(_076_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _665_ (.D(net77),
    .RN(_077_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _666_ (.D(net99),
    .RN(_078_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _667_ (.D(net152),
    .RN(_079_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _668_ (.D(net269),
    .RN(_080_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _669_ (.D(net80),
    .RN(_081_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _670_ (.D(net186),
    .RN(_082_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _671_ (.D(net82),
    .RN(_083_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _672_ (.D(net174),
    .RN(_084_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _673_ (.D(net247),
    .RN(_085_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _674_ (.D(net98),
    .RN(_086_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _675_ (.D(net45),
    .RN(_087_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _676_ (.D(net52),
    .RN(_088_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _677_ (.D(net227),
    .RN(_089_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _678_ (.D(net37),
    .RN(_090_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _679_ (.D(net96),
    .RN(_091_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _680_ (.D(net36),
    .RN(_092_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _681_ (.D(net202),
    .RN(_093_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _682_ (.D(net137),
    .RN(_094_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _683_ (.D(net131),
    .RN(_095_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _684_ (.D(net136),
    .RN(_096_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _685_ (.D(net104),
    .RN(_097_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _686_ (.D(net100),
    .RN(_098_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _687_ (.D(net44),
    .RN(_099_),
    .CLK(clknet_leaf_9_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _688_ (.D(net68),
    .RN(_100_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _689_ (.D(net157),
    .RN(_101_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _690_ (.D(net180),
    .RN(_102_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _691_ (.D(net189),
    .RN(_103_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _692_ (.D(net187),
    .RN(_104_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _693_ (.D(net251),
    .RN(_105_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _694_ (.D(net90),
    .RN(_106_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _695_ (.D(net71),
    .RN(_107_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _696_ (.D(net60),
    .RN(_108_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _697_ (.D(net245),
    .RN(_109_),
    .CLK(clknet_leaf_8_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _698_ (.D(net231),
    .RN(_110_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _699_ (.D(net24),
    .RN(_111_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _700_ (.D(net49),
    .RN(_112_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _701_ (.D(net237),
    .RN(_113_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _702_ (.D(net192),
    .RN(_114_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _703_ (.D(net185),
    .RN(_115_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _704_ (.D(net23),
    .RN(_116_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _705_ (.D(net216),
    .RN(_117_),
    .CLK(clknet_leaf_7_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _706_ (.D(net58),
    .RN(_118_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _707_ (.D(net123),
    .RN(_119_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _708_ (.D(net196),
    .RN(_120_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _709_ (.D(net145),
    .RN(_121_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _710_ (.D(net144),
    .RN(_122_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _711_ (.D(net142),
    .RN(_123_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _712_ (.D(net266),
    .RN(_124_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _713_ (.D(net120),
    .RN(_125_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _714_ (.D(net262),
    .RN(_126_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _715_ (.D(net119),
    .RN(_127_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _716_ (.D(net214),
    .RN(_128_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _717_ (.D(net209),
    .RN(_129_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _718_ (.D(net264),
    .RN(_130_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _719_ (.D(net205),
    .RN(_131_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _720_ (.D(net113),
    .RN(_132_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _721_ (.D(net179),
    .RN(_133_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _722_ (.D(net273),
    .RN(_134_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _723_ (.D(net38),
    .RN(_135_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _724_ (.D(net22),
    .RN(_136_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _725_ (.D(net181),
    .RN(_137_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _726_ (.D(net167),
    .RN(_138_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _727_ (.D(net176),
    .RN(_139_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _728_ (.D(net132),
    .RN(_140_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _729_ (.D(net225),
    .RN(_141_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _730_ (.D(net228),
    .RN(_142_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _731_ (.D(net208),
    .RN(_143_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _732_ (.D(net204),
    .RN(_144_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _733_ (.D(net160),
    .RN(_145_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _734_ (.D(net93),
    .RN(_146_),
    .CLK(clknet_leaf_10_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _735_ (.D(net54),
    .RN(_147_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _736_ (.D(net89),
    .RN(_148_),
    .CLK(clknet_leaf_6_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _737_ (.D(net57),
    .RN(_149_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _738_ (.D(net184),
    .RN(_150_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _739_ (.D(net14),
    .RN(_151_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _740_ (.D(net252),
    .RN(_152_),
    .CLK(clknet_leaf_12_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _741_ (.D(net61),
    .RN(_153_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _742_ (.D(net232),
    .RN(_154_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _743_ (.D(net130),
    .RN(_155_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _744_ (.D(net16),
    .RN(_156_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _745_ (.D(net162),
    .RN(_157_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _746_ (.D(net147),
    .RN(_158_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_8_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _747_ (.D(net13),
    .RN(_159_),
    .CLK(clknet_leaf_11_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_9_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _748_ (.D(net260),
    .RN(_160_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _749_ (.D(net46),
    .RN(_161_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _750_ (.D(net195),
    .RN(_162_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _751_ (.D(net161),
    .RN(_163_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _752_ (.D(net158),
    .RN(_164_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _753_ (.D(net168),
    .RN(_165_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _754_ (.D(net210),
    .RN(_166_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _755_ (.D(net248),
    .RN(_167_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _756_ (.D(net173),
    .RN(_168_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _757_ (.D(net139),
    .RN(_169_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _758_ (.D(net149),
    .RN(_170_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _759_ (.D(net234),
    .RN(_171_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _760_ (.D(net31),
    .RN(_172_),
    .CLK(clknet_leaf_4_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _761_ (.D(net92),
    .RN(_173_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _762_ (.D(net199),
    .RN(_174_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _763_ (.D(net188),
    .RN(_175_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _764_ (.D(net109),
    .RN(_176_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _765_ (.D(net267),
    .RN(_177_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _766_ (.D(net194),
    .RN(_178_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _767_ (.D(net29),
    .RN(_179_),
    .CLK(clknet_leaf_5_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _768_ (.D(net32),
    .RN(_180_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _769_ (.D(net261),
    .RN(_181_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _770_ (.D(net243),
    .RN(_182_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _771_ (.D(net254),
    .RN(_183_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _772_ (.D(net163),
    .RN(_184_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _773_ (.D(net201),
    .RN(_185_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _774_ (.D(net197),
    .RN(_186_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _775_ (.D(net211),
    .RN(_187_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _776_ (.D(net183),
    .RN(_188_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _777_ (.D(net175),
    .RN(_189_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _778_ (.D(net240),
    .RN(_190_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _779_ (.D(net182),
    .RN(_191_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _780_ (.D(net164),
    .RN(_192_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _781_ (.D(net88),
    .RN(_193_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _782_ (.D(net108),
    .RN(_194_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _783_ (.D(net257),
    .RN(_195_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _784_ (.D(net215),
    .RN(_196_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _785_ (.D(net244),
    .RN(_197_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _786_ (.D(net255),
    .RN(_198_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _787_ (.D(net206),
    .RN(_199_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _788_ (.D(net117),
    .RN(_200_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _789_ (.D(net48),
    .RN(_201_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _790_ (.D(net116),
    .RN(_202_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _791_ (.D(net106),
    .RN(_203_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _792_ (.D(net230),
    .RN(_204_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _793_ (.D(net128),
    .RN(_205_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _794_ (.D(net73),
    .RN(_206_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _795_ (.D(net34),
    .RN(_207_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _796_ (.D(net233),
    .RN(_208_),
    .CLK(clknet_leaf_3_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _797_ (.D(net272),
    .RN(_209_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _798_ (.D(net222),
    .RN(_210_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _799_ (.D(net18),
    .RN(_211_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _800_ (.D(net213),
    .RN(_212_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _801_ (.D(net20),
    .RN(_213_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _802_ (.D(net67),
    .RN(_214_),
    .CLK(clknet_leaf_18_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _803_ (.D(net134),
    .RN(_215_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _804_ (.D(net242),
    .RN(_216_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _805_ (.D(net219),
    .RN(_217_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _806_ (.D(net19),
    .RN(_218_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _807_ (.D(net155),
    .RN(_219_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _808_ (.D(net253),
    .RN(_220_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _809_ (.D(net41),
    .RN(_221_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _810_ (.D(net170),
    .RN(_222_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _811_ (.D(net111),
    .RN(_223_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _812_ (.D(net220),
    .RN(_224_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _813_ (.D(net55),
    .RN(_225_),
    .CLK(clknet_leaf_16_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _814_ (.D(net265),
    .RN(_226_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _815_ (.D(net97),
    .RN(_227_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _816_ (.D(net47),
    .RN(_228_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _817_ (.D(net21),
    .RN(_229_),
    .CLK(clknet_leaf_17_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _818_ (.D(net200),
    .RN(_230_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _819_ (.D(net133),
    .RN(_231_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _820_ (.D(net263),
    .RN(_232_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _821_ (.D(net114),
    .RN(_233_),
    .CLK(clknet_leaf_19_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _822_ (.D(net143),
    .RN(_234_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _823_ (.D(net256),
    .RN(_235_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _824_ (.D(net146),
    .RN(_236_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _825_ (.D(net50),
    .RN(_237_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _826_ (.D(net224),
    .RN(_238_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _827_ (.D(net39),
    .RN(_239_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _828_ (.D(net268),
    .RN(_240_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _829_ (.D(net1),
    .RN(_241_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _830_ (.D(net105),
    .RN(_242_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _831_ (.D(net246),
    .RN(_243_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _832_ (.D(net91),
    .RN(_244_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _833_ (.D(net270),
    .RN(_245_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _834_ (.D(net226),
    .RN(_246_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _835_ (.D(net53),
    .RN(_247_),
    .CLK(clknet_leaf_0_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _836_ (.D(net101),
    .RN(_248_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _837_ (.D(net124),
    .RN(_249_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _838_ (.D(net150),
    .RN(_250_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _839_ (.D(net75),
    .RN(_251_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _840_ (.D(net43),
    .RN(_252_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _841_ (.D(net74),
    .RN(_253_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _842_ (.D(net218),
    .RN(_254_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _843_ (.D(net127),
    .RN(_255_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _844_ (.D(net229),
    .RN(_256_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _845_ (.D(net223),
    .RN(_257_),
    .CLK(clknet_leaf_21_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _846_ (.D(net178),
    .RN(_258_),
    .CLK(clknet_leaf_22_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _847_ (.D(net217),
    .RN(_259_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _848_ (.D(net190),
    .RN(_260_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _849_ (.D(net122),
    .RN(_261_),
    .CLK(clknet_leaf_20_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _850_ (.D(net26),
    .RN(_262_),
    .CLK(clknet_leaf_1_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _851_ (.D(net258),
    .RN(_263_),
    .CLK(clknet_leaf_2_prog_clk),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_1_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_1_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_10_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_11_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_12_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_13_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_14_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_15_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_16_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_17_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_18_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_19_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_1_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_20_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_21_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_22_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_2_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_3_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_4_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_prog_clk (.I(clknet_1_0__leaf_prog_clk),
    .Z(clknet_leaf_5_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_6_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_7_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_8_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_prog_clk (.I(clknet_1_1__leaf_prog_clk),
    .Z(clknet_leaf_9_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_10 (.ZN(net10));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_11 (.ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_4 (.ZN(net4));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_5 (.ZN(net5));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_6 (.ZN(net6));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_7 (.ZN(net7));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_8 (.ZN(net8));
 gf180mcu_fd_sc_mcu7t5v0__tiel grid_clb_9 (.ZN(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_6_.Q ),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_2_.Q ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_1_.Q ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_3_.Q ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_1_.Q ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold108 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_6_.Q ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_4_.Q ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_5_.Q ),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold110 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_9_.Q ),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold111 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold112 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_8_.Q ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold113 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold114 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_4_.Q ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold115 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_2_.Q ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold116 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold117 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold118 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_3_.Q ),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold119 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_4_.Q ),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_5_.Q ),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold120 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_4_.Q ),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold121 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_9_.Q ),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold122 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold123 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold124 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_7_.Q ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold125 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_5_.Q ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold126 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_3_.Q ),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold127 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_5_.Q ),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold128 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold129 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_8_.Q ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_0_.Q ),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold130 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_3_.Q ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold131 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_2_.Q ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold132 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold133 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_1_.Q ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold134 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_0_.Q ),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold135 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold136 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_7_.Q ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold137 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_1_.Q ),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold138 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold139 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_0_.Q ),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold140 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_9_.Q ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold141 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_8_.Q ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold142 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_8_.Q ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold143 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_3_.Q ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold144 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold145 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_5_.Q ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold146 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_0_.Q ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold147 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold148 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_1_.Q ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold149 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_4_.Q ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold150 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold151 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_6_.Q ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold152 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold153 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold154 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_3_.Q ),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold155 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_2_.Q ),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold156 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_7_.Q ),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold157 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold158 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_7_.Q ),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold159 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_4_.Q ),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold160 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_6_.Q ),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold161 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_4_.Q ),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold162 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold163 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_3_.Q ),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold164 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold165 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_8_.Q ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold166 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_6_.Q ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold167 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold168 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_2_.Q ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold169 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_1_.Q ),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_6_.Q ),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold170 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_6_.Q ),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold171 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold172 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold173 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold174 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_4_.Q ),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold175 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_1_.Q ),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold176 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_3_.Q ),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold177 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold178 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_2_.Q ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold179 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold180 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_2_.Q ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold181 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_3_.Q ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold182 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_9_.Q ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold183 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold184 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold185 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_9_.Q ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold186 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold187 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_7_.Q ),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold188 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold189 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_2_.Q ),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold190 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold191 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_2_.Q ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold192 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_4_.Q ),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold193 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_3_.Q ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold194 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_0_.Q ),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold195 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold196 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_2_.Q ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold197 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_2_.Q ),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold198 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_8_.Q ),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold199 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_8_.Q ),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold200 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold201 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_1_.Q ),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold202 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold203 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_7_.Q ),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold204 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold205 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_6_.Q ),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold206 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold207 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold208 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold209 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold210 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_2_.Q ),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold211 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold212 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_15_.in ),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold213 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold214 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_0_.Q ),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold215 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold216 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_8_.Q ),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold217 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_1_.Q ),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold218 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold219 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_14_.in ),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_6_.Q ),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold220 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_9_.Q ),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold221 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_3_.Q ),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold222 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold223 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold224 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_9_.Q ),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold225 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_7_.Q ),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold226 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_2_.Q ),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold227 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_8_.Q ),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold228 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_6_.Q ),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold229 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold230 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_7_.Q ),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold231 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold232 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_0_.Q ),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold233 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_7_.in ),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold234 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_8_.Q ),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold235 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_1_.in ),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold236 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_4_.Q ),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold237 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold238 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_3_.Q ),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold239 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_0_.Q ),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_9_.Q ),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold240 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_4_.Q ),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold241 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_1_.Q ),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold242 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold243 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold244 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_8_.in ),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold245 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold246 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold247 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_0_.Q ),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold248 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_5_.Q ),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold249 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail ),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_1_.Q ),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold250 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.DFFR_1_.Q ),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold251 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_5_.Q ),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold252 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold253 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_9_.Q ),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold254 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold255 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFFR_3_.Q ),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold256 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold257 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold258 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_9_.Q ),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold259 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_9_.Q ),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold260 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_9_.Q ),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold261 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_2_.Q ),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold262 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_3_.Q ),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold263 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_9_.Q ),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFFR_4_.Q ),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_0_.Q ),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_0_.Q ),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_1_.Q ),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_10_.in ),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_8_.Q ),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_6_.Q ),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_1_.Q ),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_0_.Q ),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_0_.Q ),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_7_.Q ),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_5_.in ),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_6_.Q ),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_0_.Q ),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_8_.Q ),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_7_.Q ),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_4_.Q ),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_7_.Q ),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_5_.Q ),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFFR_2_.Q ),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_8_.Q ),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_4_.Q ),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_7_.Q ),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_0_.Q ),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_6_.Q ),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_1_.Q ),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFFR_9_.Q ),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFFR_8_.Q ),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_8_.Q ),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_4_.Q ),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_6_.Q ),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_1_.Q ),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail ),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_1_.Q ),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_6_.Q ),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_3_.Q ),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_8_.Q ),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_0_.Q ),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.DFFR_1_.Q ),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_5_.Q ),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_2_.Q ),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_5_.Q ),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFFR_0_.Q ),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFFR_5_.Q ),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_1_.Q ),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_2_.Q ),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_3_.in ),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_7_.Q ),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFFR_5_.Q ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_2_.in ),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_9_.in ),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFFR_5_.Q ),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFFR_7_.Q ),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFFR_4_.Q ),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_0_.Q ),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_11_.in ),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFFR_5_.Q ),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_7_.Q ),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_7_.Q ),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.DFFR_0_.Q ),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_6_.in ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFFR_5_.Q ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFFR_5_.Q ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFFR_6_.Q ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_0_.in ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_13_.in ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_3_.Q ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_4_.in ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.INVTX1_12_.in ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFFR_9_.Q ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(pReset),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output3 (.I(net3),
    .Z(ccff_tail));
 assign bottom_width_0_height_0_subtile_0__pin_O_2_ = net7;
 assign bottom_width_0_height_0_subtile_0__pin_O_6_ = net6;
 assign left_width_0_height_0_subtile_0__pin_O_3_ = net5;
 assign left_width_0_height_0_subtile_0__pin_O_7_ = net4;
 assign right_width_0_height_0_subtile_0__pin_O_1_ = net8;
 assign right_width_0_height_0_subtile_0__pin_O_5_ = net9;
 assign top_width_0_height_0_subtile_0__pin_O_0_ = net10;
 assign top_width_0_height_0_subtile_0__pin_O_4_ = net11;
endmodule

