magic
tech gf180mcuD
magscale 1 5
timestamp 1702157087
<< metal1 >>
rect 672 6285 7360 6302
rect 672 6259 2259 6285
rect 2285 6259 2311 6285
rect 2337 6259 2363 6285
rect 2389 6259 3911 6285
rect 3937 6259 3963 6285
rect 3989 6259 4015 6285
rect 4041 6259 5563 6285
rect 5589 6259 5615 6285
rect 5641 6259 5667 6285
rect 5693 6259 7215 6285
rect 7241 6259 7267 6285
rect 7293 6259 7319 6285
rect 7345 6259 7360 6285
rect 672 6242 7360 6259
rect 672 5893 7280 5910
rect 672 5867 1433 5893
rect 1459 5867 1485 5893
rect 1511 5867 1537 5893
rect 1563 5867 3085 5893
rect 3111 5867 3137 5893
rect 3163 5867 3189 5893
rect 3215 5867 4737 5893
rect 4763 5867 4789 5893
rect 4815 5867 4841 5893
rect 4867 5867 6389 5893
rect 6415 5867 6441 5893
rect 6467 5867 6493 5893
rect 6519 5867 7280 5893
rect 672 5850 7280 5867
rect 3543 5697 3569 5703
rect 3761 5671 3767 5697
rect 3793 5671 3799 5697
rect 3543 5665 3569 5671
rect 5279 5585 5305 5591
rect 4881 5559 4887 5585
rect 4913 5559 4919 5585
rect 5279 5553 5305 5559
rect 672 5501 7360 5518
rect 672 5475 2259 5501
rect 2285 5475 2311 5501
rect 2337 5475 2363 5501
rect 2389 5475 3911 5501
rect 3937 5475 3963 5501
rect 3989 5475 4015 5501
rect 4041 5475 5563 5501
rect 5589 5475 5615 5501
rect 5641 5475 5667 5501
rect 5693 5475 7215 5501
rect 7241 5475 7267 5501
rect 7293 5475 7319 5501
rect 7345 5475 7360 5501
rect 672 5458 7360 5475
rect 4489 5335 4495 5361
rect 4521 5335 4527 5361
rect 5273 5335 5279 5361
rect 5305 5335 5311 5361
rect 4327 5249 4353 5255
rect 4769 5223 4775 5249
rect 4801 5223 4807 5249
rect 4327 5217 4353 5223
rect 672 5109 7280 5126
rect 672 5083 1433 5109
rect 1459 5083 1485 5109
rect 1511 5083 1537 5109
rect 1563 5083 3085 5109
rect 3111 5083 3137 5109
rect 3163 5083 3189 5109
rect 3215 5083 4737 5109
rect 4763 5083 4789 5109
rect 4815 5083 4841 5109
rect 4867 5083 6389 5109
rect 6415 5083 6441 5109
rect 6467 5083 6493 5109
rect 6519 5083 7280 5109
rect 672 5066 7280 5083
rect 4825 4943 4831 4969
rect 4857 4943 4863 4969
rect 3481 4887 3487 4913
rect 3513 4887 3519 4913
rect 4153 4887 4159 4913
rect 4185 4887 4191 4913
rect 3487 4801 3513 4807
rect 3487 4769 3513 4775
rect 672 4717 7360 4734
rect 672 4691 2259 4717
rect 2285 4691 2311 4717
rect 2337 4691 2363 4717
rect 2389 4691 3911 4717
rect 3937 4691 3963 4717
rect 3989 4691 4015 4717
rect 4041 4691 5563 4717
rect 5589 4691 5615 4717
rect 5641 4691 5667 4717
rect 5693 4691 7215 4717
rect 7241 4691 7267 4717
rect 7293 4691 7319 4717
rect 7345 4691 7360 4717
rect 672 4674 7360 4691
rect 4271 4633 4297 4639
rect 4271 4601 4297 4607
rect 1023 4577 1049 4583
rect 1023 4545 1049 4551
rect 3879 4577 3905 4583
rect 5889 4551 5895 4577
rect 5921 4551 5927 4577
rect 7009 4551 7015 4577
rect 7041 4551 7047 4577
rect 3879 4545 3905 4551
rect 855 4521 881 4527
rect 855 4489 881 4495
rect 2423 4521 2449 4527
rect 2753 4495 2759 4521
rect 2785 4495 2791 4521
rect 6449 4495 6455 4521
rect 6481 4495 6487 4521
rect 2423 4489 2449 4495
rect 1247 4465 1273 4471
rect 5385 4439 5391 4465
rect 5417 4439 5423 4465
rect 1247 4433 1273 4439
rect 672 4325 7280 4342
rect 672 4299 1433 4325
rect 1459 4299 1485 4325
rect 1511 4299 1537 4325
rect 1563 4299 3085 4325
rect 3111 4299 3137 4325
rect 3163 4299 3189 4325
rect 3215 4299 4737 4325
rect 4763 4299 4789 4325
rect 4815 4299 4841 4325
rect 4867 4299 6389 4325
rect 6415 4299 6441 4325
rect 6467 4299 6493 4325
rect 6519 4299 7280 4325
rect 672 4282 7280 4299
rect 6511 4185 6537 4191
rect 2865 4159 2871 4185
rect 2897 4159 2903 4185
rect 6511 4153 6537 4159
rect 2591 4129 2617 4135
rect 6791 4129 6817 4135
rect 2977 4103 2983 4129
rect 3009 4103 3015 4129
rect 3201 4103 3207 4129
rect 3233 4103 3239 4129
rect 6113 4103 6119 4129
rect 6145 4103 6151 4129
rect 2591 4097 2617 4103
rect 6791 4097 6817 4103
rect 7071 4129 7097 4135
rect 7071 4097 7097 4103
rect 4209 4047 4215 4073
rect 4241 4047 4247 4073
rect 6001 4047 6007 4073
rect 6033 4047 6039 4073
rect 672 3933 7360 3950
rect 672 3907 2259 3933
rect 2285 3907 2311 3933
rect 2337 3907 2363 3933
rect 2389 3907 3911 3933
rect 3937 3907 3963 3933
rect 3989 3907 4015 3933
rect 4041 3907 5563 3933
rect 5589 3907 5615 3933
rect 5641 3907 5667 3933
rect 5693 3907 7215 3933
rect 7241 3907 7267 3933
rect 7293 3907 7319 3933
rect 7345 3907 7360 3933
rect 672 3890 7360 3907
rect 2417 3767 2423 3793
rect 2449 3767 2455 3793
rect 5945 3767 5951 3793
rect 5977 3767 5983 3793
rect 4209 3711 4215 3737
rect 4241 3711 4247 3737
rect 6449 3711 6455 3737
rect 6481 3711 6487 3737
rect 5273 3655 5279 3681
rect 5305 3655 5311 3681
rect 7009 3655 7015 3681
rect 7041 3655 7047 3681
rect 672 3541 7280 3558
rect 672 3515 1433 3541
rect 1459 3515 1485 3541
rect 1511 3515 1537 3541
rect 1563 3515 3085 3541
rect 3111 3515 3137 3541
rect 3163 3515 3189 3541
rect 3215 3515 4737 3541
rect 4763 3515 4789 3541
rect 4815 3515 4841 3541
rect 4867 3515 6389 3541
rect 6415 3515 6441 3541
rect 6467 3515 6493 3541
rect 6519 3515 7280 3541
rect 672 3498 7280 3515
rect 1073 3375 1079 3401
rect 1105 3375 1111 3401
rect 1471 3345 1497 3351
rect 5895 3345 5921 3351
rect 2473 3319 2479 3345
rect 2505 3319 2511 3345
rect 4097 3319 4103 3345
rect 4129 3319 4135 3345
rect 4377 3319 4383 3345
rect 4409 3319 4415 3345
rect 1471 3313 1497 3319
rect 5895 3313 5921 3319
rect 2367 3289 2393 3295
rect 2367 3257 2393 3263
rect 7071 3289 7097 3295
rect 7071 3257 7097 3263
rect 2983 3233 3009 3239
rect 2983 3201 3009 3207
rect 3375 3233 3401 3239
rect 3375 3201 3401 3207
rect 3543 3233 3569 3239
rect 3543 3201 3569 3207
rect 3935 3233 3961 3239
rect 6903 3233 6929 3239
rect 5609 3207 5615 3233
rect 5641 3207 5647 3233
rect 3935 3201 3961 3207
rect 6903 3201 6929 3207
rect 672 3149 7360 3166
rect 672 3123 2259 3149
rect 2285 3123 2311 3149
rect 2337 3123 2363 3149
rect 2389 3123 3911 3149
rect 3937 3123 3963 3149
rect 3989 3123 4015 3149
rect 4041 3123 5563 3149
rect 5589 3123 5615 3149
rect 5641 3123 5667 3149
rect 5693 3123 7215 3149
rect 7241 3123 7267 3149
rect 7293 3123 7319 3149
rect 7345 3123 7360 3149
rect 672 3106 7360 3123
rect 1023 3065 1049 3071
rect 1023 3033 1049 3039
rect 1247 3065 1273 3071
rect 5167 3065 5193 3071
rect 3481 3039 3487 3065
rect 3513 3039 3519 3065
rect 1247 3033 1273 3039
rect 5167 3033 5193 3039
rect 7127 3065 7153 3071
rect 7127 3033 7153 3039
rect 855 3009 881 3015
rect 855 2977 881 2983
rect 4159 3009 4185 3015
rect 4159 2977 4185 2983
rect 2143 2953 2169 2959
rect 2305 2927 2311 2953
rect 2337 2927 2343 2953
rect 4041 2927 4047 2953
rect 4073 2927 4079 2953
rect 4825 2927 4831 2953
rect 4857 2927 4863 2953
rect 2143 2921 2169 2927
rect 3879 2841 3905 2847
rect 3879 2809 3905 2815
rect 672 2757 7280 2774
rect 672 2731 1433 2757
rect 1459 2731 1485 2757
rect 1511 2731 1537 2757
rect 1563 2731 3085 2757
rect 3111 2731 3137 2757
rect 3163 2731 3189 2757
rect 3215 2731 4737 2757
rect 4763 2731 4789 2757
rect 4815 2731 4841 2757
rect 4867 2731 6389 2757
rect 6415 2731 6441 2757
rect 6467 2731 6493 2757
rect 6519 2731 7280 2757
rect 672 2714 7280 2731
rect 3033 2591 3039 2617
rect 3065 2591 3071 2617
rect 2815 2561 2841 2567
rect 2815 2529 2841 2535
rect 3375 2561 3401 2567
rect 4825 2535 4831 2561
rect 4857 2535 4863 2561
rect 3375 2529 3401 2535
rect 3543 2449 3569 2455
rect 3543 2417 3569 2423
rect 4943 2449 4969 2455
rect 4943 2417 4969 2423
rect 672 2365 7360 2382
rect 672 2339 2259 2365
rect 2285 2339 2311 2365
rect 2337 2339 2363 2365
rect 2389 2339 3911 2365
rect 3937 2339 3963 2365
rect 3989 2339 4015 2365
rect 4041 2339 5563 2365
rect 5589 2339 5615 2365
rect 5641 2339 5667 2365
rect 5693 2339 7215 2365
rect 7241 2339 7267 2365
rect 7293 2339 7319 2365
rect 7345 2339 7360 2365
rect 672 2322 7360 2339
rect 3991 2281 4017 2287
rect 3991 2249 4017 2255
rect 3823 2169 3849 2175
rect 3823 2137 3849 2143
rect 3711 2113 3737 2119
rect 3711 2081 3737 2087
rect 672 1973 7280 1990
rect 672 1947 1433 1973
rect 1459 1947 1485 1973
rect 1511 1947 1537 1973
rect 1563 1947 3085 1973
rect 3111 1947 3137 1973
rect 3163 1947 3189 1973
rect 3215 1947 4737 1973
rect 4763 1947 4789 1973
rect 4815 1947 4841 1973
rect 4867 1947 6389 1973
rect 6415 1947 6441 1973
rect 6467 1947 6493 1973
rect 6519 1947 7280 1973
rect 672 1930 7280 1947
rect 3761 1807 3767 1833
rect 3793 1807 3799 1833
rect 4881 1807 4887 1833
rect 4913 1807 4919 1833
rect 4663 1777 4689 1783
rect 3537 1751 3543 1777
rect 3569 1751 3575 1777
rect 4663 1745 4689 1751
rect 3039 1721 3065 1727
rect 3039 1689 3065 1695
rect 3151 1721 3177 1727
rect 3151 1689 3177 1695
rect 3319 1721 3345 1727
rect 3319 1689 3345 1695
rect 672 1581 7360 1598
rect 672 1555 2259 1581
rect 2285 1555 2311 1581
rect 2337 1555 2363 1581
rect 2389 1555 3911 1581
rect 3937 1555 3963 1581
rect 3989 1555 4015 1581
rect 4041 1555 5563 1581
rect 5589 1555 5615 1581
rect 5641 1555 5667 1581
rect 5693 1555 7215 1581
rect 7241 1555 7267 1581
rect 7293 1555 7319 1581
rect 7345 1555 7360 1581
rect 672 1538 7360 1555
<< via1 >>
rect 2259 6259 2285 6285
rect 2311 6259 2337 6285
rect 2363 6259 2389 6285
rect 3911 6259 3937 6285
rect 3963 6259 3989 6285
rect 4015 6259 4041 6285
rect 5563 6259 5589 6285
rect 5615 6259 5641 6285
rect 5667 6259 5693 6285
rect 7215 6259 7241 6285
rect 7267 6259 7293 6285
rect 7319 6259 7345 6285
rect 1433 5867 1459 5893
rect 1485 5867 1511 5893
rect 1537 5867 1563 5893
rect 3085 5867 3111 5893
rect 3137 5867 3163 5893
rect 3189 5867 3215 5893
rect 4737 5867 4763 5893
rect 4789 5867 4815 5893
rect 4841 5867 4867 5893
rect 6389 5867 6415 5893
rect 6441 5867 6467 5893
rect 6493 5867 6519 5893
rect 3543 5671 3569 5697
rect 3767 5671 3793 5697
rect 4887 5559 4913 5585
rect 5279 5559 5305 5585
rect 2259 5475 2285 5501
rect 2311 5475 2337 5501
rect 2363 5475 2389 5501
rect 3911 5475 3937 5501
rect 3963 5475 3989 5501
rect 4015 5475 4041 5501
rect 5563 5475 5589 5501
rect 5615 5475 5641 5501
rect 5667 5475 5693 5501
rect 7215 5475 7241 5501
rect 7267 5475 7293 5501
rect 7319 5475 7345 5501
rect 4495 5335 4521 5361
rect 5279 5335 5305 5361
rect 4327 5223 4353 5249
rect 4775 5223 4801 5249
rect 1433 5083 1459 5109
rect 1485 5083 1511 5109
rect 1537 5083 1563 5109
rect 3085 5083 3111 5109
rect 3137 5083 3163 5109
rect 3189 5083 3215 5109
rect 4737 5083 4763 5109
rect 4789 5083 4815 5109
rect 4841 5083 4867 5109
rect 6389 5083 6415 5109
rect 6441 5083 6467 5109
rect 6493 5083 6519 5109
rect 4831 4943 4857 4969
rect 3487 4887 3513 4913
rect 4159 4887 4185 4913
rect 3487 4775 3513 4801
rect 2259 4691 2285 4717
rect 2311 4691 2337 4717
rect 2363 4691 2389 4717
rect 3911 4691 3937 4717
rect 3963 4691 3989 4717
rect 4015 4691 4041 4717
rect 5563 4691 5589 4717
rect 5615 4691 5641 4717
rect 5667 4691 5693 4717
rect 7215 4691 7241 4717
rect 7267 4691 7293 4717
rect 7319 4691 7345 4717
rect 4271 4607 4297 4633
rect 1023 4551 1049 4577
rect 3879 4551 3905 4577
rect 5895 4551 5921 4577
rect 7015 4551 7041 4577
rect 855 4495 881 4521
rect 2423 4495 2449 4521
rect 2759 4495 2785 4521
rect 6455 4495 6481 4521
rect 1247 4439 1273 4465
rect 5391 4439 5417 4465
rect 1433 4299 1459 4325
rect 1485 4299 1511 4325
rect 1537 4299 1563 4325
rect 3085 4299 3111 4325
rect 3137 4299 3163 4325
rect 3189 4299 3215 4325
rect 4737 4299 4763 4325
rect 4789 4299 4815 4325
rect 4841 4299 4867 4325
rect 6389 4299 6415 4325
rect 6441 4299 6467 4325
rect 6493 4299 6519 4325
rect 2871 4159 2897 4185
rect 6511 4159 6537 4185
rect 2591 4103 2617 4129
rect 2983 4103 3009 4129
rect 3207 4103 3233 4129
rect 6119 4103 6145 4129
rect 6791 4103 6817 4129
rect 7071 4103 7097 4129
rect 4215 4047 4241 4073
rect 6007 4047 6033 4073
rect 2259 3907 2285 3933
rect 2311 3907 2337 3933
rect 2363 3907 2389 3933
rect 3911 3907 3937 3933
rect 3963 3907 3989 3933
rect 4015 3907 4041 3933
rect 5563 3907 5589 3933
rect 5615 3907 5641 3933
rect 5667 3907 5693 3933
rect 7215 3907 7241 3933
rect 7267 3907 7293 3933
rect 7319 3907 7345 3933
rect 2423 3767 2449 3793
rect 5951 3767 5977 3793
rect 4215 3711 4241 3737
rect 6455 3711 6481 3737
rect 5279 3655 5305 3681
rect 7015 3655 7041 3681
rect 1433 3515 1459 3541
rect 1485 3515 1511 3541
rect 1537 3515 1563 3541
rect 3085 3515 3111 3541
rect 3137 3515 3163 3541
rect 3189 3515 3215 3541
rect 4737 3515 4763 3541
rect 4789 3515 4815 3541
rect 4841 3515 4867 3541
rect 6389 3515 6415 3541
rect 6441 3515 6467 3541
rect 6493 3515 6519 3541
rect 1079 3375 1105 3401
rect 1471 3319 1497 3345
rect 2479 3319 2505 3345
rect 4103 3319 4129 3345
rect 4383 3319 4409 3345
rect 5895 3319 5921 3345
rect 2367 3263 2393 3289
rect 7071 3263 7097 3289
rect 2983 3207 3009 3233
rect 3375 3207 3401 3233
rect 3543 3207 3569 3233
rect 3935 3207 3961 3233
rect 5615 3207 5641 3233
rect 6903 3207 6929 3233
rect 2259 3123 2285 3149
rect 2311 3123 2337 3149
rect 2363 3123 2389 3149
rect 3911 3123 3937 3149
rect 3963 3123 3989 3149
rect 4015 3123 4041 3149
rect 5563 3123 5589 3149
rect 5615 3123 5641 3149
rect 5667 3123 5693 3149
rect 7215 3123 7241 3149
rect 7267 3123 7293 3149
rect 7319 3123 7345 3149
rect 1023 3039 1049 3065
rect 1247 3039 1273 3065
rect 3487 3039 3513 3065
rect 5167 3039 5193 3065
rect 7127 3039 7153 3065
rect 855 2983 881 3009
rect 4159 2983 4185 3009
rect 2143 2927 2169 2953
rect 2311 2927 2337 2953
rect 4047 2927 4073 2953
rect 4831 2927 4857 2953
rect 3879 2815 3905 2841
rect 1433 2731 1459 2757
rect 1485 2731 1511 2757
rect 1537 2731 1563 2757
rect 3085 2731 3111 2757
rect 3137 2731 3163 2757
rect 3189 2731 3215 2757
rect 4737 2731 4763 2757
rect 4789 2731 4815 2757
rect 4841 2731 4867 2757
rect 6389 2731 6415 2757
rect 6441 2731 6467 2757
rect 6493 2731 6519 2757
rect 3039 2591 3065 2617
rect 2815 2535 2841 2561
rect 3375 2535 3401 2561
rect 4831 2535 4857 2561
rect 3543 2423 3569 2449
rect 4943 2423 4969 2449
rect 2259 2339 2285 2365
rect 2311 2339 2337 2365
rect 2363 2339 2389 2365
rect 3911 2339 3937 2365
rect 3963 2339 3989 2365
rect 4015 2339 4041 2365
rect 5563 2339 5589 2365
rect 5615 2339 5641 2365
rect 5667 2339 5693 2365
rect 7215 2339 7241 2365
rect 7267 2339 7293 2365
rect 7319 2339 7345 2365
rect 3991 2255 4017 2281
rect 3823 2143 3849 2169
rect 3711 2087 3737 2113
rect 1433 1947 1459 1973
rect 1485 1947 1511 1973
rect 1537 1947 1563 1973
rect 3085 1947 3111 1973
rect 3137 1947 3163 1973
rect 3189 1947 3215 1973
rect 4737 1947 4763 1973
rect 4789 1947 4815 1973
rect 4841 1947 4867 1973
rect 6389 1947 6415 1973
rect 6441 1947 6467 1973
rect 6493 1947 6519 1973
rect 3767 1807 3793 1833
rect 4887 1807 4913 1833
rect 3543 1751 3569 1777
rect 4663 1751 4689 1777
rect 3039 1695 3065 1721
rect 3151 1695 3177 1721
rect 3319 1695 3345 1721
rect 2259 1555 2285 1581
rect 2311 1555 2337 1581
rect 2363 1555 2389 1581
rect 3911 1555 3937 1581
rect 3963 1555 3989 1581
rect 4015 1555 4041 1581
rect 5563 1555 5589 1581
rect 5615 1555 5641 1581
rect 5667 1555 5693 1581
rect 7215 1555 7241 1581
rect 7267 1555 7293 1581
rect 7319 1555 7345 1581
<< metal2 >>
rect 2258 6286 2390 6291
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2258 6253 2390 6258
rect 3910 6286 4042 6291
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 3910 6253 4042 6258
rect 5562 6286 5694 6291
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5562 6253 5694 6258
rect 7214 6286 7346 6291
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7214 6253 7346 6258
rect 1432 5894 1564 5899
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1432 5861 1564 5866
rect 3084 5894 3216 5899
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3084 5861 3216 5866
rect 4736 5894 4868 5899
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4736 5861 4868 5866
rect 6388 5894 6520 5899
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6388 5861 6520 5866
rect 3542 5697 3570 5703
rect 3542 5671 3543 5697
rect 3569 5671 3570 5697
rect 2258 5502 2390 5507
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2258 5469 2390 5474
rect 1432 5110 1564 5115
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1432 5077 1564 5082
rect 3084 5110 3216 5115
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3084 5077 3216 5082
rect 3542 4970 3570 5671
rect 3766 5697 3794 5703
rect 3766 5671 3767 5697
rect 3793 5671 3794 5697
rect 3766 5250 3794 5671
rect 4886 5586 4914 5591
rect 4494 5585 4914 5586
rect 4494 5559 4887 5585
rect 4913 5559 4914 5585
rect 4494 5558 4914 5559
rect 3910 5502 4042 5507
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 3910 5469 4042 5474
rect 3766 5217 3794 5222
rect 4270 5362 4298 5367
rect 3542 4937 3570 4942
rect 4102 4970 4130 4975
rect 2982 4914 3010 4919
rect 2258 4718 2390 4723
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2258 4685 2390 4690
rect 1022 4577 1050 4583
rect 1022 4551 1023 4577
rect 1049 4551 1050 4577
rect 854 4521 882 4527
rect 854 4495 855 4521
rect 881 4495 882 4521
rect 854 4410 882 4495
rect 854 4377 882 4382
rect 1022 3626 1050 4551
rect 2478 4578 2506 4583
rect 2422 4521 2450 4527
rect 2422 4495 2423 4521
rect 2449 4495 2450 4521
rect 1246 4465 1274 4471
rect 1246 4439 1247 4465
rect 1273 4439 1274 4465
rect 1246 4410 1274 4439
rect 1246 4377 1274 4382
rect 1432 4326 1564 4331
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1432 4293 1564 4298
rect 2258 3934 2390 3939
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2258 3901 2390 3906
rect 2422 3794 2450 4495
rect 2478 4214 2506 4550
rect 2870 4578 2898 4583
rect 2758 4521 2786 4527
rect 2758 4495 2759 4521
rect 2785 4495 2786 4521
rect 2758 4242 2786 4495
rect 2478 4186 2618 4214
rect 2758 4209 2786 4214
rect 2590 4130 2618 4186
rect 2870 4185 2898 4550
rect 2870 4159 2871 4185
rect 2897 4159 2898 4185
rect 2870 4153 2898 4159
rect 2590 4083 2618 4102
rect 2982 4129 3010 4886
rect 3486 4914 3514 4933
rect 3486 4881 3514 4886
rect 3486 4801 3514 4807
rect 3486 4775 3487 4801
rect 3513 4775 3514 4801
rect 3084 4326 3216 4331
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3084 4293 3216 4298
rect 2982 4103 2983 4129
rect 3009 4103 3010 4129
rect 2982 4097 3010 4103
rect 3206 4130 3234 4135
rect 3206 4083 3234 4102
rect 2142 3793 2450 3794
rect 2142 3767 2423 3793
rect 2449 3767 2450 3793
rect 2142 3766 2450 3767
rect 1022 3593 1050 3598
rect 2030 3738 2058 3743
rect 1432 3542 1564 3547
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1432 3509 1564 3514
rect 1078 3402 1106 3407
rect 1078 3355 1106 3374
rect 1470 3402 1498 3407
rect 1470 3345 1498 3374
rect 1470 3319 1471 3345
rect 1497 3319 1498 3345
rect 1470 3313 1498 3319
rect 1022 3290 1050 3295
rect 854 3066 882 3071
rect 854 3009 882 3038
rect 1022 3065 1050 3262
rect 1022 3039 1023 3065
rect 1049 3039 1050 3065
rect 1022 3033 1050 3039
rect 1246 3066 1274 3071
rect 1246 3019 1274 3038
rect 854 2983 855 3009
rect 881 2983 882 3009
rect 854 2977 882 2983
rect 1432 2758 1564 2763
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1432 2725 1564 2730
rect 2030 2674 2058 3710
rect 2142 2953 2170 3766
rect 2422 3761 2450 3766
rect 2142 2927 2143 2953
rect 2169 2927 2170 2953
rect 2142 2921 2170 2927
rect 2198 3626 2226 3631
rect 2198 2954 2226 3598
rect 3084 3542 3216 3547
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3084 3509 3216 3514
rect 2366 3402 2394 3407
rect 2366 3289 2394 3374
rect 2366 3263 2367 3289
rect 2393 3263 2394 3289
rect 2366 3257 2394 3263
rect 2478 3345 2506 3351
rect 2478 3319 2479 3345
rect 2505 3319 2506 3345
rect 2478 3290 2506 3319
rect 2478 3257 2506 3262
rect 2814 3290 2842 3295
rect 2258 3150 2390 3155
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2258 3117 2390 3122
rect 2310 2954 2338 2959
rect 2198 2953 2338 2954
rect 2198 2927 2311 2953
rect 2337 2927 2338 2953
rect 2198 2926 2338 2927
rect 2310 2921 2338 2926
rect 2030 2641 2058 2646
rect 2814 2561 2842 3262
rect 2982 3234 3010 3239
rect 2814 2535 2815 2561
rect 2841 2535 2842 2561
rect 2814 2529 2842 2535
rect 2870 3233 3010 3234
rect 2870 3207 2983 3233
rect 3009 3207 3010 3233
rect 2870 3206 3010 3207
rect 2258 2366 2390 2371
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2258 2333 2390 2338
rect 1432 1974 1564 1979
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1432 1941 1564 1946
rect 2258 1582 2390 1587
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2258 1549 2390 1554
rect 2870 490 2898 3206
rect 2982 3201 3010 3206
rect 3374 3233 3402 3239
rect 3374 3207 3375 3233
rect 3401 3207 3402 3233
rect 3084 2758 3216 2763
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3084 2725 3216 2730
rect 3038 2674 3066 2679
rect 3038 2617 3066 2646
rect 3038 2591 3039 2617
rect 3065 2591 3066 2617
rect 3038 2585 3066 2591
rect 3374 2562 3402 3207
rect 3486 3065 3514 4775
rect 3910 4718 4042 4723
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 3910 4685 4042 4690
rect 3878 4578 3906 4583
rect 3878 4531 3906 4550
rect 3910 3934 4042 3939
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 3910 3901 4042 3906
rect 4102 3345 4130 4942
rect 4158 4913 4186 4919
rect 4158 4887 4159 4913
rect 4185 4887 4186 4913
rect 4158 4074 4186 4887
rect 4270 4633 4298 5334
rect 4494 5361 4522 5558
rect 4886 5553 4914 5558
rect 5278 5586 5306 5591
rect 5278 5585 5362 5586
rect 5278 5559 5279 5585
rect 5305 5559 5362 5585
rect 5278 5558 5362 5559
rect 5278 5553 5306 5558
rect 4494 5335 4495 5361
rect 4521 5335 4522 5361
rect 4494 5329 4522 5335
rect 5278 5362 5306 5367
rect 5278 5315 5306 5334
rect 4270 4607 4271 4633
rect 4297 4607 4298 4633
rect 4270 4601 4298 4607
rect 4326 5249 4354 5255
rect 4326 5223 4327 5249
rect 4353 5223 4354 5249
rect 4326 4914 4354 5223
rect 4774 5250 4802 5255
rect 4774 5203 4802 5222
rect 4736 5110 4868 5115
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4736 5077 4868 5082
rect 4830 4970 4858 4975
rect 4830 4923 4858 4942
rect 4326 4214 4354 4886
rect 5334 4578 5362 5558
rect 5562 5502 5694 5507
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5562 5469 5694 5474
rect 7214 5502 7346 5507
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7214 5469 7346 5474
rect 6388 5110 6520 5115
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6388 5077 6520 5082
rect 5562 4718 5694 4723
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5562 4685 5694 4690
rect 7214 4718 7346 4723
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7214 4685 7346 4690
rect 7014 4634 7042 4639
rect 5334 4545 5362 4550
rect 5894 4578 5922 4583
rect 5894 4531 5922 4550
rect 7014 4577 7042 4606
rect 7014 4551 7015 4577
rect 7041 4551 7042 4577
rect 7014 4545 7042 4551
rect 6454 4522 6482 4527
rect 5950 4521 6482 4522
rect 5950 4495 6455 4521
rect 6481 4495 6482 4521
rect 5950 4494 6482 4495
rect 5390 4465 5418 4471
rect 5390 4439 5391 4465
rect 5417 4439 5418 4465
rect 4736 4326 4868 4331
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4736 4293 4868 4298
rect 5278 4242 5306 4247
rect 4326 4186 4410 4214
rect 4382 4130 4410 4186
rect 4382 4097 4410 4102
rect 4214 4074 4242 4079
rect 4158 4073 4242 4074
rect 4158 4047 4215 4073
rect 4241 4047 4242 4073
rect 4158 4046 4242 4047
rect 4214 3737 4242 4046
rect 4214 3711 4215 3737
rect 4241 3711 4242 3737
rect 4214 3705 4242 3711
rect 4382 3794 4410 3799
rect 4102 3319 4103 3345
rect 4129 3319 4130 3345
rect 4102 3313 4130 3319
rect 4382 3345 4410 3766
rect 4998 3738 5026 3743
rect 4736 3542 4868 3547
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4736 3509 4868 3514
rect 4382 3319 4383 3345
rect 4409 3319 4410 3345
rect 4382 3313 4410 3319
rect 3542 3234 3570 3239
rect 3934 3234 3962 3239
rect 4830 3234 4858 3239
rect 3542 3233 3626 3234
rect 3542 3207 3543 3233
rect 3569 3207 3626 3233
rect 3542 3206 3626 3207
rect 3542 3201 3570 3206
rect 3486 3039 3487 3065
rect 3513 3039 3514 3065
rect 3486 3033 3514 3039
rect 3318 2561 3402 2562
rect 3318 2535 3375 2561
rect 3401 2535 3402 2561
rect 3318 2534 3402 2535
rect 3084 1974 3216 1979
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3084 1941 3216 1946
rect 2702 462 2898 490
rect 3038 1722 3066 1727
rect 3150 1722 3178 1727
rect 3038 1721 3178 1722
rect 3038 1695 3039 1721
rect 3065 1695 3151 1721
rect 3177 1695 3178 1721
rect 3038 1694 3178 1695
rect 2702 400 2730 462
rect 3038 400 3066 1694
rect 3150 1689 3178 1694
rect 3318 1721 3346 2534
rect 3374 2529 3402 2534
rect 3542 2449 3570 2455
rect 3542 2423 3543 2449
rect 3569 2423 3570 2449
rect 3486 1834 3514 1839
rect 3318 1695 3319 1721
rect 3345 1695 3346 1721
rect 3318 1689 3346 1695
rect 3374 1806 3486 1834
rect 3374 400 3402 1806
rect 3486 1801 3514 1806
rect 3542 1777 3570 2423
rect 3598 1946 3626 3206
rect 3934 3233 4130 3234
rect 3934 3207 3935 3233
rect 3961 3207 4130 3233
rect 3934 3206 4130 3207
rect 3934 3201 3962 3206
rect 3910 3150 4042 3155
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 3910 3117 4042 3122
rect 4046 2954 4074 2959
rect 4102 2954 4130 3206
rect 4046 2953 4130 2954
rect 4046 2927 4047 2953
rect 4073 2927 4130 2953
rect 4046 2926 4130 2927
rect 4046 2921 4074 2926
rect 3878 2842 3906 2847
rect 3878 2795 3906 2814
rect 3910 2366 4042 2371
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 3910 2333 4042 2338
rect 3990 2282 4018 2287
rect 4102 2282 4130 2926
rect 3990 2281 4130 2282
rect 3990 2255 3991 2281
rect 4017 2255 4130 2281
rect 3990 2254 4130 2255
rect 4158 3009 4186 3015
rect 4158 2983 4159 3009
rect 4185 2983 4186 3009
rect 3990 2249 4018 2254
rect 3822 2169 3850 2175
rect 3822 2143 3823 2169
rect 3849 2143 3850 2169
rect 3710 2114 3738 2119
rect 3822 2114 3850 2143
rect 3710 2113 3850 2114
rect 3710 2087 3711 2113
rect 3737 2087 3850 2113
rect 3710 2086 3850 2087
rect 3710 2081 3738 2086
rect 3598 1913 3626 1918
rect 3766 1834 3794 1839
rect 3766 1787 3794 1806
rect 3542 1751 3543 1777
rect 3569 1751 3570 1777
rect 3542 1745 3570 1751
rect 3822 1442 3850 2086
rect 4102 1834 4130 1839
rect 3910 1582 4042 1587
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 3910 1549 4042 1554
rect 3710 1414 3850 1442
rect 3710 400 3738 1414
rect 4102 602 4130 1806
rect 4158 1778 4186 2983
rect 4830 2954 4858 3206
rect 4830 2953 4970 2954
rect 4830 2927 4831 2953
rect 4857 2927 4970 2953
rect 4830 2926 4970 2927
rect 4830 2921 4858 2926
rect 4736 2758 4868 2763
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4736 2725 4868 2730
rect 4830 2562 4858 2567
rect 4942 2562 4970 2926
rect 4830 2561 4970 2562
rect 4830 2535 4831 2561
rect 4857 2535 4970 2561
rect 4830 2534 4970 2535
rect 4830 2529 4858 2534
rect 4942 2450 4970 2455
rect 4998 2450 5026 3710
rect 5166 3682 5194 3687
rect 5166 3065 5194 3654
rect 5278 3681 5306 4214
rect 5390 3794 5418 4439
rect 5950 4214 5978 4494
rect 6454 4489 6482 4494
rect 6388 4326 6520 4331
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6388 4293 6520 4298
rect 5894 4186 5978 4214
rect 6510 4186 6538 4191
rect 5562 3934 5694 3939
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5562 3901 5694 3906
rect 5390 3761 5418 3766
rect 5278 3655 5279 3681
rect 5305 3655 5306 3681
rect 5278 3649 5306 3655
rect 5614 3626 5642 3631
rect 5614 3233 5642 3598
rect 5894 3345 5922 4186
rect 6510 4139 6538 4158
rect 7070 4186 7098 4191
rect 6118 4130 6146 4135
rect 6118 4083 6146 4102
rect 6790 4130 6818 4135
rect 6790 4083 6818 4102
rect 7070 4129 7098 4158
rect 7070 4103 7071 4129
rect 7097 4103 7098 4129
rect 7070 4097 7098 4103
rect 6006 4073 6034 4079
rect 6006 4047 6007 4073
rect 6033 4047 6034 4073
rect 5894 3319 5895 3345
rect 5921 3319 5922 3345
rect 5894 3313 5922 3319
rect 5950 3793 5978 3799
rect 5950 3767 5951 3793
rect 5977 3767 5978 3793
rect 5614 3207 5615 3233
rect 5641 3207 5642 3233
rect 5614 3201 5642 3207
rect 5562 3150 5694 3155
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5562 3117 5694 3122
rect 5166 3039 5167 3065
rect 5193 3039 5194 3065
rect 5166 3033 5194 3039
rect 5950 2842 5978 3767
rect 6006 3626 6034 4047
rect 7214 3934 7346 3939
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7214 3901 7346 3906
rect 6454 3738 6482 3743
rect 6454 3691 6482 3710
rect 6006 3593 6034 3598
rect 7014 3681 7042 3687
rect 7014 3655 7015 3681
rect 7041 3655 7042 3681
rect 6388 3542 6520 3547
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6388 3509 6520 3514
rect 7014 3402 7042 3655
rect 7014 3369 7042 3374
rect 7070 3289 7098 3295
rect 7070 3263 7071 3289
rect 7097 3263 7098 3289
rect 6902 3234 6930 3239
rect 6902 3187 6930 3206
rect 7070 3066 7098 3263
rect 7214 3150 7346 3155
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7214 3117 7346 3122
rect 7126 3066 7154 3071
rect 7070 3038 7126 3066
rect 7126 3019 7154 3038
rect 5950 2809 5978 2814
rect 6388 2758 6520 2763
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6388 2725 6520 2730
rect 4942 2449 5026 2450
rect 4942 2423 4943 2449
rect 4969 2423 5026 2449
rect 4942 2422 5026 2423
rect 4942 2417 4970 2422
rect 5562 2366 5694 2371
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5562 2333 5694 2338
rect 7214 2366 7346 2371
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7214 2333 7346 2338
rect 4736 1974 4868 1979
rect 4158 1745 4186 1750
rect 4382 1946 4410 1951
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4736 1941 4868 1946
rect 6388 1974 6520 1979
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6388 1941 6520 1946
rect 4046 574 4130 602
rect 4046 400 4074 574
rect 4382 400 4410 1918
rect 4886 1834 4914 1839
rect 4886 1787 4914 1806
rect 4662 1778 4690 1783
rect 4662 1731 4690 1750
rect 5562 1582 5694 1587
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5562 1549 5694 1554
rect 7214 1582 7346 1587
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7214 1549 7346 1554
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
<< via2 >>
rect 2258 6285 2286 6286
rect 2258 6259 2259 6285
rect 2259 6259 2285 6285
rect 2285 6259 2286 6285
rect 2258 6258 2286 6259
rect 2310 6285 2338 6286
rect 2310 6259 2311 6285
rect 2311 6259 2337 6285
rect 2337 6259 2338 6285
rect 2310 6258 2338 6259
rect 2362 6285 2390 6286
rect 2362 6259 2363 6285
rect 2363 6259 2389 6285
rect 2389 6259 2390 6285
rect 2362 6258 2390 6259
rect 3910 6285 3938 6286
rect 3910 6259 3911 6285
rect 3911 6259 3937 6285
rect 3937 6259 3938 6285
rect 3910 6258 3938 6259
rect 3962 6285 3990 6286
rect 3962 6259 3963 6285
rect 3963 6259 3989 6285
rect 3989 6259 3990 6285
rect 3962 6258 3990 6259
rect 4014 6285 4042 6286
rect 4014 6259 4015 6285
rect 4015 6259 4041 6285
rect 4041 6259 4042 6285
rect 4014 6258 4042 6259
rect 5562 6285 5590 6286
rect 5562 6259 5563 6285
rect 5563 6259 5589 6285
rect 5589 6259 5590 6285
rect 5562 6258 5590 6259
rect 5614 6285 5642 6286
rect 5614 6259 5615 6285
rect 5615 6259 5641 6285
rect 5641 6259 5642 6285
rect 5614 6258 5642 6259
rect 5666 6285 5694 6286
rect 5666 6259 5667 6285
rect 5667 6259 5693 6285
rect 5693 6259 5694 6285
rect 5666 6258 5694 6259
rect 7214 6285 7242 6286
rect 7214 6259 7215 6285
rect 7215 6259 7241 6285
rect 7241 6259 7242 6285
rect 7214 6258 7242 6259
rect 7266 6285 7294 6286
rect 7266 6259 7267 6285
rect 7267 6259 7293 6285
rect 7293 6259 7294 6285
rect 7266 6258 7294 6259
rect 7318 6285 7346 6286
rect 7318 6259 7319 6285
rect 7319 6259 7345 6285
rect 7345 6259 7346 6285
rect 7318 6258 7346 6259
rect 1432 5893 1460 5894
rect 1432 5867 1433 5893
rect 1433 5867 1459 5893
rect 1459 5867 1460 5893
rect 1432 5866 1460 5867
rect 1484 5893 1512 5894
rect 1484 5867 1485 5893
rect 1485 5867 1511 5893
rect 1511 5867 1512 5893
rect 1484 5866 1512 5867
rect 1536 5893 1564 5894
rect 1536 5867 1537 5893
rect 1537 5867 1563 5893
rect 1563 5867 1564 5893
rect 1536 5866 1564 5867
rect 3084 5893 3112 5894
rect 3084 5867 3085 5893
rect 3085 5867 3111 5893
rect 3111 5867 3112 5893
rect 3084 5866 3112 5867
rect 3136 5893 3164 5894
rect 3136 5867 3137 5893
rect 3137 5867 3163 5893
rect 3163 5867 3164 5893
rect 3136 5866 3164 5867
rect 3188 5893 3216 5894
rect 3188 5867 3189 5893
rect 3189 5867 3215 5893
rect 3215 5867 3216 5893
rect 3188 5866 3216 5867
rect 4736 5893 4764 5894
rect 4736 5867 4737 5893
rect 4737 5867 4763 5893
rect 4763 5867 4764 5893
rect 4736 5866 4764 5867
rect 4788 5893 4816 5894
rect 4788 5867 4789 5893
rect 4789 5867 4815 5893
rect 4815 5867 4816 5893
rect 4788 5866 4816 5867
rect 4840 5893 4868 5894
rect 4840 5867 4841 5893
rect 4841 5867 4867 5893
rect 4867 5867 4868 5893
rect 4840 5866 4868 5867
rect 6388 5893 6416 5894
rect 6388 5867 6389 5893
rect 6389 5867 6415 5893
rect 6415 5867 6416 5893
rect 6388 5866 6416 5867
rect 6440 5893 6468 5894
rect 6440 5867 6441 5893
rect 6441 5867 6467 5893
rect 6467 5867 6468 5893
rect 6440 5866 6468 5867
rect 6492 5893 6520 5894
rect 6492 5867 6493 5893
rect 6493 5867 6519 5893
rect 6519 5867 6520 5893
rect 6492 5866 6520 5867
rect 2258 5501 2286 5502
rect 2258 5475 2259 5501
rect 2259 5475 2285 5501
rect 2285 5475 2286 5501
rect 2258 5474 2286 5475
rect 2310 5501 2338 5502
rect 2310 5475 2311 5501
rect 2311 5475 2337 5501
rect 2337 5475 2338 5501
rect 2310 5474 2338 5475
rect 2362 5501 2390 5502
rect 2362 5475 2363 5501
rect 2363 5475 2389 5501
rect 2389 5475 2390 5501
rect 2362 5474 2390 5475
rect 1432 5109 1460 5110
rect 1432 5083 1433 5109
rect 1433 5083 1459 5109
rect 1459 5083 1460 5109
rect 1432 5082 1460 5083
rect 1484 5109 1512 5110
rect 1484 5083 1485 5109
rect 1485 5083 1511 5109
rect 1511 5083 1512 5109
rect 1484 5082 1512 5083
rect 1536 5109 1564 5110
rect 1536 5083 1537 5109
rect 1537 5083 1563 5109
rect 1563 5083 1564 5109
rect 1536 5082 1564 5083
rect 3084 5109 3112 5110
rect 3084 5083 3085 5109
rect 3085 5083 3111 5109
rect 3111 5083 3112 5109
rect 3084 5082 3112 5083
rect 3136 5109 3164 5110
rect 3136 5083 3137 5109
rect 3137 5083 3163 5109
rect 3163 5083 3164 5109
rect 3136 5082 3164 5083
rect 3188 5109 3216 5110
rect 3188 5083 3189 5109
rect 3189 5083 3215 5109
rect 3215 5083 3216 5109
rect 3188 5082 3216 5083
rect 3910 5501 3938 5502
rect 3910 5475 3911 5501
rect 3911 5475 3937 5501
rect 3937 5475 3938 5501
rect 3910 5474 3938 5475
rect 3962 5501 3990 5502
rect 3962 5475 3963 5501
rect 3963 5475 3989 5501
rect 3989 5475 3990 5501
rect 3962 5474 3990 5475
rect 4014 5501 4042 5502
rect 4014 5475 4015 5501
rect 4015 5475 4041 5501
rect 4041 5475 4042 5501
rect 4014 5474 4042 5475
rect 3766 5222 3794 5250
rect 4270 5334 4298 5362
rect 3542 4942 3570 4970
rect 4102 4942 4130 4970
rect 2982 4886 3010 4914
rect 2258 4717 2286 4718
rect 2258 4691 2259 4717
rect 2259 4691 2285 4717
rect 2285 4691 2286 4717
rect 2258 4690 2286 4691
rect 2310 4717 2338 4718
rect 2310 4691 2311 4717
rect 2311 4691 2337 4717
rect 2337 4691 2338 4717
rect 2310 4690 2338 4691
rect 2362 4717 2390 4718
rect 2362 4691 2363 4717
rect 2363 4691 2389 4717
rect 2389 4691 2390 4717
rect 2362 4690 2390 4691
rect 854 4382 882 4410
rect 2478 4550 2506 4578
rect 1246 4382 1274 4410
rect 1432 4325 1460 4326
rect 1432 4299 1433 4325
rect 1433 4299 1459 4325
rect 1459 4299 1460 4325
rect 1432 4298 1460 4299
rect 1484 4325 1512 4326
rect 1484 4299 1485 4325
rect 1485 4299 1511 4325
rect 1511 4299 1512 4325
rect 1484 4298 1512 4299
rect 1536 4325 1564 4326
rect 1536 4299 1537 4325
rect 1537 4299 1563 4325
rect 1563 4299 1564 4325
rect 1536 4298 1564 4299
rect 2258 3933 2286 3934
rect 2258 3907 2259 3933
rect 2259 3907 2285 3933
rect 2285 3907 2286 3933
rect 2258 3906 2286 3907
rect 2310 3933 2338 3934
rect 2310 3907 2311 3933
rect 2311 3907 2337 3933
rect 2337 3907 2338 3933
rect 2310 3906 2338 3907
rect 2362 3933 2390 3934
rect 2362 3907 2363 3933
rect 2363 3907 2389 3933
rect 2389 3907 2390 3933
rect 2362 3906 2390 3907
rect 2870 4550 2898 4578
rect 2758 4214 2786 4242
rect 2590 4129 2618 4130
rect 2590 4103 2591 4129
rect 2591 4103 2617 4129
rect 2617 4103 2618 4129
rect 2590 4102 2618 4103
rect 3486 4913 3514 4914
rect 3486 4887 3487 4913
rect 3487 4887 3513 4913
rect 3513 4887 3514 4913
rect 3486 4886 3514 4887
rect 3084 4325 3112 4326
rect 3084 4299 3085 4325
rect 3085 4299 3111 4325
rect 3111 4299 3112 4325
rect 3084 4298 3112 4299
rect 3136 4325 3164 4326
rect 3136 4299 3137 4325
rect 3137 4299 3163 4325
rect 3163 4299 3164 4325
rect 3136 4298 3164 4299
rect 3188 4325 3216 4326
rect 3188 4299 3189 4325
rect 3189 4299 3215 4325
rect 3215 4299 3216 4325
rect 3188 4298 3216 4299
rect 3206 4129 3234 4130
rect 3206 4103 3207 4129
rect 3207 4103 3233 4129
rect 3233 4103 3234 4129
rect 3206 4102 3234 4103
rect 1022 3598 1050 3626
rect 2030 3710 2058 3738
rect 1432 3541 1460 3542
rect 1432 3515 1433 3541
rect 1433 3515 1459 3541
rect 1459 3515 1460 3541
rect 1432 3514 1460 3515
rect 1484 3541 1512 3542
rect 1484 3515 1485 3541
rect 1485 3515 1511 3541
rect 1511 3515 1512 3541
rect 1484 3514 1512 3515
rect 1536 3541 1564 3542
rect 1536 3515 1537 3541
rect 1537 3515 1563 3541
rect 1563 3515 1564 3541
rect 1536 3514 1564 3515
rect 1078 3401 1106 3402
rect 1078 3375 1079 3401
rect 1079 3375 1105 3401
rect 1105 3375 1106 3401
rect 1078 3374 1106 3375
rect 1470 3374 1498 3402
rect 1022 3262 1050 3290
rect 854 3038 882 3066
rect 1246 3065 1274 3066
rect 1246 3039 1247 3065
rect 1247 3039 1273 3065
rect 1273 3039 1274 3065
rect 1246 3038 1274 3039
rect 1432 2757 1460 2758
rect 1432 2731 1433 2757
rect 1433 2731 1459 2757
rect 1459 2731 1460 2757
rect 1432 2730 1460 2731
rect 1484 2757 1512 2758
rect 1484 2731 1485 2757
rect 1485 2731 1511 2757
rect 1511 2731 1512 2757
rect 1484 2730 1512 2731
rect 1536 2757 1564 2758
rect 1536 2731 1537 2757
rect 1537 2731 1563 2757
rect 1563 2731 1564 2757
rect 1536 2730 1564 2731
rect 2198 3598 2226 3626
rect 3084 3541 3112 3542
rect 3084 3515 3085 3541
rect 3085 3515 3111 3541
rect 3111 3515 3112 3541
rect 3084 3514 3112 3515
rect 3136 3541 3164 3542
rect 3136 3515 3137 3541
rect 3137 3515 3163 3541
rect 3163 3515 3164 3541
rect 3136 3514 3164 3515
rect 3188 3541 3216 3542
rect 3188 3515 3189 3541
rect 3189 3515 3215 3541
rect 3215 3515 3216 3541
rect 3188 3514 3216 3515
rect 2366 3374 2394 3402
rect 2478 3262 2506 3290
rect 2814 3262 2842 3290
rect 2258 3149 2286 3150
rect 2258 3123 2259 3149
rect 2259 3123 2285 3149
rect 2285 3123 2286 3149
rect 2258 3122 2286 3123
rect 2310 3149 2338 3150
rect 2310 3123 2311 3149
rect 2311 3123 2337 3149
rect 2337 3123 2338 3149
rect 2310 3122 2338 3123
rect 2362 3149 2390 3150
rect 2362 3123 2363 3149
rect 2363 3123 2389 3149
rect 2389 3123 2390 3149
rect 2362 3122 2390 3123
rect 2030 2646 2058 2674
rect 2258 2365 2286 2366
rect 2258 2339 2259 2365
rect 2259 2339 2285 2365
rect 2285 2339 2286 2365
rect 2258 2338 2286 2339
rect 2310 2365 2338 2366
rect 2310 2339 2311 2365
rect 2311 2339 2337 2365
rect 2337 2339 2338 2365
rect 2310 2338 2338 2339
rect 2362 2365 2390 2366
rect 2362 2339 2363 2365
rect 2363 2339 2389 2365
rect 2389 2339 2390 2365
rect 2362 2338 2390 2339
rect 1432 1973 1460 1974
rect 1432 1947 1433 1973
rect 1433 1947 1459 1973
rect 1459 1947 1460 1973
rect 1432 1946 1460 1947
rect 1484 1973 1512 1974
rect 1484 1947 1485 1973
rect 1485 1947 1511 1973
rect 1511 1947 1512 1973
rect 1484 1946 1512 1947
rect 1536 1973 1564 1974
rect 1536 1947 1537 1973
rect 1537 1947 1563 1973
rect 1563 1947 1564 1973
rect 1536 1946 1564 1947
rect 2258 1581 2286 1582
rect 2258 1555 2259 1581
rect 2259 1555 2285 1581
rect 2285 1555 2286 1581
rect 2258 1554 2286 1555
rect 2310 1581 2338 1582
rect 2310 1555 2311 1581
rect 2311 1555 2337 1581
rect 2337 1555 2338 1581
rect 2310 1554 2338 1555
rect 2362 1581 2390 1582
rect 2362 1555 2363 1581
rect 2363 1555 2389 1581
rect 2389 1555 2390 1581
rect 2362 1554 2390 1555
rect 3084 2757 3112 2758
rect 3084 2731 3085 2757
rect 3085 2731 3111 2757
rect 3111 2731 3112 2757
rect 3084 2730 3112 2731
rect 3136 2757 3164 2758
rect 3136 2731 3137 2757
rect 3137 2731 3163 2757
rect 3163 2731 3164 2757
rect 3136 2730 3164 2731
rect 3188 2757 3216 2758
rect 3188 2731 3189 2757
rect 3189 2731 3215 2757
rect 3215 2731 3216 2757
rect 3188 2730 3216 2731
rect 3038 2646 3066 2674
rect 3910 4717 3938 4718
rect 3910 4691 3911 4717
rect 3911 4691 3937 4717
rect 3937 4691 3938 4717
rect 3910 4690 3938 4691
rect 3962 4717 3990 4718
rect 3962 4691 3963 4717
rect 3963 4691 3989 4717
rect 3989 4691 3990 4717
rect 3962 4690 3990 4691
rect 4014 4717 4042 4718
rect 4014 4691 4015 4717
rect 4015 4691 4041 4717
rect 4041 4691 4042 4717
rect 4014 4690 4042 4691
rect 3878 4577 3906 4578
rect 3878 4551 3879 4577
rect 3879 4551 3905 4577
rect 3905 4551 3906 4577
rect 3878 4550 3906 4551
rect 3910 3933 3938 3934
rect 3910 3907 3911 3933
rect 3911 3907 3937 3933
rect 3937 3907 3938 3933
rect 3910 3906 3938 3907
rect 3962 3933 3990 3934
rect 3962 3907 3963 3933
rect 3963 3907 3989 3933
rect 3989 3907 3990 3933
rect 3962 3906 3990 3907
rect 4014 3933 4042 3934
rect 4014 3907 4015 3933
rect 4015 3907 4041 3933
rect 4041 3907 4042 3933
rect 4014 3906 4042 3907
rect 5278 5361 5306 5362
rect 5278 5335 5279 5361
rect 5279 5335 5305 5361
rect 5305 5335 5306 5361
rect 5278 5334 5306 5335
rect 4774 5249 4802 5250
rect 4774 5223 4775 5249
rect 4775 5223 4801 5249
rect 4801 5223 4802 5249
rect 4774 5222 4802 5223
rect 4736 5109 4764 5110
rect 4736 5083 4737 5109
rect 4737 5083 4763 5109
rect 4763 5083 4764 5109
rect 4736 5082 4764 5083
rect 4788 5109 4816 5110
rect 4788 5083 4789 5109
rect 4789 5083 4815 5109
rect 4815 5083 4816 5109
rect 4788 5082 4816 5083
rect 4840 5109 4868 5110
rect 4840 5083 4841 5109
rect 4841 5083 4867 5109
rect 4867 5083 4868 5109
rect 4840 5082 4868 5083
rect 4830 4969 4858 4970
rect 4830 4943 4831 4969
rect 4831 4943 4857 4969
rect 4857 4943 4858 4969
rect 4830 4942 4858 4943
rect 4326 4886 4354 4914
rect 5562 5501 5590 5502
rect 5562 5475 5563 5501
rect 5563 5475 5589 5501
rect 5589 5475 5590 5501
rect 5562 5474 5590 5475
rect 5614 5501 5642 5502
rect 5614 5475 5615 5501
rect 5615 5475 5641 5501
rect 5641 5475 5642 5501
rect 5614 5474 5642 5475
rect 5666 5501 5694 5502
rect 5666 5475 5667 5501
rect 5667 5475 5693 5501
rect 5693 5475 5694 5501
rect 5666 5474 5694 5475
rect 7214 5501 7242 5502
rect 7214 5475 7215 5501
rect 7215 5475 7241 5501
rect 7241 5475 7242 5501
rect 7214 5474 7242 5475
rect 7266 5501 7294 5502
rect 7266 5475 7267 5501
rect 7267 5475 7293 5501
rect 7293 5475 7294 5501
rect 7266 5474 7294 5475
rect 7318 5501 7346 5502
rect 7318 5475 7319 5501
rect 7319 5475 7345 5501
rect 7345 5475 7346 5501
rect 7318 5474 7346 5475
rect 6388 5109 6416 5110
rect 6388 5083 6389 5109
rect 6389 5083 6415 5109
rect 6415 5083 6416 5109
rect 6388 5082 6416 5083
rect 6440 5109 6468 5110
rect 6440 5083 6441 5109
rect 6441 5083 6467 5109
rect 6467 5083 6468 5109
rect 6440 5082 6468 5083
rect 6492 5109 6520 5110
rect 6492 5083 6493 5109
rect 6493 5083 6519 5109
rect 6519 5083 6520 5109
rect 6492 5082 6520 5083
rect 5562 4717 5590 4718
rect 5562 4691 5563 4717
rect 5563 4691 5589 4717
rect 5589 4691 5590 4717
rect 5562 4690 5590 4691
rect 5614 4717 5642 4718
rect 5614 4691 5615 4717
rect 5615 4691 5641 4717
rect 5641 4691 5642 4717
rect 5614 4690 5642 4691
rect 5666 4717 5694 4718
rect 5666 4691 5667 4717
rect 5667 4691 5693 4717
rect 5693 4691 5694 4717
rect 5666 4690 5694 4691
rect 7214 4717 7242 4718
rect 7214 4691 7215 4717
rect 7215 4691 7241 4717
rect 7241 4691 7242 4717
rect 7214 4690 7242 4691
rect 7266 4717 7294 4718
rect 7266 4691 7267 4717
rect 7267 4691 7293 4717
rect 7293 4691 7294 4717
rect 7266 4690 7294 4691
rect 7318 4717 7346 4718
rect 7318 4691 7319 4717
rect 7319 4691 7345 4717
rect 7345 4691 7346 4717
rect 7318 4690 7346 4691
rect 7014 4606 7042 4634
rect 5334 4550 5362 4578
rect 5894 4577 5922 4578
rect 5894 4551 5895 4577
rect 5895 4551 5921 4577
rect 5921 4551 5922 4577
rect 5894 4550 5922 4551
rect 4736 4325 4764 4326
rect 4736 4299 4737 4325
rect 4737 4299 4763 4325
rect 4763 4299 4764 4325
rect 4736 4298 4764 4299
rect 4788 4325 4816 4326
rect 4788 4299 4789 4325
rect 4789 4299 4815 4325
rect 4815 4299 4816 4325
rect 4788 4298 4816 4299
rect 4840 4325 4868 4326
rect 4840 4299 4841 4325
rect 4841 4299 4867 4325
rect 4867 4299 4868 4325
rect 4840 4298 4868 4299
rect 5278 4214 5306 4242
rect 4382 4102 4410 4130
rect 4382 3766 4410 3794
rect 4998 3710 5026 3738
rect 4736 3541 4764 3542
rect 4736 3515 4737 3541
rect 4737 3515 4763 3541
rect 4763 3515 4764 3541
rect 4736 3514 4764 3515
rect 4788 3541 4816 3542
rect 4788 3515 4789 3541
rect 4789 3515 4815 3541
rect 4815 3515 4816 3541
rect 4788 3514 4816 3515
rect 4840 3541 4868 3542
rect 4840 3515 4841 3541
rect 4841 3515 4867 3541
rect 4867 3515 4868 3541
rect 4840 3514 4868 3515
rect 3084 1973 3112 1974
rect 3084 1947 3085 1973
rect 3085 1947 3111 1973
rect 3111 1947 3112 1973
rect 3084 1946 3112 1947
rect 3136 1973 3164 1974
rect 3136 1947 3137 1973
rect 3137 1947 3163 1973
rect 3163 1947 3164 1973
rect 3136 1946 3164 1947
rect 3188 1973 3216 1974
rect 3188 1947 3189 1973
rect 3189 1947 3215 1973
rect 3215 1947 3216 1973
rect 3188 1946 3216 1947
rect 3486 1806 3514 1834
rect 3910 3149 3938 3150
rect 3910 3123 3911 3149
rect 3911 3123 3937 3149
rect 3937 3123 3938 3149
rect 3910 3122 3938 3123
rect 3962 3149 3990 3150
rect 3962 3123 3963 3149
rect 3963 3123 3989 3149
rect 3989 3123 3990 3149
rect 3962 3122 3990 3123
rect 4014 3149 4042 3150
rect 4014 3123 4015 3149
rect 4015 3123 4041 3149
rect 4041 3123 4042 3149
rect 4014 3122 4042 3123
rect 4830 3206 4858 3234
rect 3878 2841 3906 2842
rect 3878 2815 3879 2841
rect 3879 2815 3905 2841
rect 3905 2815 3906 2841
rect 3878 2814 3906 2815
rect 3910 2365 3938 2366
rect 3910 2339 3911 2365
rect 3911 2339 3937 2365
rect 3937 2339 3938 2365
rect 3910 2338 3938 2339
rect 3962 2365 3990 2366
rect 3962 2339 3963 2365
rect 3963 2339 3989 2365
rect 3989 2339 3990 2365
rect 3962 2338 3990 2339
rect 4014 2365 4042 2366
rect 4014 2339 4015 2365
rect 4015 2339 4041 2365
rect 4041 2339 4042 2365
rect 4014 2338 4042 2339
rect 3598 1918 3626 1946
rect 3766 1833 3794 1834
rect 3766 1807 3767 1833
rect 3767 1807 3793 1833
rect 3793 1807 3794 1833
rect 3766 1806 3794 1807
rect 4102 1806 4130 1834
rect 3910 1581 3938 1582
rect 3910 1555 3911 1581
rect 3911 1555 3937 1581
rect 3937 1555 3938 1581
rect 3910 1554 3938 1555
rect 3962 1581 3990 1582
rect 3962 1555 3963 1581
rect 3963 1555 3989 1581
rect 3989 1555 3990 1581
rect 3962 1554 3990 1555
rect 4014 1581 4042 1582
rect 4014 1555 4015 1581
rect 4015 1555 4041 1581
rect 4041 1555 4042 1581
rect 4014 1554 4042 1555
rect 4736 2757 4764 2758
rect 4736 2731 4737 2757
rect 4737 2731 4763 2757
rect 4763 2731 4764 2757
rect 4736 2730 4764 2731
rect 4788 2757 4816 2758
rect 4788 2731 4789 2757
rect 4789 2731 4815 2757
rect 4815 2731 4816 2757
rect 4788 2730 4816 2731
rect 4840 2757 4868 2758
rect 4840 2731 4841 2757
rect 4841 2731 4867 2757
rect 4867 2731 4868 2757
rect 4840 2730 4868 2731
rect 5166 3654 5194 3682
rect 6388 4325 6416 4326
rect 6388 4299 6389 4325
rect 6389 4299 6415 4325
rect 6415 4299 6416 4325
rect 6388 4298 6416 4299
rect 6440 4325 6468 4326
rect 6440 4299 6441 4325
rect 6441 4299 6467 4325
rect 6467 4299 6468 4325
rect 6440 4298 6468 4299
rect 6492 4325 6520 4326
rect 6492 4299 6493 4325
rect 6493 4299 6519 4325
rect 6519 4299 6520 4325
rect 6492 4298 6520 4299
rect 5562 3933 5590 3934
rect 5562 3907 5563 3933
rect 5563 3907 5589 3933
rect 5589 3907 5590 3933
rect 5562 3906 5590 3907
rect 5614 3933 5642 3934
rect 5614 3907 5615 3933
rect 5615 3907 5641 3933
rect 5641 3907 5642 3933
rect 5614 3906 5642 3907
rect 5666 3933 5694 3934
rect 5666 3907 5667 3933
rect 5667 3907 5693 3933
rect 5693 3907 5694 3933
rect 5666 3906 5694 3907
rect 5390 3766 5418 3794
rect 5614 3598 5642 3626
rect 6510 4185 6538 4186
rect 6510 4159 6511 4185
rect 6511 4159 6537 4185
rect 6537 4159 6538 4185
rect 6510 4158 6538 4159
rect 7070 4158 7098 4186
rect 6118 4129 6146 4130
rect 6118 4103 6119 4129
rect 6119 4103 6145 4129
rect 6145 4103 6146 4129
rect 6118 4102 6146 4103
rect 6790 4129 6818 4130
rect 6790 4103 6791 4129
rect 6791 4103 6817 4129
rect 6817 4103 6818 4129
rect 6790 4102 6818 4103
rect 5562 3149 5590 3150
rect 5562 3123 5563 3149
rect 5563 3123 5589 3149
rect 5589 3123 5590 3149
rect 5562 3122 5590 3123
rect 5614 3149 5642 3150
rect 5614 3123 5615 3149
rect 5615 3123 5641 3149
rect 5641 3123 5642 3149
rect 5614 3122 5642 3123
rect 5666 3149 5694 3150
rect 5666 3123 5667 3149
rect 5667 3123 5693 3149
rect 5693 3123 5694 3149
rect 5666 3122 5694 3123
rect 7214 3933 7242 3934
rect 7214 3907 7215 3933
rect 7215 3907 7241 3933
rect 7241 3907 7242 3933
rect 7214 3906 7242 3907
rect 7266 3933 7294 3934
rect 7266 3907 7267 3933
rect 7267 3907 7293 3933
rect 7293 3907 7294 3933
rect 7266 3906 7294 3907
rect 7318 3933 7346 3934
rect 7318 3907 7319 3933
rect 7319 3907 7345 3933
rect 7345 3907 7346 3933
rect 7318 3906 7346 3907
rect 6454 3737 6482 3738
rect 6454 3711 6455 3737
rect 6455 3711 6481 3737
rect 6481 3711 6482 3737
rect 6454 3710 6482 3711
rect 6006 3598 6034 3626
rect 6388 3541 6416 3542
rect 6388 3515 6389 3541
rect 6389 3515 6415 3541
rect 6415 3515 6416 3541
rect 6388 3514 6416 3515
rect 6440 3541 6468 3542
rect 6440 3515 6441 3541
rect 6441 3515 6467 3541
rect 6467 3515 6468 3541
rect 6440 3514 6468 3515
rect 6492 3541 6520 3542
rect 6492 3515 6493 3541
rect 6493 3515 6519 3541
rect 6519 3515 6520 3541
rect 6492 3514 6520 3515
rect 7014 3374 7042 3402
rect 6902 3233 6930 3234
rect 6902 3207 6903 3233
rect 6903 3207 6929 3233
rect 6929 3207 6930 3233
rect 6902 3206 6930 3207
rect 7214 3149 7242 3150
rect 7214 3123 7215 3149
rect 7215 3123 7241 3149
rect 7241 3123 7242 3149
rect 7214 3122 7242 3123
rect 7266 3149 7294 3150
rect 7266 3123 7267 3149
rect 7267 3123 7293 3149
rect 7293 3123 7294 3149
rect 7266 3122 7294 3123
rect 7318 3149 7346 3150
rect 7318 3123 7319 3149
rect 7319 3123 7345 3149
rect 7345 3123 7346 3149
rect 7318 3122 7346 3123
rect 7126 3065 7154 3066
rect 7126 3039 7127 3065
rect 7127 3039 7153 3065
rect 7153 3039 7154 3065
rect 7126 3038 7154 3039
rect 5950 2814 5978 2842
rect 6388 2757 6416 2758
rect 6388 2731 6389 2757
rect 6389 2731 6415 2757
rect 6415 2731 6416 2757
rect 6388 2730 6416 2731
rect 6440 2757 6468 2758
rect 6440 2731 6441 2757
rect 6441 2731 6467 2757
rect 6467 2731 6468 2757
rect 6440 2730 6468 2731
rect 6492 2757 6520 2758
rect 6492 2731 6493 2757
rect 6493 2731 6519 2757
rect 6519 2731 6520 2757
rect 6492 2730 6520 2731
rect 5562 2365 5590 2366
rect 5562 2339 5563 2365
rect 5563 2339 5589 2365
rect 5589 2339 5590 2365
rect 5562 2338 5590 2339
rect 5614 2365 5642 2366
rect 5614 2339 5615 2365
rect 5615 2339 5641 2365
rect 5641 2339 5642 2365
rect 5614 2338 5642 2339
rect 5666 2365 5694 2366
rect 5666 2339 5667 2365
rect 5667 2339 5693 2365
rect 5693 2339 5694 2365
rect 5666 2338 5694 2339
rect 7214 2365 7242 2366
rect 7214 2339 7215 2365
rect 7215 2339 7241 2365
rect 7241 2339 7242 2365
rect 7214 2338 7242 2339
rect 7266 2365 7294 2366
rect 7266 2339 7267 2365
rect 7267 2339 7293 2365
rect 7293 2339 7294 2365
rect 7266 2338 7294 2339
rect 7318 2365 7346 2366
rect 7318 2339 7319 2365
rect 7319 2339 7345 2365
rect 7345 2339 7346 2365
rect 7318 2338 7346 2339
rect 4736 1973 4764 1974
rect 4158 1750 4186 1778
rect 4382 1918 4410 1946
rect 4736 1947 4737 1973
rect 4737 1947 4763 1973
rect 4763 1947 4764 1973
rect 4736 1946 4764 1947
rect 4788 1973 4816 1974
rect 4788 1947 4789 1973
rect 4789 1947 4815 1973
rect 4815 1947 4816 1973
rect 4788 1946 4816 1947
rect 4840 1973 4868 1974
rect 4840 1947 4841 1973
rect 4841 1947 4867 1973
rect 4867 1947 4868 1973
rect 4840 1946 4868 1947
rect 6388 1973 6416 1974
rect 6388 1947 6389 1973
rect 6389 1947 6415 1973
rect 6415 1947 6416 1973
rect 6388 1946 6416 1947
rect 6440 1973 6468 1974
rect 6440 1947 6441 1973
rect 6441 1947 6467 1973
rect 6467 1947 6468 1973
rect 6440 1946 6468 1947
rect 6492 1973 6520 1974
rect 6492 1947 6493 1973
rect 6493 1947 6519 1973
rect 6519 1947 6520 1973
rect 6492 1946 6520 1947
rect 4886 1833 4914 1834
rect 4886 1807 4887 1833
rect 4887 1807 4913 1833
rect 4913 1807 4914 1833
rect 4886 1806 4914 1807
rect 4662 1777 4690 1778
rect 4662 1751 4663 1777
rect 4663 1751 4689 1777
rect 4689 1751 4690 1777
rect 4662 1750 4690 1751
rect 5562 1581 5590 1582
rect 5562 1555 5563 1581
rect 5563 1555 5589 1581
rect 5589 1555 5590 1581
rect 5562 1554 5590 1555
rect 5614 1581 5642 1582
rect 5614 1555 5615 1581
rect 5615 1555 5641 1581
rect 5641 1555 5642 1581
rect 5614 1554 5642 1555
rect 5666 1581 5694 1582
rect 5666 1555 5667 1581
rect 5667 1555 5693 1581
rect 5693 1555 5694 1581
rect 5666 1554 5694 1555
rect 7214 1581 7242 1582
rect 7214 1555 7215 1581
rect 7215 1555 7241 1581
rect 7241 1555 7242 1581
rect 7214 1554 7242 1555
rect 7266 1581 7294 1582
rect 7266 1555 7267 1581
rect 7267 1555 7293 1581
rect 7293 1555 7294 1581
rect 7266 1554 7294 1555
rect 7318 1581 7346 1582
rect 7318 1555 7319 1581
rect 7319 1555 7345 1581
rect 7345 1555 7346 1581
rect 7318 1554 7346 1555
<< metal3 >>
rect 2253 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2395 6286
rect 3905 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4047 6286
rect 5557 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5699 6286
rect 7209 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7351 6286
rect 1427 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1569 5894
rect 3079 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3221 5894
rect 4731 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4873 5894
rect 6383 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6525 5894
rect 2253 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2395 5502
rect 3905 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4047 5502
rect 5557 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5699 5502
rect 7209 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7351 5502
rect 4265 5334 4270 5362
rect 4298 5334 5278 5362
rect 5306 5334 5311 5362
rect 3761 5222 3766 5250
rect 3794 5222 4774 5250
rect 4802 5222 4807 5250
rect 1427 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1569 5110
rect 3079 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3221 5110
rect 4731 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4873 5110
rect 6383 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6525 5110
rect 3537 4942 3542 4970
rect 3570 4942 4102 4970
rect 4130 4942 4830 4970
rect 4858 4942 4863 4970
rect 2977 4886 2982 4914
rect 3010 4886 3486 4914
rect 3514 4886 4326 4914
rect 4354 4886 4359 4914
rect 0 4746 400 4760
rect 7600 4746 8000 4760
rect 0 4718 1694 4746
rect 7406 4718 8000 4746
rect 0 4704 400 4718
rect 1666 4578 1694 4718
rect 2253 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2395 4718
rect 3905 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4047 4718
rect 5557 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5699 4718
rect 7209 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7351 4718
rect 7406 4634 7434 4718
rect 7600 4704 8000 4718
rect 7009 4606 7014 4634
rect 7042 4606 7434 4634
rect 1666 4550 2478 4578
rect 2506 4550 2511 4578
rect 2865 4550 2870 4578
rect 2898 4550 3878 4578
rect 3906 4550 3911 4578
rect 5329 4550 5334 4578
rect 5362 4550 5894 4578
rect 5922 4550 5927 4578
rect 0 4410 400 4424
rect 7600 4410 8000 4424
rect 0 4382 854 4410
rect 882 4382 1246 4410
rect 1274 4382 1279 4410
rect 7518 4382 8000 4410
rect 0 4368 400 4382
rect 1427 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1569 4326
rect 3079 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3221 4326
rect 4731 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4873 4326
rect 6383 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6525 4326
rect 7518 4242 7546 4382
rect 7600 4368 8000 4382
rect 2753 4214 2758 4242
rect 2786 4214 5278 4242
rect 5306 4214 5311 4242
rect 7518 4214 7658 4242
rect 7630 4186 7658 4214
rect 6505 4158 6510 4186
rect 6538 4158 7070 4186
rect 7098 4158 7658 4186
rect 2585 4102 2590 4130
rect 2618 4102 3206 4130
rect 3234 4102 3239 4130
rect 4377 4102 4382 4130
rect 4410 4102 6118 4130
rect 6146 4102 6790 4130
rect 6818 4102 6823 4130
rect 2253 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2395 3934
rect 3905 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4047 3934
rect 5557 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5699 3934
rect 7209 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7351 3934
rect 4377 3766 4382 3794
rect 4410 3766 5390 3794
rect 5418 3766 5423 3794
rect 0 3738 400 3752
rect 7600 3738 8000 3752
rect 0 3710 2030 3738
rect 2058 3710 2063 3738
rect 4993 3710 4998 3738
rect 5026 3710 6454 3738
rect 6482 3710 6487 3738
rect 6566 3710 8000 3738
rect 0 3696 400 3710
rect 6566 3682 6594 3710
rect 7600 3696 8000 3710
rect 5161 3654 5166 3682
rect 5194 3654 6594 3682
rect 1017 3598 1022 3626
rect 1050 3598 2198 3626
rect 2226 3598 2231 3626
rect 5609 3598 5614 3626
rect 5642 3598 6006 3626
rect 6034 3598 6039 3626
rect 1427 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1569 3542
rect 3079 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3221 3542
rect 4731 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4873 3542
rect 6383 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6525 3542
rect 0 3402 400 3416
rect 7600 3402 8000 3416
rect 0 3374 1078 3402
rect 1106 3374 1111 3402
rect 1465 3374 1470 3402
rect 1498 3374 2366 3402
rect 2394 3374 2399 3402
rect 7009 3374 7014 3402
rect 7042 3374 8000 3402
rect 0 3360 400 3374
rect 7600 3360 8000 3374
rect 1017 3262 1022 3290
rect 1050 3262 2478 3290
rect 2506 3262 2814 3290
rect 2842 3262 2847 3290
rect 4825 3206 4830 3234
rect 4858 3206 6902 3234
rect 6930 3206 6935 3234
rect 2253 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2395 3150
rect 3905 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4047 3150
rect 5557 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5699 3150
rect 7209 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7351 3150
rect 0 3066 400 3080
rect 7600 3066 8000 3080
rect 0 3038 854 3066
rect 882 3038 1246 3066
rect 1274 3038 1279 3066
rect 7121 3038 7126 3066
rect 7154 3038 8000 3066
rect 0 3024 400 3038
rect 7600 3024 8000 3038
rect 3873 2814 3878 2842
rect 3906 2814 5950 2842
rect 5978 2814 5983 2842
rect 1427 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1569 2758
rect 3079 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3221 2758
rect 4731 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4873 2758
rect 6383 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6525 2758
rect 2025 2646 2030 2674
rect 2058 2646 3038 2674
rect 3066 2646 3071 2674
rect 2253 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2395 2366
rect 3905 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4047 2366
rect 5557 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5699 2366
rect 7209 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7351 2366
rect 1427 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1569 1974
rect 3079 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3221 1974
rect 4731 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4873 1974
rect 6383 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6525 1974
rect 3593 1918 3598 1946
rect 3626 1918 4382 1946
rect 4410 1918 4415 1946
rect 3481 1806 3486 1834
rect 3514 1806 3766 1834
rect 3794 1806 3799 1834
rect 4097 1806 4102 1834
rect 4130 1806 4886 1834
rect 4914 1806 4919 1834
rect 4153 1750 4158 1778
rect 4186 1750 4662 1778
rect 4690 1750 4695 1778
rect 2253 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2395 1582
rect 3905 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4047 1582
rect 5557 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5699 1582
rect 7209 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7351 1582
<< via3 >>
rect 2258 6258 2286 6286
rect 2310 6258 2338 6286
rect 2362 6258 2390 6286
rect 3910 6258 3938 6286
rect 3962 6258 3990 6286
rect 4014 6258 4042 6286
rect 5562 6258 5590 6286
rect 5614 6258 5642 6286
rect 5666 6258 5694 6286
rect 7214 6258 7242 6286
rect 7266 6258 7294 6286
rect 7318 6258 7346 6286
rect 1432 5866 1460 5894
rect 1484 5866 1512 5894
rect 1536 5866 1564 5894
rect 3084 5866 3112 5894
rect 3136 5866 3164 5894
rect 3188 5866 3216 5894
rect 4736 5866 4764 5894
rect 4788 5866 4816 5894
rect 4840 5866 4868 5894
rect 6388 5866 6416 5894
rect 6440 5866 6468 5894
rect 6492 5866 6520 5894
rect 2258 5474 2286 5502
rect 2310 5474 2338 5502
rect 2362 5474 2390 5502
rect 3910 5474 3938 5502
rect 3962 5474 3990 5502
rect 4014 5474 4042 5502
rect 5562 5474 5590 5502
rect 5614 5474 5642 5502
rect 5666 5474 5694 5502
rect 7214 5474 7242 5502
rect 7266 5474 7294 5502
rect 7318 5474 7346 5502
rect 1432 5082 1460 5110
rect 1484 5082 1512 5110
rect 1536 5082 1564 5110
rect 3084 5082 3112 5110
rect 3136 5082 3164 5110
rect 3188 5082 3216 5110
rect 4736 5082 4764 5110
rect 4788 5082 4816 5110
rect 4840 5082 4868 5110
rect 6388 5082 6416 5110
rect 6440 5082 6468 5110
rect 6492 5082 6520 5110
rect 2258 4690 2286 4718
rect 2310 4690 2338 4718
rect 2362 4690 2390 4718
rect 3910 4690 3938 4718
rect 3962 4690 3990 4718
rect 4014 4690 4042 4718
rect 5562 4690 5590 4718
rect 5614 4690 5642 4718
rect 5666 4690 5694 4718
rect 7214 4690 7242 4718
rect 7266 4690 7294 4718
rect 7318 4690 7346 4718
rect 1432 4298 1460 4326
rect 1484 4298 1512 4326
rect 1536 4298 1564 4326
rect 3084 4298 3112 4326
rect 3136 4298 3164 4326
rect 3188 4298 3216 4326
rect 4736 4298 4764 4326
rect 4788 4298 4816 4326
rect 4840 4298 4868 4326
rect 6388 4298 6416 4326
rect 6440 4298 6468 4326
rect 6492 4298 6520 4326
rect 2258 3906 2286 3934
rect 2310 3906 2338 3934
rect 2362 3906 2390 3934
rect 3910 3906 3938 3934
rect 3962 3906 3990 3934
rect 4014 3906 4042 3934
rect 5562 3906 5590 3934
rect 5614 3906 5642 3934
rect 5666 3906 5694 3934
rect 7214 3906 7242 3934
rect 7266 3906 7294 3934
rect 7318 3906 7346 3934
rect 1432 3514 1460 3542
rect 1484 3514 1512 3542
rect 1536 3514 1564 3542
rect 3084 3514 3112 3542
rect 3136 3514 3164 3542
rect 3188 3514 3216 3542
rect 4736 3514 4764 3542
rect 4788 3514 4816 3542
rect 4840 3514 4868 3542
rect 6388 3514 6416 3542
rect 6440 3514 6468 3542
rect 6492 3514 6520 3542
rect 2258 3122 2286 3150
rect 2310 3122 2338 3150
rect 2362 3122 2390 3150
rect 3910 3122 3938 3150
rect 3962 3122 3990 3150
rect 4014 3122 4042 3150
rect 5562 3122 5590 3150
rect 5614 3122 5642 3150
rect 5666 3122 5694 3150
rect 7214 3122 7242 3150
rect 7266 3122 7294 3150
rect 7318 3122 7346 3150
rect 1432 2730 1460 2758
rect 1484 2730 1512 2758
rect 1536 2730 1564 2758
rect 3084 2730 3112 2758
rect 3136 2730 3164 2758
rect 3188 2730 3216 2758
rect 4736 2730 4764 2758
rect 4788 2730 4816 2758
rect 4840 2730 4868 2758
rect 6388 2730 6416 2758
rect 6440 2730 6468 2758
rect 6492 2730 6520 2758
rect 2258 2338 2286 2366
rect 2310 2338 2338 2366
rect 2362 2338 2390 2366
rect 3910 2338 3938 2366
rect 3962 2338 3990 2366
rect 4014 2338 4042 2366
rect 5562 2338 5590 2366
rect 5614 2338 5642 2366
rect 5666 2338 5694 2366
rect 7214 2338 7242 2366
rect 7266 2338 7294 2366
rect 7318 2338 7346 2366
rect 1432 1946 1460 1974
rect 1484 1946 1512 1974
rect 1536 1946 1564 1974
rect 3084 1946 3112 1974
rect 3136 1946 3164 1974
rect 3188 1946 3216 1974
rect 4736 1946 4764 1974
rect 4788 1946 4816 1974
rect 4840 1946 4868 1974
rect 6388 1946 6416 1974
rect 6440 1946 6468 1974
rect 6492 1946 6520 1974
rect 2258 1554 2286 1582
rect 2310 1554 2338 1582
rect 2362 1554 2390 1582
rect 3910 1554 3938 1582
rect 3962 1554 3990 1582
rect 4014 1554 4042 1582
rect 5562 1554 5590 1582
rect 5614 1554 5642 1582
rect 5666 1554 5694 1582
rect 7214 1554 7242 1582
rect 7266 1554 7294 1582
rect 7318 1554 7346 1582
<< metal4 >>
rect 1418 5894 1578 6302
rect 1418 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1578 5894
rect 1418 5110 1578 5866
rect 1418 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1578 5110
rect 1418 4326 1578 5082
rect 1418 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1578 4326
rect 1418 3542 1578 4298
rect 1418 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1578 3542
rect 1418 2758 1578 3514
rect 1418 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1578 2758
rect 1418 1974 1578 2730
rect 1418 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1578 1974
rect 1418 1538 1578 1946
rect 2244 6286 2404 6302
rect 2244 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2404 6286
rect 2244 5502 2404 6258
rect 2244 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2404 5502
rect 2244 4718 2404 5474
rect 2244 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2404 4718
rect 2244 3934 2404 4690
rect 2244 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2404 3934
rect 2244 3150 2404 3906
rect 2244 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2404 3150
rect 2244 2366 2404 3122
rect 2244 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2404 2366
rect 2244 1582 2404 2338
rect 2244 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2404 1582
rect 2244 1538 2404 1554
rect 3070 5894 3230 6302
rect 3070 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3230 5894
rect 3070 5110 3230 5866
rect 3070 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3230 5110
rect 3070 4326 3230 5082
rect 3070 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3230 4326
rect 3070 3542 3230 4298
rect 3070 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3230 3542
rect 3070 2758 3230 3514
rect 3070 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3230 2758
rect 3070 1974 3230 2730
rect 3070 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3230 1974
rect 3070 1538 3230 1946
rect 3896 6286 4056 6302
rect 3896 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4056 6286
rect 3896 5502 4056 6258
rect 3896 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4056 5502
rect 3896 4718 4056 5474
rect 3896 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4056 4718
rect 3896 3934 4056 4690
rect 3896 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4056 3934
rect 3896 3150 4056 3906
rect 3896 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4056 3150
rect 3896 2366 4056 3122
rect 3896 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4056 2366
rect 3896 1582 4056 2338
rect 3896 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4056 1582
rect 3896 1538 4056 1554
rect 4722 5894 4882 6302
rect 4722 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4882 5894
rect 4722 5110 4882 5866
rect 4722 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4882 5110
rect 4722 4326 4882 5082
rect 4722 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4882 4326
rect 4722 3542 4882 4298
rect 4722 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4882 3542
rect 4722 2758 4882 3514
rect 4722 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4882 2758
rect 4722 1974 4882 2730
rect 4722 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4882 1974
rect 4722 1538 4882 1946
rect 5548 6286 5708 6302
rect 5548 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5708 6286
rect 5548 5502 5708 6258
rect 5548 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5708 5502
rect 5548 4718 5708 5474
rect 5548 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5708 4718
rect 5548 3934 5708 4690
rect 5548 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5708 3934
rect 5548 3150 5708 3906
rect 5548 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5708 3150
rect 5548 2366 5708 3122
rect 5548 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5708 2366
rect 5548 1582 5708 2338
rect 5548 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5708 1582
rect 5548 1538 5708 1554
rect 6374 5894 6534 6302
rect 6374 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6534 5894
rect 6374 5110 6534 5866
rect 6374 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6534 5110
rect 6374 4326 6534 5082
rect 6374 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6534 4326
rect 6374 3542 6534 4298
rect 6374 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6534 3542
rect 6374 2758 6534 3514
rect 6374 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6534 2758
rect 6374 1974 6534 2730
rect 6374 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6534 1974
rect 6374 1538 6534 1946
rect 7200 6286 7360 6302
rect 7200 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7360 6286
rect 7200 5502 7360 6258
rect 7200 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7360 5502
rect 7200 4718 7360 5474
rect 7200 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7360 4718
rect 7200 3934 7360 4690
rect 7200 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7360 3934
rect 7200 3150 7360 3906
rect 7200 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7360 3150
rect 7200 2366 7360 3122
rect 7200 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7360 2366
rect 7200 1582 7360 2338
rect 7200 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7360 1582
rect 7200 1538 7360 1554
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _04_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _05_
timestamp 1698431365
transform -1 0 3136 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _06_
timestamp 1698431365
transform 1 0 4256 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _07_
timestamp 1698431365
transform -1 0 6272 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _08_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 -1 3136
box -43 -43 1947 435
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _09_
timestamp 1698431365
transform 1 0 2408 0 -1 4704
box -43 -43 1947 435
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _10_
timestamp 1698431365
transform 1 0 3416 0 1 5488
box -43 -43 1947 435
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _11_
timestamp 1698431365
transform 1 0 4032 0 1 3136
box -43 -43 1947 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _12_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3472 0 1 3136
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _13_
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _14_
timestamp 1698431365
transform -1 0 4032 0 1 3136
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _15_
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _16_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _17_
timestamp 1698431365
transform 1 0 3920 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _18_
timestamp 1698431365
transform -1 0 2632 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _19_
timestamp 1698431365
transform 1 0 3304 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1232 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 7168 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 3752 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 1232 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 3080 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 1 3920
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1698431365
transform -1 0 4312 0 -1 3920
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1698431365
transform 1 0 3752 0 1 4704
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_40 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_59 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3976 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 4424 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_80 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_96
timestamp 1698431365
transform 1 0 6048 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_100 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_104
timestamp 1698431365
transform 1 0 6496 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_112
timestamp 1698431365
transform 1 0 6944 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_2
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_34
timestamp 1698431365
transform 1 0 2576 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_50
timestamp 1698431365
transform 1 0 3472 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_52
timestamp 1698431365
transform 1 0 3584 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_61
timestamp 1698431365
transform 1 0 4088 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 4536 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_104
timestamp 1698431365
transform 1 0 6496 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_112
timestamp 1698431365
transform 1 0 6944 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_53
timestamp 1698431365
transform 1 0 3640 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_69
timestamp 1698431365
transform 1 0 4536 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_71
timestamp 1698431365
transform 1 0 4648 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_78
timestamp 1698431365
transform 1 0 5040 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_94
timestamp 1698431365
transform 1 0 5936 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 6384 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 6496 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_107
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_115
timestamp 1698431365
transform 1 0 7112 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1698431365
transform 1 0 1120 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_12
timestamp 1698431365
transform 1 0 1344 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_20
timestamp 1698431365
transform 1 0 1792 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_64
timestamp 1698431365
transform 1 0 4256 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 4480 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_82
timestamp 1698431365
transform 1 0 5264 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_16
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_24
timestamp 1698431365
transform 1 0 2016 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_28
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_39
timestamp 1698431365
transform 1 0 2856 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_94
timestamp 1698431365
transform 1 0 5936 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_102
timestamp 1698431365
transform 1 0 6384 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_109
timestamp 1698431365
transform 1 0 6776 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_10
timestamp 1698431365
transform 1 0 1232 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_14
timestamp 1698431365
transform 1 0 1456 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_65
timestamp 1698431365
transform 1 0 4312 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 4536 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_72
timestamp 1698431365
transform 1 0 4704 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_80
timestamp 1698431365
transform 1 0 5152 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_97
timestamp 1698431365
transform 1 0 6104 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_101
timestamp 1698431365
transform 1 0 6328 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_18
timestamp 1698431365
transform 1 0 1680 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_26
timestamp 1698431365
transform 1 0 2128 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_30
timestamp 1698431365
transform 1 0 2352 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_32
timestamp 1698431365
transform 1 0 2464 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_100
timestamp 1698431365
transform 1 0 6272 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_102
timestamp 1698431365
transform 1 0 6384 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_107
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 1120 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_12
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_28
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_30
timestamp 1698431365
transform 1 0 2352 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_65
timestamp 1698431365
transform 1 0 4312 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 4536 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_72
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_80
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_82
timestamp 1698431365
transform 1 0 5264 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_99
timestamp 1698431365
transform 1 0 6216 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_101
timestamp 1698431365
transform 1 0 6328 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_45
timestamp 1698431365
transform 1 0 3192 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_47
timestamp 1698431365
transform 1 0 3304 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_54
timestamp 1698431365
transform 1 0 3696 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_115
timestamp 1698431365
transform 1 0 7112 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 2576 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_50
timestamp 1698431365
transform 1 0 3472 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_58
timestamp 1698431365
transform 1 0 3920 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_62
timestamp 1698431365
transform 1 0 4144 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_88
timestamp 1698431365
transform 1 0 5600 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_104
timestamp 1698431365
transform 1 0 6496 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_112
timestamp 1698431365
transform 1 0 6944 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_45
timestamp 1698431365
transform 1 0 3192 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_83
timestamp 1698431365
transform 1 0 5320 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_99
timestamp 1698431365
transform 1 0 6216 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 6440 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_115
timestamp 1698431365
transform 1 0 7112 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_36
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_70
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_104
timestamp 1698431365
transform 1 0 6496 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_112
timestamp 1698431365
transform 1 0 6944 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5600 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 6104 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 6216 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7168 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 7168 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 3752 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 3080 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6384 0 -1 4704
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1698431365
transform 1 0 6384 0 -1 3920
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output9
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output10
timestamp 1698431365
transform -1 0 1568 0 1 3136
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output11
timestamp 1698431365
transform 1 0 3416 0 1 1568
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 7280 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_13
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 7280 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_14
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 7280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_15
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 7280 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_16
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_17
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 7280 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_18
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 7280 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_19
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 7280 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_20
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 7280 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_21
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 7280 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_22
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 7280 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_23
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 7280 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_25
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_26
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_27
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_28
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_29
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_30
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_31
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_32
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_33
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_34
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_35
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_36
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_37
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_38
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_39
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_40
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_41
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_42
timestamp 1698431365
transform 1 0 2576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_43
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_44
timestamp 1698431365
transform 1 0 6384 0 -1 6272
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 4368 400 4424 0 FreeSans 224 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 7600 4704 8000 4760 0 FreeSans 224 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 7600 3696 8000 3752 0 FreeSans 224 0 0 0 gfpga_pad_GPIO_PAD[0]
port 2 nsew signal bidirectional
flabel metal2 s 4368 0 4424 400 0 FreeSans 224 90 0 0 gfpga_pad_GPIO_PAD[1]
port 3 nsew signal bidirectional
flabel metal3 s 0 3696 400 3752 0 FreeSans 224 0 0 0 gfpga_pad_GPIO_PAD[2]
port 4 nsew signal bidirectional
flabel metal2 s 2688 0 2744 400 0 FreeSans 224 90 0 0 gfpga_pad_GPIO_PAD[3]
port 5 nsew signal bidirectional
flabel metal3 s 7600 4368 8000 4424 0 FreeSans 224 0 0 0 pReset
port 6 nsew signal input
flabel metal3 s 0 4704 400 4760 0 FreeSans 224 0 0 0 prog_clk
port 7 nsew signal input
flabel metal3 s 7600 3360 8000 3416 0 FreeSans 224 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 8 nsew signal tristate
flabel metal3 s 7600 3024 8000 3080 0 FreeSans 224 0 0 0 right_width_0_height_0_subtile_0__pin_outpad_0_
port 9 nsew signal input
flabel metal2 s 4032 0 4088 400 0 FreeSans 224 90 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 10 nsew signal tristate
flabel metal2 s 3696 0 3752 400 0 FreeSans 224 90 0 0 right_width_0_height_0_subtile_1__pin_outpad_0_
port 11 nsew signal input
flabel metal3 s 0 3360 400 3416 0 FreeSans 224 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 12 nsew signal tristate
flabel metal3 s 0 3024 400 3080 0 FreeSans 224 0 0 0 right_width_0_height_0_subtile_2__pin_outpad_0_
port 13 nsew signal input
flabel metal2 s 3360 0 3416 400 0 FreeSans 224 90 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 14 nsew signal tristate
flabel metal2 s 3024 0 3080 400 0 FreeSans 224 90 0 0 right_width_0_height_0_subtile_3__pin_outpad_0_
port 15 nsew signal input
flabel metal4 s 1418 1538 1578 6302 0 FreeSans 640 90 0 0 vdd
port 16 nsew power bidirectional
flabel metal4 s 3070 1538 3230 6302 0 FreeSans 640 90 0 0 vdd
port 16 nsew power bidirectional
flabel metal4 s 4722 1538 4882 6302 0 FreeSans 640 90 0 0 vdd
port 16 nsew power bidirectional
flabel metal4 s 6374 1538 6534 6302 0 FreeSans 640 90 0 0 vdd
port 16 nsew power bidirectional
flabel metal4 s 2244 1538 2404 6302 0 FreeSans 640 90 0 0 vss
port 17 nsew ground bidirectional
flabel metal4 s 3896 1538 4056 6302 0 FreeSans 640 90 0 0 vss
port 17 nsew ground bidirectional
flabel metal4 s 5548 1538 5708 6302 0 FreeSans 640 90 0 0 vss
port 17 nsew ground bidirectional
flabel metal4 s 7200 1538 7360 6302 0 FreeSans 640 90 0 0 vss
port 17 nsew ground bidirectional
rlabel metal1 3976 5880 3976 5880 0 vdd
rlabel via1 4016 6272 4016 6272 0 vss
rlabel metal2 3500 3920 3500 3920 0 _00_
rlabel metal3 3388 4564 3388 4564 0 _01_
rlabel metal2 4508 5460 4508 5460 0 _02_
rlabel metal2 5628 3416 5628 3416 0 _03_
rlabel metal2 868 4452 868 4452 0 ccff_head
rlabel metal2 7028 4592 7028 4592 0 ccff_tail
rlabel metal2 4172 4480 4172 4480 0 clknet_0_prog_clk
rlabel metal2 2156 3360 2156 3360 0 clknet_1_0__leaf_prog_clk
rlabel metal2 3556 5320 3556 5320 0 clknet_1_1__leaf_prog_clk
rlabel metal2 5180 3360 5180 3360 0 gfpga_pad_GPIO_PAD[0]
rlabel metal2 3612 2576 3612 2576 0 gfpga_pad_GPIO_PAD[1]
rlabel metal2 3052 2632 3052 2632 0 gfpga_pad_GPIO_PAD[2]
rlabel metal2 2716 427 2716 427 0 gfpga_pad_GPIO_PAD[3]
rlabel metal2 5964 3304 5964 3304 0 logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 4284 4984 4284 4984 0 logical_tile_io_mode_io__1.ccff_tail
rlabel metal3 5628 4564 5628 4564 0 logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 2212 3276 2212 3276 0 net1
rlabel metal2 2380 3332 2380 3332 0 net10
rlabel metal2 3556 2100 3556 2100 0 net11
rlabel metal2 3780 5460 3780 5460 0 net12
rlabel metal2 2772 4368 2772 4368 0 net13
rlabel metal3 4900 3780 4900 3780 0 net14
rlabel metal3 3248 4900 3248 4900 0 net2
rlabel metal2 4844 3080 4844 3080 0 net3
rlabel metal2 4088 2940 4088 2940 0 net4
rlabel metal2 2492 3304 2492 3304 0 net5
rlabel metal2 3388 2884 3388 2884 0 net6
rlabel metal2 5908 3766 5908 3766 0 net7
rlabel metal2 4984 2436 4984 2436 0 net8
rlabel metal2 4172 2380 4172 2380 0 net9
rlabel metal2 7084 4144 7084 4144 0 pReset
rlabel metal3 2912 4116 2912 4116 0 prog_clk
rlabel metal2 7028 3528 7028 3528 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 7385 3052 7385 3052 0 right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 4060 483 4060 483 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 3836 1792 3836 1792 0 right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal3 735 3388 735 3388 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 868 3024 868 3024 0 right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 3388 1099 3388 1099 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 3052 1043 3052 1043 0 right_width_0_height_0_subtile_3__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 8000 8000
<< end >>
