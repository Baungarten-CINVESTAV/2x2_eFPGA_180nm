magic
tech gf180mcuD
magscale 1 5
timestamp 1702149426
<< obsm1 >>
rect 672 463 23296 22609
<< metal2 >>
rect 3696 23600 3752 24000
rect 4032 23600 4088 24000
rect 6720 23600 6776 24000
rect 7056 23600 7112 24000
rect 7392 23600 7448 24000
rect 8400 23600 8456 24000
rect 8736 23600 8792 24000
rect 9072 23600 9128 24000
rect 9408 23600 9464 24000
rect 9744 23600 9800 24000
rect 10080 23600 10136 24000
rect 10416 23600 10472 24000
rect 10752 23600 10808 24000
rect 11088 23600 11144 24000
rect 11424 23600 11480 24000
rect 11760 23600 11816 24000
rect 12096 23600 12152 24000
rect 12432 23600 12488 24000
rect 12768 23600 12824 24000
rect 13104 23600 13160 24000
rect 13440 23600 13496 24000
rect 13776 23600 13832 24000
rect 14112 23600 14168 24000
rect 14448 23600 14504 24000
rect 14784 23600 14840 24000
rect 15120 23600 15176 24000
rect 15456 23600 15512 24000
rect 15792 23600 15848 24000
rect 16128 23600 16184 24000
rect 17136 23600 17192 24000
rect 17472 23600 17528 24000
rect 17808 23600 17864 24000
rect 18144 23600 18200 24000
rect 18480 23600 18536 24000
rect 18816 23600 18872 24000
rect 19152 23600 19208 24000
rect 19488 23600 19544 24000
rect 19824 23600 19880 24000
rect 20160 23600 20216 24000
rect 20496 23600 20552 24000
rect 20832 23600 20888 24000
rect 21168 23600 21224 24000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
rect 13104 0 13160 400
rect 13440 0 13496 400
rect 13776 0 13832 400
rect 14112 0 14168 400
rect 14448 0 14504 400
rect 14784 0 14840 400
rect 15120 0 15176 400
rect 15456 0 15512 400
rect 15792 0 15848 400
rect 16128 0 16184 400
rect 16464 0 16520 400
rect 16800 0 16856 400
rect 17136 0 17192 400
rect 17472 0 17528 400
rect 17808 0 17864 400
rect 18144 0 18200 400
rect 18480 0 18536 400
rect 18816 0 18872 400
rect 19152 0 19208 400
rect 19488 0 19544 400
rect 19824 0 19880 400
rect 20160 0 20216 400
rect 20496 0 20552 400
rect 20832 0 20888 400
rect 21168 0 21224 400
rect 21504 0 21560 400
rect 21840 0 21896 400
rect 22176 0 22232 400
rect 22512 0 22568 400
rect 22848 0 22904 400
rect 23184 0 23240 400
rect 23520 0 23576 400
rect 23856 0 23912 400
<< obsm2 >>
rect 742 23570 3666 23600
rect 3782 23570 4002 23600
rect 4118 23570 6690 23600
rect 6806 23570 7026 23600
rect 7142 23570 7362 23600
rect 7478 23570 8370 23600
rect 8486 23570 8706 23600
rect 8822 23570 9042 23600
rect 9158 23570 9378 23600
rect 9494 23570 9714 23600
rect 9830 23570 10050 23600
rect 10166 23570 10386 23600
rect 10502 23570 10722 23600
rect 10838 23570 11058 23600
rect 11174 23570 11394 23600
rect 11510 23570 11730 23600
rect 11846 23570 12066 23600
rect 12182 23570 12402 23600
rect 12518 23570 12738 23600
rect 12854 23570 13074 23600
rect 13190 23570 13410 23600
rect 13526 23570 13746 23600
rect 13862 23570 14082 23600
rect 14198 23570 14418 23600
rect 14534 23570 14754 23600
rect 14870 23570 15090 23600
rect 15206 23570 15426 23600
rect 15542 23570 15762 23600
rect 15878 23570 16098 23600
rect 16214 23570 17106 23600
rect 17222 23570 17442 23600
rect 17558 23570 17778 23600
rect 17894 23570 18114 23600
rect 18230 23570 18450 23600
rect 18566 23570 18786 23600
rect 18902 23570 19122 23600
rect 19238 23570 19458 23600
rect 19574 23570 19794 23600
rect 19910 23570 20130 23600
rect 20246 23570 20466 23600
rect 20582 23570 20802 23600
rect 20918 23570 21138 23600
rect 21254 23570 23338 23600
rect 742 430 23338 23570
rect 758 9 978 430
rect 1094 9 1314 430
rect 1430 9 1650 430
rect 1766 9 1986 430
rect 2102 9 2322 430
rect 2438 9 2658 430
rect 2774 9 2994 430
rect 3110 9 3330 430
rect 3446 9 3666 430
rect 3782 9 4002 430
rect 4118 9 4338 430
rect 4454 9 4674 430
rect 4790 9 5010 430
rect 5126 9 5346 430
rect 5462 9 5682 430
rect 5798 9 6018 430
rect 6134 9 6354 430
rect 6470 9 6690 430
rect 6806 9 7026 430
rect 7142 9 7362 430
rect 7478 9 7698 430
rect 7814 9 8034 430
rect 8150 9 8370 430
rect 8486 9 8706 430
rect 8822 9 9042 430
rect 9158 9 9378 430
rect 9494 9 9714 430
rect 9830 9 10050 430
rect 10166 9 10386 430
rect 10502 9 10722 430
rect 10838 9 11058 430
rect 11174 9 11394 430
rect 11510 9 11730 430
rect 11846 9 12066 430
rect 12182 9 12402 430
rect 12518 9 12738 430
rect 12854 9 13074 430
rect 13190 9 13410 430
rect 13526 9 13746 430
rect 13862 9 14082 430
rect 14198 9 14418 430
rect 14534 9 14754 430
rect 14870 9 15090 430
rect 15206 9 15426 430
rect 15542 9 15762 430
rect 15878 9 16098 430
rect 16214 9 16434 430
rect 16550 9 16770 430
rect 16886 9 17106 430
rect 17222 9 17442 430
rect 17558 9 17778 430
rect 17894 9 18114 430
rect 18230 9 18450 430
rect 18566 9 18786 430
rect 18902 9 19122 430
rect 19238 9 19458 430
rect 19574 9 19794 430
rect 19910 9 20130 430
rect 20246 9 20466 430
rect 20582 9 20802 430
rect 20918 9 21138 430
rect 21254 9 21474 430
rect 21590 9 21810 430
rect 21926 9 22146 430
rect 22262 9 22482 430
rect 22598 9 22818 430
rect 22934 9 23154 430
rect 23270 9 23338 430
<< metal3 >>
rect 23600 22176 24000 22232
rect 23600 21840 24000 21896
rect 23600 21504 24000 21560
rect 0 21168 400 21224
rect 23600 21168 24000 21224
rect 23600 20832 24000 20888
rect 23600 20496 24000 20552
rect 23600 16128 24000 16184
rect 0 15792 400 15848
rect 23600 15792 24000 15848
rect 23600 15456 24000 15512
rect 23600 15120 24000 15176
rect 23600 14784 24000 14840
rect 23600 14448 24000 14504
rect 23600 14112 24000 14168
rect 23600 13776 24000 13832
rect 23600 13440 24000 13496
rect 23600 13104 24000 13160
rect 23600 12768 24000 12824
rect 23600 12432 24000 12488
rect 23600 12096 24000 12152
rect 23600 11760 24000 11816
rect 23600 11424 24000 11480
rect 23600 11088 24000 11144
rect 23600 10752 24000 10808
rect 23600 10416 24000 10472
rect 23600 10080 24000 10136
rect 23600 9744 24000 9800
rect 23600 9408 24000 9464
rect 23600 9072 24000 9128
rect 0 8736 400 8792
rect 23600 8736 24000 8792
rect 23600 8400 24000 8456
rect 23600 8064 24000 8120
rect 23600 7728 24000 7784
rect 23600 7392 24000 7448
rect 23600 7056 24000 7112
rect 23600 6720 24000 6776
rect 23600 6384 24000 6440
rect 23600 6048 24000 6104
rect 23600 5712 24000 5768
rect 23600 5376 24000 5432
rect 23600 5040 24000 5096
rect 23600 4704 24000 4760
rect 23600 4368 24000 4424
rect 23600 4032 24000 4088
rect 0 3696 400 3752
rect 23600 3696 24000 3752
rect 0 3360 400 3416
rect 23600 3360 24000 3416
rect 0 3024 400 3080
rect 23600 3024 24000 3080
rect 0 2688 400 2744
rect 23600 2688 24000 2744
rect 0 2352 400 2408
rect 23600 2352 24000 2408
rect 0 2016 400 2072
rect 23600 2016 24000 2072
rect 0 1680 400 1736
rect 23600 1680 24000 1736
rect 0 1344 400 1400
rect 23600 1344 24000 1400
rect 23600 1008 24000 1064
rect 23600 672 24000 728
rect 23600 336 24000 392
rect 23600 0 24000 56
<< obsm3 >>
rect 400 22262 23600 22666
rect 400 22146 23570 22262
rect 400 21926 23600 22146
rect 400 21810 23570 21926
rect 400 21590 23600 21810
rect 400 21474 23570 21590
rect 400 21254 23600 21474
rect 430 21138 23570 21254
rect 400 20918 23600 21138
rect 400 20802 23570 20918
rect 400 20582 23600 20802
rect 400 20466 23570 20582
rect 400 16214 23600 20466
rect 400 16098 23570 16214
rect 400 15878 23600 16098
rect 430 15762 23570 15878
rect 400 15542 23600 15762
rect 400 15426 23570 15542
rect 400 15206 23600 15426
rect 400 15090 23570 15206
rect 400 14870 23600 15090
rect 400 14754 23570 14870
rect 400 14534 23600 14754
rect 400 14418 23570 14534
rect 400 14198 23600 14418
rect 400 14082 23570 14198
rect 400 13862 23600 14082
rect 400 13746 23570 13862
rect 400 13526 23600 13746
rect 400 13410 23570 13526
rect 400 13190 23600 13410
rect 400 13074 23570 13190
rect 400 12854 23600 13074
rect 400 12738 23570 12854
rect 400 12518 23600 12738
rect 400 12402 23570 12518
rect 400 12182 23600 12402
rect 400 12066 23570 12182
rect 400 11846 23600 12066
rect 400 11730 23570 11846
rect 400 11510 23600 11730
rect 400 11394 23570 11510
rect 400 11174 23600 11394
rect 400 11058 23570 11174
rect 400 10838 23600 11058
rect 400 10722 23570 10838
rect 400 10502 23600 10722
rect 400 10386 23570 10502
rect 400 10166 23600 10386
rect 400 10050 23570 10166
rect 400 9830 23600 10050
rect 400 9714 23570 9830
rect 400 9494 23600 9714
rect 400 9378 23570 9494
rect 400 9158 23600 9378
rect 400 9042 23570 9158
rect 400 8822 23600 9042
rect 430 8706 23570 8822
rect 400 8486 23600 8706
rect 400 8370 23570 8486
rect 400 8150 23600 8370
rect 400 8034 23570 8150
rect 400 7814 23600 8034
rect 400 7698 23570 7814
rect 400 7478 23600 7698
rect 400 7362 23570 7478
rect 400 7142 23600 7362
rect 400 7026 23570 7142
rect 400 6806 23600 7026
rect 400 6690 23570 6806
rect 400 6470 23600 6690
rect 400 6354 23570 6470
rect 400 6134 23600 6354
rect 400 6018 23570 6134
rect 400 5798 23600 6018
rect 400 5682 23570 5798
rect 400 5462 23600 5682
rect 400 5346 23570 5462
rect 400 5126 23600 5346
rect 400 5010 23570 5126
rect 400 4790 23600 5010
rect 400 4674 23570 4790
rect 400 4454 23600 4674
rect 400 4338 23570 4454
rect 400 4118 23600 4338
rect 400 4002 23570 4118
rect 400 3782 23600 4002
rect 430 3666 23570 3782
rect 400 3446 23600 3666
rect 430 3330 23570 3446
rect 400 3110 23600 3330
rect 430 2994 23570 3110
rect 400 2774 23600 2994
rect 430 2658 23570 2774
rect 400 2438 23600 2658
rect 430 2322 23570 2438
rect 400 2102 23600 2322
rect 430 1986 23570 2102
rect 400 1766 23600 1986
rect 430 1650 23570 1766
rect 400 1430 23600 1650
rect 430 1314 23570 1430
rect 400 1094 23600 1314
rect 400 978 23570 1094
rect 400 758 23600 978
rect 400 642 23570 758
rect 400 422 23600 642
rect 400 306 23570 422
rect 400 86 23600 306
rect 400 14 23570 86
<< metal4 >>
rect 2224 1538 2384 22374
rect 9904 1538 10064 22374
rect 17584 1538 17744 22374
<< obsm4 >>
rect 18326 4433 22386 10911
<< labels >>
rlabel metal2 s 23520 0 23576 400 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 2 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 3 nsew signal input
rlabel metal2 s 336 0 392 400 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 4 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 ccff_head
port 5 nsew signal input
rlabel metal3 s 23600 13104 24000 13160 6 ccff_tail
port 6 nsew signal output
rlabel metal2 s 20832 0 20888 400 6 chanx_left_in[0]
port 7 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 chanx_left_in[10]
port 8 nsew signal input
rlabel metal2 s 0 0 56 400 6 chanx_left_in[11]
port 9 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 chanx_left_in[12]
port 10 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 chanx_left_in[13]
port 11 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 chanx_left_in[14]
port 12 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 chanx_left_in[15]
port 13 nsew signal input
rlabel metal2 s 12096 23600 12152 24000 6 chanx_left_in[16]
port 14 nsew signal input
rlabel metal2 s 6720 23600 6776 24000 6 chanx_left_in[17]
port 15 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 chanx_left_in[18]
port 16 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 chanx_left_in[19]
port 17 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 chanx_left_in[1]
port 18 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 chanx_left_in[2]
port 19 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 chanx_left_in[3]
port 20 nsew signal input
rlabel metal2 s 13440 23600 13496 24000 6 chanx_left_in[4]
port 21 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 chanx_left_in[5]
port 22 nsew signal input
rlabel metal2 s 16128 23600 16184 24000 6 chanx_left_in[6]
port 23 nsew signal input
rlabel metal2 s 672 0 728 400 6 chanx_left_in[7]
port 24 nsew signal input
rlabel metal2 s 15120 23600 15176 24000 6 chanx_left_in[8]
port 25 nsew signal input
rlabel metal2 s 11424 23600 11480 24000 6 chanx_left_in[9]
port 26 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 chanx_left_out[0]
port 27 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 chanx_left_out[10]
port 28 nsew signal output
rlabel metal2 s 8400 23600 8456 24000 6 chanx_left_out[11]
port 29 nsew signal output
rlabel metal2 s 9072 0 9128 400 6 chanx_left_out[12]
port 30 nsew signal output
rlabel metal2 s 3696 0 3752 400 6 chanx_left_out[13]
port 31 nsew signal output
rlabel metal3 s 23600 22176 24000 22232 6 chanx_left_out[14]
port 32 nsew signal output
rlabel metal2 s 20496 0 20552 400 6 chanx_left_out[15]
port 33 nsew signal output
rlabel metal2 s 7392 23600 7448 24000 6 chanx_left_out[16]
port 34 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 chanx_left_out[17]
port 35 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 chanx_left_out[18]
port 36 nsew signal output
rlabel metal2 s 10752 0 10808 400 6 chanx_left_out[19]
port 37 nsew signal output
rlabel metal3 s 23600 21504 24000 21560 6 chanx_left_out[1]
port 38 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 chanx_left_out[2]
port 39 nsew signal output
rlabel metal2 s 14784 0 14840 400 6 chanx_left_out[3]
port 40 nsew signal output
rlabel metal3 s 23600 1344 24000 1400 6 chanx_left_out[4]
port 41 nsew signal output
rlabel metal2 s 10080 23600 10136 24000 6 chanx_left_out[5]
port 42 nsew signal output
rlabel metal2 s 18144 0 18200 400 6 chanx_left_out[6]
port 43 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 chanx_left_out[7]
port 44 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 chanx_left_out[8]
port 45 nsew signal output
rlabel metal2 s 13104 23600 13160 24000 6 chanx_left_out[9]
port 46 nsew signal output
rlabel metal3 s 23600 20496 24000 20552 6 chanx_right_in[0]
port 47 nsew signal input
rlabel metal2 s 9408 23600 9464 24000 6 chanx_right_in[10]
port 48 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 chanx_right_in[11]
port 49 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 chanx_right_in[12]
port 50 nsew signal input
rlabel metal3 s 23600 21840 24000 21896 6 chanx_right_in[13]
port 51 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 chanx_right_in[14]
port 52 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 chanx_right_in[15]
port 53 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 chanx_right_in[16]
port 54 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 chanx_right_in[17]
port 55 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 chanx_right_in[18]
port 56 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 chanx_right_in[19]
port 57 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 chanx_right_in[1]
port 58 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 chanx_right_in[2]
port 59 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 chanx_right_in[3]
port 60 nsew signal input
rlabel metal2 s 10416 23600 10472 24000 6 chanx_right_in[4]
port 61 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 chanx_right_in[5]
port 62 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 chanx_right_in[6]
port 63 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 chanx_right_in[7]
port 64 nsew signal input
rlabel metal2 s 12768 23600 12824 24000 6 chanx_right_in[8]
port 65 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 chanx_right_in[9]
port 66 nsew signal input
rlabel metal3 s 23600 21168 24000 21224 6 chanx_right_out[0]
port 67 nsew signal output
rlabel metal2 s 11760 23600 11816 24000 6 chanx_right_out[10]
port 68 nsew signal output
rlabel metal2 s 14112 0 14168 400 6 chanx_right_out[11]
port 69 nsew signal output
rlabel metal2 s 14448 23600 14504 24000 6 chanx_right_out[12]
port 70 nsew signal output
rlabel metal2 s 6048 0 6104 400 6 chanx_right_out[13]
port 71 nsew signal output
rlabel metal2 s 7392 0 7448 400 6 chanx_right_out[14]
port 72 nsew signal output
rlabel metal2 s 8736 0 8792 400 6 chanx_right_out[15]
port 73 nsew signal output
rlabel metal3 s 23600 2016 24000 2072 6 chanx_right_out[16]
port 74 nsew signal output
rlabel metal2 s 12432 23600 12488 24000 6 chanx_right_out[17]
port 75 nsew signal output
rlabel metal2 s 7056 23600 7112 24000 6 chanx_right_out[18]
port 76 nsew signal output
rlabel metal2 s 4368 0 4424 400 6 chanx_right_out[19]
port 77 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 chanx_right_out[1]
port 78 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 chanx_right_out[2]
port 79 nsew signal output
rlabel metal2 s 7728 0 7784 400 6 chanx_right_out[3]
port 80 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 chanx_right_out[4]
port 81 nsew signal output
rlabel metal2 s 14784 23600 14840 24000 6 chanx_right_out[5]
port 82 nsew signal output
rlabel metal2 s 4032 0 4088 400 6 chanx_right_out[6]
port 83 nsew signal output
rlabel metal2 s 13776 23600 13832 24000 6 chanx_right_out[7]
port 84 nsew signal output
rlabel metal3 s 0 1344 400 1400 6 chanx_right_out[8]
port 85 nsew signal output
rlabel metal2 s 15456 23600 15512 24000 6 chanx_right_out[9]
port 86 nsew signal output
rlabel metal2 s 17136 23600 17192 24000 6 chany_bottom_in[0]
port 87 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 chany_bottom_in[10]
port 88 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 chany_bottom_in[11]
port 89 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 chany_bottom_in[12]
port 90 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 chany_bottom_in[13]
port 91 nsew signal input
rlabel metal2 s 17472 23600 17528 24000 6 chany_bottom_in[14]
port 92 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 chany_bottom_in[15]
port 93 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 chany_bottom_in[16]
port 94 nsew signal input
rlabel metal3 s 23600 9744 24000 9800 6 chany_bottom_in[17]
port 95 nsew signal input
rlabel metal3 s 23600 5376 24000 5432 6 chany_bottom_in[18]
port 96 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 chany_bottom_in[19]
port 97 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 chany_bottom_in[1]
port 98 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 chany_bottom_in[2]
port 99 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 chany_bottom_in[3]
port 100 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 chany_bottom_in[4]
port 101 nsew signal input
rlabel metal3 s 23600 2688 24000 2744 6 chany_bottom_in[5]
port 102 nsew signal input
rlabel metal2 s 20832 23600 20888 24000 6 chany_bottom_in[6]
port 103 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 chany_bottom_in[7]
port 104 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 chany_bottom_in[8]
port 105 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 chany_bottom_in[9]
port 106 nsew signal input
rlabel metal2 s 17472 0 17528 400 6 chany_bottom_out[0]
port 107 nsew signal output
rlabel metal2 s 6384 0 6440 400 6 chany_bottom_out[10]
port 108 nsew signal output
rlabel metal2 s 19488 23600 19544 24000 6 chany_bottom_out[11]
port 109 nsew signal output
rlabel metal3 s 23600 2352 24000 2408 6 chany_bottom_out[12]
port 110 nsew signal output
rlabel metal2 s 14112 23600 14168 24000 6 chany_bottom_out[13]
port 111 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 chany_bottom_out[14]
port 112 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 chany_bottom_out[15]
port 113 nsew signal output
rlabel metal3 s 23600 672 24000 728 6 chany_bottom_out[16]
port 114 nsew signal output
rlabel metal3 s 23600 7056 24000 7112 6 chany_bottom_out[17]
port 115 nsew signal output
rlabel metal3 s 23600 7728 24000 7784 6 chany_bottom_out[18]
port 116 nsew signal output
rlabel metal2 s 9744 23600 9800 24000 6 chany_bottom_out[19]
port 117 nsew signal output
rlabel metal2 s 4032 23600 4088 24000 6 chany_bottom_out[1]
port 118 nsew signal output
rlabel metal2 s 11088 23600 11144 24000 6 chany_bottom_out[2]
port 119 nsew signal output
rlabel metal3 s 23600 9072 24000 9128 6 chany_bottom_out[3]
port 120 nsew signal output
rlabel metal3 s 23600 336 24000 392 6 chany_bottom_out[4]
port 121 nsew signal output
rlabel metal3 s 23600 6720 24000 6776 6 chany_bottom_out[5]
port 122 nsew signal output
rlabel metal2 s 21168 23600 21224 24000 6 chany_bottom_out[6]
port 123 nsew signal output
rlabel metal3 s 0 2688 400 2744 6 chany_bottom_out[7]
port 124 nsew signal output
rlabel metal3 s 23600 20832 24000 20888 6 chany_bottom_out[8]
port 125 nsew signal output
rlabel metal2 s 20160 23600 20216 24000 6 chany_bottom_out[9]
port 126 nsew signal output
rlabel metal2 s 3696 23600 3752 24000 6 chany_top_in[0]
port 127 nsew signal input
rlabel metal2 s 19152 23600 19208 24000 6 chany_top_in[10]
port 128 nsew signal input
rlabel metal3 s 23600 12096 24000 12152 6 chany_top_in[11]
port 129 nsew signal input
rlabel metal2 s 15792 23600 15848 24000 6 chany_top_in[12]
port 130 nsew signal input
rlabel metal3 s 23600 4704 24000 4760 6 chany_top_in[13]
port 131 nsew signal input
rlabel metal3 s 0 2352 400 2408 6 chany_top_in[14]
port 132 nsew signal input
rlabel metal3 s 23600 16128 24000 16184 6 chany_top_in[15]
port 133 nsew signal input
rlabel metal3 s 23600 6384 24000 6440 6 chany_top_in[16]
port 134 nsew signal input
rlabel metal3 s 23600 3024 24000 3080 6 chany_top_in[17]
port 135 nsew signal input
rlabel metal2 s 9072 23600 9128 24000 6 chany_top_in[18]
port 136 nsew signal input
rlabel metal3 s 23600 12768 24000 12824 6 chany_top_in[19]
port 137 nsew signal input
rlabel metal2 s 10752 23600 10808 24000 6 chany_top_in[1]
port 138 nsew signal input
rlabel metal3 s 23600 5040 24000 5096 6 chany_top_in[2]
port 139 nsew signal input
rlabel metal3 s 23600 11424 24000 11480 6 chany_top_in[3]
port 140 nsew signal input
rlabel metal3 s 23600 4368 24000 4424 6 chany_top_in[4]
port 141 nsew signal input
rlabel metal2 s 18480 23600 18536 24000 6 chany_top_in[5]
port 142 nsew signal input
rlabel metal3 s 0 1680 400 1736 6 chany_top_in[6]
port 143 nsew signal input
rlabel metal3 s 23600 14112 24000 14168 6 chany_top_in[7]
port 144 nsew signal input
rlabel metal2 s 19824 23600 19880 24000 6 chany_top_in[8]
port 145 nsew signal input
rlabel metal3 s 0 2016 400 2072 6 chany_top_in[9]
port 146 nsew signal input
rlabel metal2 s 8736 23600 8792 24000 6 chany_top_out[0]
port 147 nsew signal output
rlabel metal3 s 23600 3696 24000 3752 6 chany_top_out[10]
port 148 nsew signal output
rlabel metal3 s 0 3024 400 3080 6 chany_top_out[11]
port 149 nsew signal output
rlabel metal3 s 23600 1680 24000 1736 6 chany_top_out[12]
port 150 nsew signal output
rlabel metal3 s 0 3360 400 3416 6 chany_top_out[13]
port 151 nsew signal output
rlabel metal3 s 23600 6048 24000 6104 6 chany_top_out[14]
port 152 nsew signal output
rlabel metal2 s 18144 23600 18200 24000 6 chany_top_out[15]
port 153 nsew signal output
rlabel metal3 s 23600 0 24000 56 6 chany_top_out[16]
port 154 nsew signal output
rlabel metal3 s 23600 3360 24000 3416 6 chany_top_out[17]
port 155 nsew signal output
rlabel metal3 s 23600 8736 24000 8792 6 chany_top_out[18]
port 156 nsew signal output
rlabel metal3 s 23600 8064 24000 8120 6 chany_top_out[19]
port 157 nsew signal output
rlabel metal2 s 18816 23600 18872 24000 6 chany_top_out[1]
port 158 nsew signal output
rlabel metal3 s 23600 7392 24000 7448 6 chany_top_out[2]
port 159 nsew signal output
rlabel metal3 s 23600 4032 24000 4088 6 chany_top_out[3]
port 160 nsew signal output
rlabel metal3 s 23600 1008 24000 1064 6 chany_top_out[4]
port 161 nsew signal output
rlabel metal3 s 23600 5712 24000 5768 6 chany_top_out[5]
port 162 nsew signal output
rlabel metal3 s 23600 8400 24000 8456 6 chany_top_out[6]
port 163 nsew signal output
rlabel metal2 s 20496 23600 20552 24000 6 chany_top_out[7]
port 164 nsew signal output
rlabel metal2 s 17808 23600 17864 24000 6 chany_top_out[8]
port 165 nsew signal output
rlabel metal3 s 23600 9408 24000 9464 6 chany_top_out[9]
port 166 nsew signal output
rlabel metal3 s 23600 10752 24000 10808 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 167 nsew signal input
rlabel metal3 s 23600 15456 24000 15512 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 168 nsew signal input
rlabel metal3 s 23600 15120 24000 15176 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 169 nsew signal input
rlabel metal3 s 23600 14448 24000 14504 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 170 nsew signal input
rlabel metal3 s 23600 13440 24000 13496 6 pReset
port 171 nsew signal input
rlabel metal3 s 0 15792 400 15848 6 prog_clk
port 172 nsew signal input
rlabel metal3 s 23600 15792 24000 15848 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 173 nsew signal input
rlabel metal3 s 23600 13776 24000 13832 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 174 nsew signal input
rlabel metal3 s 23600 14784 24000 14840 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 175 nsew signal input
rlabel metal3 s 23600 10416 24000 10472 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 176 nsew signal input
rlabel metal3 s 23600 11088 24000 11144 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 177 nsew signal input
rlabel metal3 s 23600 11760 24000 11816 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 178 nsew signal input
rlabel metal3 s 23600 10080 24000 10136 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 179 nsew signal input
rlabel metal3 s 23600 12432 24000 12488 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 180 nsew signal input
rlabel metal4 s 2224 1538 2384 22374 6 vdd
port 181 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 22374 6 vdd
port 181 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 22374 6 vss
port 182 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1114600
string GDS_FILE /home/baungarten/Desktop/2x2_FPGA_180nmD/openlane/sb_1__1_/runs/23_12_09_13_16/results/signoff/sb_1__1_.magic.gds
string GDS_START 126026
<< end >>

