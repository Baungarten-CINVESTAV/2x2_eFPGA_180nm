// This is the unpowered netlist.
module sb_1__0_ (ccff_head,
    ccff_tail,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
    right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
    right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
    right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out,
    chany_top_in,
    chany_top_out);
 input ccff_head;
 output ccff_tail;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input [19:0] chanx_left_in;
 output [19:0] chanx_left_out;
 input [19:0] chanx_right_in;
 output [19:0] chanx_right_out;
 input [19:0] chany_top_in;
 output [19:0] chany_top_out;

 wire net96;
 wire net93;
 wire net92;
 wire net95;
 wire net94;
 wire net91;
 wire net88;
 wire net87;
 wire net90;
 wire net89;
 wire net86;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire clknet_0_prog_clk;
 wire clknet_3_0__leaf_prog_clk;
 wire clknet_3_1__leaf_prog_clk;
 wire clknet_3_2__leaf_prog_clk;
 wire clknet_3_3__leaf_prog_clk;
 wire clknet_3_4__leaf_prog_clk;
 wire clknet_3_5__leaf_prog_clk;
 wire clknet_3_6__leaf_prog_clk;
 wire clknet_3_7__leaf_prog_clk;
 wire \mem_left_track_1.DFFR_0_.D ;
 wire \mem_left_track_1.DFFR_0_.Q ;
 wire \mem_left_track_1.DFFR_1_.Q ;
 wire \mem_left_track_1.DFFR_2_.Q ;
 wire \mem_left_track_1.DFFR_3_.Q ;
 wire \mem_left_track_1.DFFR_4_.Q ;
 wire \mem_left_track_1.DFFR_5_.Q ;
 wire \mem_left_track_1.DFFR_6_.Q ;
 wire \mem_left_track_1.DFFR_7_.Q ;
 wire \mem_left_track_17.DFFR_0_.D ;
 wire \mem_left_track_17.DFFR_0_.Q ;
 wire \mem_left_track_17.DFFR_1_.Q ;
 wire \mem_left_track_17.DFFR_2_.Q ;
 wire \mem_left_track_17.DFFR_3_.Q ;
 wire \mem_left_track_17.DFFR_4_.Q ;
 wire \mem_left_track_17.DFFR_5_.Q ;
 wire \mem_left_track_25.DFFR_0_.Q ;
 wire \mem_left_track_25.DFFR_1_.Q ;
 wire \mem_left_track_25.DFFR_2_.Q ;
 wire \mem_left_track_25.DFFR_3_.Q ;
 wire \mem_left_track_25.DFFR_4_.Q ;
 wire \mem_left_track_25.DFFR_5_.Q ;
 wire \mem_left_track_33.DFFR_0_.Q ;
 wire \mem_left_track_33.DFFR_1_.Q ;
 wire \mem_left_track_33.DFFR_2_.Q ;
 wire \mem_left_track_33.DFFR_3_.Q ;
 wire \mem_left_track_33.DFFR_4_.Q ;
 wire \mem_left_track_9.DFFR_0_.Q ;
 wire \mem_left_track_9.DFFR_1_.Q ;
 wire \mem_left_track_9.DFFR_2_.Q ;
 wire \mem_left_track_9.DFFR_3_.Q ;
 wire \mem_left_track_9.DFFR_4_.Q ;
 wire \mem_right_track_0.DFFR_0_.D ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_0.DFFR_2_.Q ;
 wire \mem_right_track_0.DFFR_3_.Q ;
 wire \mem_right_track_0.DFFR_4_.Q ;
 wire \mem_right_track_0.DFFR_5_.Q ;
 wire \mem_right_track_0.DFFR_6_.Q ;
 wire \mem_right_track_0.DFFR_7_.Q ;
 wire \mem_right_track_16.DFFR_0_.D ;
 wire \mem_right_track_16.DFFR_0_.Q ;
 wire \mem_right_track_16.DFFR_1_.Q ;
 wire \mem_right_track_16.DFFR_2_.Q ;
 wire \mem_right_track_16.DFFR_3_.Q ;
 wire \mem_right_track_16.DFFR_4_.Q ;
 wire \mem_right_track_16.DFFR_5_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_2_.Q ;
 wire \mem_right_track_24.DFFR_3_.Q ;
 wire \mem_right_track_24.DFFR_4_.Q ;
 wire \mem_right_track_24.DFFR_5_.Q ;
 wire \mem_right_track_32.DFFR_0_.Q ;
 wire \mem_right_track_32.DFFR_1_.Q ;
 wire \mem_right_track_32.DFFR_2_.Q ;
 wire \mem_right_track_32.DFFR_3_.Q ;
 wire \mem_right_track_32.DFFR_4_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire \mem_right_track_8.DFFR_1_.Q ;
 wire \mem_right_track_8.DFFR_2_.Q ;
 wire \mem_right_track_8.DFFR_3_.Q ;
 wire \mem_right_track_8.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_0.DFFR_2_.Q ;
 wire \mem_top_track_0.DFFR_3_.Q ;
 wire \mem_top_track_0.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_5_.Q ;
 wire \mem_top_track_10.DFFR_0_.D ;
 wire \mem_top_track_10.DFFR_0_.Q ;
 wire \mem_top_track_10.DFFR_1_.Q ;
 wire \mem_top_track_12.DFFR_0_.Q ;
 wire \mem_top_track_12.DFFR_1_.Q ;
 wire \mem_top_track_14.DFFR_0_.Q ;
 wire \mem_top_track_14.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_18.DFFR_0_.Q ;
 wire \mem_top_track_18.DFFR_1_.Q ;
 wire \mem_top_track_2.DFFR_0_.Q ;
 wire \mem_top_track_2.DFFR_1_.Q ;
 wire \mem_top_track_2.DFFR_2_.Q ;
 wire \mem_top_track_2.DFFR_3_.Q ;
 wire \mem_top_track_2.DFFR_4_.Q ;
 wire \mem_top_track_2.DFFR_5_.Q ;
 wire \mem_top_track_20.DFFR_0_.Q ;
 wire \mem_top_track_20.DFFR_1_.Q ;
 wire \mem_top_track_22.DFFR_0_.Q ;
 wire \mem_top_track_22.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_26.DFFR_0_.Q ;
 wire \mem_top_track_26.DFFR_1_.Q ;
 wire \mem_top_track_28.DFFR_0_.Q ;
 wire \mem_top_track_28.DFFR_1_.Q ;
 wire \mem_top_track_38.DFFR_0_.Q ;
 wire \mem_top_track_4.DFFR_0_.Q ;
 wire \mem_top_track_4.DFFR_1_.Q ;
 wire \mem_top_track_4.DFFR_2_.Q ;
 wire \mem_top_track_4.DFFR_3_.Q ;
 wire \mem_top_track_4.DFFR_4_.Q ;
 wire \mem_top_track_4.DFFR_5_.Q ;
 wire \mem_top_track_6.DFFR_0_.Q ;
 wire \mem_top_track_6.DFFR_1_.Q ;
 wire \mem_top_track_6.DFFR_2_.Q ;
 wire \mem_top_track_6.DFFR_3_.Q ;
 wire \mem_top_track_6.DFFR_4_.Q ;
 wire \mem_top_track_6.DFFR_5_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net8;
 wire net9;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__213__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__CLK (.I(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__CLK (.I(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(chanx_left_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(chanx_left_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(chanx_left_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(chanx_left_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(chanx_left_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(chanx_left_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(chanx_left_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(chanx_left_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(chanx_left_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(chanx_left_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(chanx_right_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(chanx_right_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(chanx_right_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(chanx_right_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(chanx_right_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(chanx_right_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(chanx_right_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(chanx_right_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(chanx_right_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(chanx_right_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(chanx_left_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(chanx_right_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(chanx_right_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(chanx_right_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(chanx_right_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(chanx_right_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(chanx_left_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(chanx_left_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(chanx_left_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(chanx_left_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(chanx_left_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(chanx_left_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(chanx_left_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _125_ (.I(net35),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _126_ (.I(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _127_ (.I(_113_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _128_ (.I(_114_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _129_ (.I(_114_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _130_ (.I(_114_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _131_ (.I(_114_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _132_ (.I(_114_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _133_ (.I(_114_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _134_ (.I(_114_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _135_ (.I(_114_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _136_ (.I(_114_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _137_ (.I(_114_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _138_ (.I(_113_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _139_ (.I(_115_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _140_ (.I(_115_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _141_ (.I(_115_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _142_ (.I(_115_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _143_ (.I(_115_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _144_ (.I(_115_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _145_ (.I(_115_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _146_ (.I(_115_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _147_ (.I(_115_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _148_ (.I(_115_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _149_ (.I(_113_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _150_ (.I(_116_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _151_ (.I(_116_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _152_ (.I(_116_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _153_ (.I(_116_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _154_ (.I(_116_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _155_ (.I(_116_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _156_ (.I(_116_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _157_ (.I(_116_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _158_ (.I(_116_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _159_ (.I(_116_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _160_ (.I(_113_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _161_ (.I(_117_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _162_ (.I(_117_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _163_ (.I(_117_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _164_ (.I(_117_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _165_ (.I(_117_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _166_ (.I(_117_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _167_ (.I(_117_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _168_ (.I(_117_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _169_ (.I(_117_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _170_ (.I(_117_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _171_ (.I(_113_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _172_ (.I(_118_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _173_ (.I(_118_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _174_ (.I(_118_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _175_ (.I(_118_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _176_ (.I(_118_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _177_ (.I(_118_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _178_ (.I(_118_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _179_ (.I(_118_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _180_ (.I(_118_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _181_ (.I(_118_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _182_ (.I(_113_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _183_ (.I(_119_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _184_ (.I(_119_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _185_ (.I(_119_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _186_ (.I(_119_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _187_ (.I(_119_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _188_ (.I(_119_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _189_ (.I(_119_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _190_ (.I(_119_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _191_ (.I(_119_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _192_ (.I(_119_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _193_ (.I(_113_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _194_ (.I(_120_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _195_ (.I(_120_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _196_ (.I(_120_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _197_ (.I(_120_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _198_ (.I(_120_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _199_ (.I(_120_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _200_ (.I(_120_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _201_ (.I(_120_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _202_ (.I(_120_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _203_ (.I(_120_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _204_ (.I(_113_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _205_ (.I(_121_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _206_ (.I(_121_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _207_ (.I(_121_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _208_ (.I(_121_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _209_ (.I(_121_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _210_ (.I(_121_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _211_ (.I(_121_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _212_ (.I(_121_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _213_ (.I(_121_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _214_ (.I(_121_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _215_ (.I(_112_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _216_ (.I(_122_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _217_ (.I(_122_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _218_ (.I(_122_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _219_ (.I(_122_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _220_ (.I(_122_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _221_ (.I(_122_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _222_ (.I(_122_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _223_ (.I(_122_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _224_ (.I(_122_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _225_ (.I(_122_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _226_ (.I(_112_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _227_ (.I(_123_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _228_ (.I(_123_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _229_ (.I(_123_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _230_ (.I(_123_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _231_ (.I(_123_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _232_ (.I(_123_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _233_ (.I(_123_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _234_ (.I(_123_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _235_ (.I(_123_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _236_ (.I(_123_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _237_ (.I(_112_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _238_ (.I(_124_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _239_ (.I(_124_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _240_ (.I(_124_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _241_ (.I(_124_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _242_ (.I(_124_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _243_ (.I(_124_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _244_ (.I(_124_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _245_ (.I(_124_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _246_ (.I(_124_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _247_ (.I(_124_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _248_ (.I(_113_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _249_ (.I(_113_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _250_ (.D(net105),
    .RN(_000_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _251_ (.D(net121),
    .RN(_001_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _252_ (.D(net133),
    .RN(_002_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _253_ (.D(net166),
    .RN(_003_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _254_ (.D(net156),
    .RN(_004_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _255_ (.D(net1),
    .RN(_005_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _256_ (.D(net127),
    .RN(_006_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _257_ (.D(net203),
    .RN(_007_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _258_ (.D(net201),
    .RN(_008_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _259_ (.D(net151),
    .RN(_009_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _260_ (.D(net116),
    .RN(_010_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _261_ (.D(net167),
    .RN(_011_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _262_ (.D(net107),
    .RN(_012_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_4.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _263_ (.D(net180),
    .RN(_013_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_4.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _264_ (.D(net192),
    .RN(_014_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_4.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _265_ (.D(net146),
    .RN(_015_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_4.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _266_ (.D(net145),
    .RN(_016_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_4.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _267_ (.D(net149),
    .RN(_017_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_4.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _268_ (.D(net131),
    .RN(_018_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_6.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _269_ (.D(net170),
    .RN(_019_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_6.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _270_ (.D(net119),
    .RN(_020_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_6.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _271_ (.D(net144),
    .RN(_021_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_6.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _272_ (.D(net172),
    .RN(_022_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_6.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _273_ (.D(net137),
    .RN(_023_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_6.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _274_ (.D(net138),
    .RN(_024_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_10.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _275_ (.D(net182),
    .RN(_025_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _276_ (.D(net191),
    .RN(_026_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_10.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _277_ (.D(net157),
    .RN(_027_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_10.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _278_ (.D(net108),
    .RN(_028_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_12.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _279_ (.D(net117),
    .RN(_029_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_12.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _280_ (.D(net143),
    .RN(_030_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_14.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _281_ (.D(net114),
    .RN(_031_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_14.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _282_ (.D(net102),
    .RN(_032_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _283_ (.D(net178),
    .RN(_033_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _284_ (.D(net161),
    .RN(_034_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_18.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _285_ (.D(net135),
    .RN(_035_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_18.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _286_ (.D(net158),
    .RN(_036_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_28.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _287_ (.D(net204),
    .RN(_037_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_28.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _288_ (.D(net103),
    .RN(_038_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _289_ (.D(net190),
    .RN(_039_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_38.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _290_ (.D(net183),
    .RN(_040_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_20.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _291_ (.D(net162),
    .RN(_041_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_20.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _292_ (.D(net132),
    .RN(_042_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_22.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _293_ (.D(net195),
    .RN(_043_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_22.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _294_ (.D(net169),
    .RN(_044_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _295_ (.D(net126),
    .RN(_045_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _296_ (.D(net194),
    .RN(_046_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_26.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _297_ (.D(net179),
    .RN(_047_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_26.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _298_ (.D(net124),
    .RN(_048_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _299_ (.D(net129),
    .RN(_049_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _300_ (.D(net98),
    .RN(_050_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _301_ (.D(net115),
    .RN(_051_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _302_ (.D(net109),
    .RN(_052_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _303_ (.D(net181),
    .RN(_053_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _304_ (.D(net113),
    .RN(_054_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _305_ (.D(net198),
    .RN(_055_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _306_ (.D(net99),
    .RN(_056_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _307_ (.D(net148),
    .RN(_057_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _308_ (.D(net185),
    .RN(_058_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _309_ (.D(net202),
    .RN(_059_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _310_ (.D(net177),
    .RN(_060_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _311_ (.D(net173),
    .RN(_061_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _312_ (.D(net150),
    .RN(_062_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _313_ (.D(net104),
    .RN(_063_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _314_ (.D(net197),
    .RN(_064_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _315_ (.D(net147),
    .RN(_065_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _316_ (.D(net171),
    .RN(_066_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _317_ (.D(net101),
    .RN(_067_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _318_ (.D(net125),
    .RN(_068_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _319_ (.D(net100),
    .RN(_069_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _320_ (.D(net139),
    .RN(_070_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _321_ (.D(net128),
    .RN(_071_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _322_ (.D(net154),
    .RN(_072_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _323_ (.D(net134),
    .RN(_073_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _324_ (.D(net153),
    .RN(_074_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _325_ (.D(net174),
    .RN(_075_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _326_ (.D(net97),
    .RN(_076_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _327_ (.D(net141),
    .RN(_077_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _328_ (.D(net184),
    .RN(_078_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _329_ (.D(net136),
    .RN(_079_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _330_ (.D(net142),
    .RN(_080_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _331_ (.D(net205),
    .RN(_081_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _332_ (.D(net168),
    .RN(_082_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _333_ (.D(net159),
    .RN(_083_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_32.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _334_ (.D(net106),
    .RN(_084_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_32.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _335_ (.D(net110),
    .RN(_085_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_32.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _336_ (.D(net111),
    .RN(_086_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_32.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _337_ (.D(net207),
    .RN(_087_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_32.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _338_ (.D(net155),
    .RN(_088_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _339_ (.D(net118),
    .RN(_089_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_9.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _340_ (.D(net176),
    .RN(_090_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_9.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _341_ (.D(net140),
    .RN(_091_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_9.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _342_ (.D(net152),
    .RN(_092_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_9.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _343_ (.D(net206),
    .RN(_093_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _344_ (.D(net112),
    .RN(_094_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _345_ (.D(net123),
    .RN(_095_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _346_ (.D(net164),
    .RN(_096_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _347_ (.D(net186),
    .RN(_097_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _348_ (.D(net163),
    .RN(_098_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _349_ (.D(net196),
    .RN(_099_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _350_ (.D(net160),
    .RN(_100_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _351_ (.D(net193),
    .RN(_101_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _352_ (.D(net200),
    .RN(_102_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _353_ (.D(net165),
    .RN(_103_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _354_ (.D(net189),
    .RN(_104_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _355_ (.D(net120),
    .RN(_105_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _356_ (.D(net175),
    .RN(_106_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _357_ (.D(net199),
    .RN(_107_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_33.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _358_ (.D(net122),
    .RN(_108_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_33.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _359_ (.D(net130),
    .RN(_109_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_33.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _360_ (.D(net188),
    .RN(_110_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_33.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _361_ (.D(net187),
    .RN(_111_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_left_track_33.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _389_ (.I(net27),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _390_ (.I(net26),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _391_ (.I(net25),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _392_ (.I(net24),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _393_ (.I(net23),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _394_ (.I(net22),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _395_ (.I(net21),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _396_ (.I(net34),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _397_ (.I(net33),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _398_ (.I(net32),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _399_ (.I(net31),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _400_ (.I(net30),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _401_ (.I(net29),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _402_ (.I(net28),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _403_ (.I(net20),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _404_ (.I(net11),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _405_ (.I(net10),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _406_ (.I(net9),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _407_ (.I(net7),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _408_ (.I(net6),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _409_ (.I(net5),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _410_ (.I(net3),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _411_ (.I(net19),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _412_ (.I(net18),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _413_ (.I(net17),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _414_ (.I(net16),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _415_ (.I(net15),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _416_ (.I(net14),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _417_ (.I(net13),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _418_ (.I(net2),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _419_ (.I(net4),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _420_ (.I(net8),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _421_ (.I(net12),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_4__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\mem_right_track_24.DFFR_4_.Q ),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\mem_right_track_32.DFFR_2_.Q ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(\mem_left_track_17.DFFR_0_.D ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(\mem_right_track_8.DFFR_4_.Q ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(\mem_right_track_0.DFFR_0_.D ),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(\mem_left_track_33.DFFR_3_.Q ),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(\mem_left_track_25.DFFR_2_.Q ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(\mem_top_track_2.DFFR_2_.Q ),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(\mem_left_track_1.DFFR_3_.Q ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(\mem_top_track_2.DFFR_3_.Q ),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold108 (.I(\mem_top_track_26.DFFR_1_.Q ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(\mem_right_track_16.DFFR_5_.Q ),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\mem_top_track_4.DFFR_4_.Q ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold110 (.I(\mem_left_track_1.DFFR_7_.Q ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold111 (.I(\mem_right_track_24.DFFR_5_.Q ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\mem_top_track_12.DFFR_0_.Q ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\mem_right_track_0.DFFR_2_.Q ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\mem_right_track_32.DFFR_1_.Q ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\mem_right_track_32.DFFR_0_.Q ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\mem_left_track_17.DFFR_4_.Q ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\mem_right_track_0.DFFR_0_.Q ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\mem_top_track_12.DFFR_1_.Q ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\mem_right_track_0.DFFR_3_.Q ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\mem_right_track_0.DFFR_4_.Q ),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\mem_top_track_2.DFFR_0_.Q ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\mem_top_track_10.DFFR_1_.Q ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\mem_left_track_9.DFFR_3_.Q ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\mem_top_track_6.DFFR_2_.Q ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\mem_left_track_17.DFFR_5_.Q ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\mem_top_track_0.DFFR_4_.Q ),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\mem_left_track_33.DFFR_2_.Q ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\mem_left_track_17.DFFR_3_.Q ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\mem_right_track_0.DFFR_6_.Q ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\mem_right_track_8.DFFR_0_.Q ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\mem_left_track_1.DFFR_6_.Q ),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\mem_top_track_22.DFFR_1_.Q ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\mem_top_track_2.DFFR_4_.Q ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\mem_right_track_16.DFFR_3_.Q ),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\mem_right_track_0.DFFR_5_.Q ),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\mem_left_track_33.DFFR_1_.Q ),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\mem_top_track_6.DFFR_4_.Q ),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\mem_top_track_22.DFFR_0_.Q ),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\mem_top_track_0.DFFR_1_.Q ),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\mem_right_track_16.DFFR_1_.Q ),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\mem_top_track_16.DFFR_1_.Q ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\mem_right_track_0.DFFR_7_.Q ),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\mem_right_track_24.DFFR_1_.Q ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\mem_top_track_4.DFFR_5_.Q ),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\mem_top_track_8.DFFR_0_.Q ),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\mem_right_track_16.DFFR_4_.Q ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\mem_left_track_9.DFFR_1_.Q ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\mem_right_track_24.DFFR_3_.Q ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\mem_right_track_24.DFFR_0_.Q ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\mem_top_track_14.DFFR_0_.Q ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(\mem_top_track_6.DFFR_1_.Q ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\mem_top_track_4.DFFR_0_.Q ),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\mem_right_track_8.DFFR_1_.Q ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(\mem_top_track_4.DFFR_1_.Q ),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\mem_right_track_8.DFFR_3_.Q ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(\mem_left_track_1.DFFR_5_.Q ),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\mem_top_track_2.DFFR_5_.Q ),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(\mem_left_track_1.DFFR_0_.Q ),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\mem_top_track_2.DFFR_1_.Q ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(\mem_left_track_9.DFFR_0_.Q ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\mem_right_track_16.DFFR_0_.Q ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(\mem_right_track_16.DFFR_2_.Q ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\mem_left_track_9.DFFR_4_.Q ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\mem_top_track_16.DFFR_0_.Q ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(\mem_top_track_0.DFFR_0_.Q ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\mem_top_track_10.DFFR_0_.D ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(\mem_top_track_28.DFFR_0_.Q ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\mem_right_track_32.DFFR_3_.Q ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(\mem_left_track_25.DFFR_4_.Q ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\mem_top_track_18.DFFR_0_.Q ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(\mem_top_track_18.DFFR_1_.Q ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\mem_left_track_17.DFFR_0_.Q ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(\mem_left_track_17.DFFR_2_.Q ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\mem_left_track_25.DFFR_1_.Q ),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\mem_top_track_38.DFFR_0_.Q ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(\mem_top_track_0.DFFR_2_.Q ),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\mem_top_track_0.DFFR_5_.Q ),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(\mem_right_track_32.DFFR_4_.Q ),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\mem_top_track_24.DFFR_0_.Q ),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(\mem_top_track_6.DFFR_3_.Q ),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\mem_right_track_8.DFFR_2_.Q ),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(\mem_top_track_6.DFFR_0_.Q ),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\mem_left_track_1.DFFR_1_.Q ),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(\mem_right_track_16.DFFR_0_.D ),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\mem_left_track_33.DFFR_4_.Q ),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\mem_left_track_1.DFFR_0_.D ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(\mem_left_track_9.DFFR_2_.Q ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\mem_left_track_1.DFFR_2_.Q ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(\mem_top_track_14.DFFR_1_.Q ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\mem_top_track_24.DFFR_1_.Q ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(\mem_top_track_4.DFFR_3_.Q ),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\mem_right_track_0.DFFR_1_.Q ),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(\mem_top_track_6.DFFR_5_.Q ),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\mem_top_track_20.DFFR_0_.Q ),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(\mem_right_track_24.DFFR_2_.Q ),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\mem_left_track_1.DFFR_4_.Q ),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\mem_top_track_0.DFFR_3_.Q ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(\mem_left_track_17.DFFR_1_.Q ),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\mem_left_track_25.DFFR_5_.Q ),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(\mem_left_track_33.DFFR_0_.Q ),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\mem_left_track_25.DFFR_0_.Q ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(\mem_top_track_28.DFFR_1_.Q ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(\mem_top_track_10.DFFR_0_.Q ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(\mem_top_track_4.DFFR_2_.Q ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(\mem_left_track_25.DFFR_3_.Q ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(\mem_top_track_26.DFFR_0_.Q ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(\mem_top_track_20.DFFR_1_.Q ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(chanx_left_in[17]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(chanx_left_in[18]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(chanx_left_in[19]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(chanx_left_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(chanx_left_in[2]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(chanx_left_in[4]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(chanx_left_in[5]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(chanx_left_in[6]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(chanx_left_in[8]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(chanx_left_in[9]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(chanx_left_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(chanx_right_in[0]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(chanx_right_in[10]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(chanx_right_in[12]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(chanx_right_in[13]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(chanx_right_in[14]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(chanx_right_in[16]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(chanx_right_in[17]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(chanx_right_in[18]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(chanx_right_in[1]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(chanx_right_in[2]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(chanx_left_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(chanx_right_in[4]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(chanx_right_in[5]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(chanx_right_in[6]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(chanx_right_in[8]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(chanx_right_in[9]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(pReset),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(chanx_left_in[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(chanx_left_in[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(chanx_left_in[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(chanx_left_in[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(chanx_left_in[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(chanx_left_in[16]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output36 (.I(net36),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(chanx_left_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(chanx_left_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output39 (.I(net39),
    .Z(chanx_left_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output40 (.I(net40),
    .Z(chanx_left_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output41 (.I(net41),
    .Z(chanx_left_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(chanx_left_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output43 (.I(net43),
    .Z(chanx_left_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output44 (.I(net44),
    .Z(chanx_left_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(chanx_left_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(chanx_left_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output47 (.I(net47),
    .Z(chanx_left_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output48 (.I(net48),
    .Z(chanx_left_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(chanx_left_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output50 (.I(net50),
    .Z(chanx_left_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(chanx_left_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output52 (.I(net52),
    .Z(chanx_right_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output53 (.I(net53),
    .Z(chanx_right_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output54 (.I(net54),
    .Z(chanx_right_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output55 (.I(net55),
    .Z(chanx_right_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output56 (.I(net56),
    .Z(chanx_right_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(chanx_right_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output58 (.I(net58),
    .Z(chanx_right_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output59 (.I(net59),
    .Z(chanx_right_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output60 (.I(net60),
    .Z(chanx_right_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output61 (.I(net61),
    .Z(chanx_right_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output62 (.I(net62),
    .Z(chanx_right_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output63 (.I(net63),
    .Z(chanx_right_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(chanx_right_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output65 (.I(net65),
    .Z(chanx_right_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output66 (.I(net66),
    .Z(chanx_right_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output67 (.I(net67),
    .Z(chany_top_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(chany_top_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output69 (.I(net69),
    .Z(chany_top_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_1__0__96 (.ZN(net96));
 assign chanx_left_out[0] = net96;
 assign chanx_left_out[12] = net93;
 assign chanx_left_out[16] = net92;
 assign chanx_left_out[4] = net95;
 assign chanx_left_out[8] = net94;
 assign chanx_right_out[0] = net91;
 assign chanx_right_out[12] = net88;
 assign chanx_right_out[16] = net87;
 assign chanx_right_out[4] = net90;
 assign chanx_right_out[8] = net89;
 assign chany_top_out[0] = net86;
 assign chany_top_out[10] = net76;
 assign chany_top_out[11] = net75;
 assign chany_top_out[12] = net74;
 assign chany_top_out[13] = net73;
 assign chany_top_out[14] = net72;
 assign chany_top_out[15] = net71;
 assign chany_top_out[19] = net70;
 assign chany_top_out[1] = net85;
 assign chany_top_out[2] = net84;
 assign chany_top_out[3] = net83;
 assign chany_top_out[4] = net82;
 assign chany_top_out[5] = net81;
 assign chany_top_out[6] = net80;
 assign chany_top_out[7] = net79;
 assign chany_top_out[8] = net78;
 assign chany_top_out[9] = net77;
endmodule

