// This is the unpowered netlist.
module cby_1__1_ (ccff_head,
    ccff_tail,
    left_grid_right_width_0_height_0_subtile_0__pin_I_1_,
    left_grid_right_width_0_height_0_subtile_0__pin_I_5_,
    left_grid_right_width_0_height_0_subtile_0__pin_I_9_,
    pReset,
    prog_clk,
    right_grid_left_width_0_height_0_subtile_0__pin_I_11_,
    right_grid_left_width_0_height_0_subtile_0__pin_I_3_,
    right_grid_left_width_0_height_0_subtile_0__pin_I_7_,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input ccff_head;
 output ccff_tail;
 output left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
 output left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
 output left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
 input pReset;
 input prog_clk;
 output right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
 output right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
 output right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
 input [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;
 input [19:0] chany_top_in;
 output [19:0] chany_top_out;

 wire net86;
 wire net85;
 wire net84;
 wire net87;
 wire net88;
 wire net89;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire clknet_0_prog_clk;
 wire clknet_2_0__leaf_prog_clk;
 wire clknet_2_1__leaf_prog_clk;
 wire clknet_2_2__leaf_prog_clk;
 wire clknet_2_3__leaf_prog_clk;
 wire \mem_left_ipin_0.DFFR_0_.Q ;
 wire \mem_left_ipin_0.DFFR_1_.Q ;
 wire \mem_left_ipin_0.DFFR_2_.Q ;
 wire \mem_left_ipin_0.DFFR_3_.Q ;
 wire \mem_left_ipin_0.DFFR_4_.Q ;
 wire \mem_left_ipin_0.DFFR_5_.Q ;
 wire \mem_left_ipin_1.DFFR_0_.Q ;
 wire \mem_left_ipin_1.DFFR_1_.Q ;
 wire \mem_left_ipin_1.DFFR_2_.Q ;
 wire \mem_left_ipin_1.DFFR_3_.Q ;
 wire \mem_left_ipin_1.DFFR_4_.Q ;
 wire \mem_left_ipin_1.DFFR_5_.Q ;
 wire \mem_left_ipin_2.DFFR_0_.Q ;
 wire \mem_left_ipin_2.DFFR_1_.Q ;
 wire \mem_left_ipin_2.DFFR_2_.Q ;
 wire \mem_left_ipin_2.DFFR_3_.Q ;
 wire \mem_left_ipin_2.DFFR_4_.Q ;
 wire \mem_left_ipin_2.DFFR_5_.Q ;
 wire \mem_right_ipin_0.DFFR_0_.Q ;
 wire \mem_right_ipin_0.DFFR_1_.Q ;
 wire \mem_right_ipin_0.DFFR_2_.Q ;
 wire \mem_right_ipin_0.DFFR_3_.Q ;
 wire \mem_right_ipin_0.DFFR_4_.Q ;
 wire \mem_right_ipin_0.DFFR_5_.Q ;
 wire \mem_right_ipin_1.DFFR_0_.Q ;
 wire \mem_right_ipin_1.DFFR_1_.Q ;
 wire \mem_right_ipin_1.DFFR_2_.Q ;
 wire \mem_right_ipin_1.DFFR_3_.Q ;
 wire \mem_right_ipin_1.DFFR_4_.Q ;
 wire \mem_right_ipin_1.DFFR_5_.Q ;
 wire \mem_right_ipin_2.DFFR_0_.Q ;
 wire \mem_right_ipin_2.DFFR_1_.Q ;
 wire \mem_right_ipin_2.DFFR_2_.Q ;
 wire \mem_right_ipin_2.DFFR_3_.Q ;
 wire \mem_right_ipin_2.DFFR_4_.Q ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__064__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__065__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__066__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__067__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__068__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__069__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__070__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__071__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__072__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__073__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__CLK (.I(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(chany_bottom_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(chany_bottom_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(chany_bottom_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(chany_bottom_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(chany_bottom_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(chany_bottom_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(chany_bottom_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(chany_bottom_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(chany_bottom_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(chany_bottom_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(chany_bottom_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(chany_bottom_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(chany_top_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(chany_top_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(chany_top_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(chany_top_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(chany_top_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(chany_top_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(chany_top_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(chany_top_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(chany_bottom_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(chany_top_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(chany_top_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(chany_top_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(chany_top_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(chany_top_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(chany_top_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(chany_top_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(chany_top_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(chany_top_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(chany_top_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(chany_bottom_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(chany_top_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(chany_top_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(chany_bottom_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(chany_bottom_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(chany_bottom_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(chany_bottom_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(chany_bottom_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(chany_bottom_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_93 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _040_ (.I(net42),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _041_ (.I(_036_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _042_ (.I(_037_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _043_ (.I(_037_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _044_ (.I(_037_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _045_ (.I(_037_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _046_ (.I(_037_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _047_ (.I(_037_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _048_ (.I(_037_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _049_ (.I(_037_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _050_ (.I(_037_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _051_ (.I(_037_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _052_ (.I(_036_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _053_ (.I(_038_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _054_ (.I(_038_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _055_ (.I(_038_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _056_ (.I(_038_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _057_ (.I(_038_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _058_ (.I(_038_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _059_ (.I(_038_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _060_ (.I(_038_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _061_ (.I(_038_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _062_ (.I(_038_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _063_ (.I(_036_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _064_ (.I(_039_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _065_ (.I(_039_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _066_ (.I(_039_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _067_ (.I(_039_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _068_ (.I(_039_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _069_ (.I(_039_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _070_ (.I(_039_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _071_ (.I(_039_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _072_ (.I(_039_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _073_ (.I(_039_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _074_ (.I(_036_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _075_ (.I(_036_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _076_ (.I(_036_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _077_ (.I(_036_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _078_ (.I(_036_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _079_ (.I(_036_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _080_ (.D(net98),
    .RN(_000_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_left_ipin_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _081_ (.D(net108),
    .RN(_001_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_left_ipin_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _082_ (.D(net112),
    .RN(_002_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_left_ipin_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _083_ (.D(net117),
    .RN(_003_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_left_ipin_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _084_ (.D(net123),
    .RN(_004_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_left_ipin_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _085_ (.D(net1),
    .RN(_005_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_left_ipin_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _086_ (.D(net99),
    .RN(_006_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _087_ (.D(net107),
    .RN(_007_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _088_ (.D(net111),
    .RN(_008_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _089_ (.D(net95),
    .RN(_009_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _090_ (.D(net91),
    .RN(_010_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_left_ipin_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _091_ (.D(net93),
    .RN(_011_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _092_ (.D(net103),
    .RN(_012_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_left_ipin_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _093_ (.D(net110),
    .RN(_013_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_left_ipin_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _094_ (.D(net90),
    .RN(_014_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_left_ipin_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _095_ (.D(net106),
    .RN(_015_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _096_ (.D(net105),
    .RN(_016_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _097_ (.D(net100),
    .RN(_017_),
    .CLK(clknet_2_1__leaf_prog_clk),
    .Q(\mem_left_ipin_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _098_ (.D(net94),
    .RN(_018_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _099_ (.D(net104),
    .RN(_019_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_ipin_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _100_ (.D(net116),
    .RN(_020_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_ipin_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _101_ (.D(net119),
    .RN(_021_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_ipin_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _102_ (.D(net120),
    .RN(_022_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_ipin_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _103_ (.D(net97),
    .RN(_023_),
    .CLK(clknet_2_3__leaf_prog_clk),
    .Q(\mem_right_ipin_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _104_ (.D(net122),
    .RN(_024_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _105_ (.D(net118),
    .RN(_025_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _106_ (.D(net102),
    .RN(_026_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _107_ (.D(net121),
    .RN(_027_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _108_ (.D(net114),
    .RN(_028_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _109_ (.D(net109),
    .RN(_029_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _110_ (.D(net101),
    .RN(_030_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _111_ (.D(net92),
    .RN(_031_),
    .CLK(clknet_2_2__leaf_prog_clk),
    .Q(\mem_right_ipin_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _112_ (.D(net115),
    .RN(_032_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_ipin_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _113_ (.D(net96),
    .RN(_033_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_ipin_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _114_ (.D(net113),
    .RN(_034_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_ipin_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _115_ (.D(net124),
    .RN(_035_),
    .CLK(clknet_2_0__leaf_prog_clk),
    .Q(\mem_right_ipin_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _122_ (.I(net32),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _123_ (.I(net31),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _124_ (.I(net30),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _125_ (.I(net29),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _126_ (.I(net28),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _127_ (.I(net27),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _128_ (.I(net26),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _129_ (.I(net25),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _130_ (.I(net24),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _131_ (.I(net23),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _132_ (.I(net41),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _133_ (.I(net40),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _134_ (.I(net39),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _135_ (.I(net38),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _136_ (.I(net37),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _137_ (.I(net36),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _138_ (.I(net35),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _139_ (.I(net34),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _140_ (.I(net33),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _141_ (.I(net22),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _142_ (.I(net12),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _143_ (.I(net11),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _144_ (.I(net10),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _145_ (.I(net9),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _146_ (.I(net8),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _147_ (.I(net7),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _148_ (.I(net6),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _149_ (.I(net5),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _150_ (.I(net4),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _151_ (.I(net3),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _152_ (.I(net21),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _153_ (.I(net20),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _154_ (.I(net19),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _155_ (.I(net18),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _156_ (.I(net17),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _157_ (.I(net16),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _158_ (.I(net15),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _159_ (.I(net14),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _160_ (.I(net13),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _161_ (.I(net2),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel cby_1__1__84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel cby_1__1__85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel cby_1__1__86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel cby_1__1__87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel cby_1__1__88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel cby_1__1__89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_2_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\mem_left_ipin_2.DFFR_2_.Q ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\mem_left_ipin_1.DFFR_4_.Q ),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\mem_left_ipin_1.DFFR_5_.Q ),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\mem_right_ipin_2.DFFR_4_.Q ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\mem_right_ipin_1.DFFR_2_.Q ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\mem_left_ipin_2.DFFR_4_.Q ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\mem_right_ipin_0.DFFR_3_.Q ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\mem_left_ipin_2.DFFR_0_.Q ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\mem_left_ipin_2.DFFR_1_.Q ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\mem_left_ipin_1.DFFR_3_.Q ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\mem_left_ipin_0.DFFR_3_.Q ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\mem_left_ipin_1.DFFR_0_.Q ),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\mem_right_ipin_0.DFFR_5_.Q ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\mem_left_ipin_2.DFFR_3_.Q ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\mem_left_ipin_1.DFFR_2_.Q ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\mem_left_ipin_0.DFFR_2_.Q ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\mem_right_ipin_2.DFFR_0_.Q ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\mem_right_ipin_1.DFFR_0_.Q ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\mem_right_ipin_2.DFFR_2_.Q ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\mem_right_ipin_0.DFFR_2_.Q ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\mem_left_ipin_0.DFFR_1_.Q ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\mem_right_ipin_1.DFFR_3_.Q ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\mem_right_ipin_2.DFFR_3_.Q ),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\mem_right_ipin_0.DFFR_1_.Q ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\mem_right_ipin_0.DFFR_0_.Q ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\mem_right_ipin_1.DFFR_1_.Q ),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\mem_right_ipin_1.DFFR_4_.Q ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\mem_left_ipin_0.DFFR_0_.Q ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\mem_right_ipin_1.DFFR_5_.Q ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\mem_left_ipin_0.DFFR_5_.Q ),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\mem_right_ipin_0.DFFR_4_.Q ),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\mem_left_ipin_1.DFFR_1_.Q ),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\mem_right_ipin_2.DFFR_1_.Q ),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\mem_left_ipin_2.DFFR_5_.Q ),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\mem_left_ipin_0.DFFR_4_.Q ),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(chany_bottom_in[17]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(chany_bottom_in[18]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(chany_bottom_in[19]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(chany_bottom_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(chany_bottom_in[2]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(chany_bottom_in[3]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(chany_bottom_in[4]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(chany_bottom_in[5]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(chany_bottom_in[6]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(chany_bottom_in[7]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(chany_bottom_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(chany_bottom_in[8]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(chany_bottom_in[9]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(chany_top_in[0]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(chany_top_in[10]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(chany_top_in[11]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(chany_top_in[12]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(chany_top_in[13]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(chany_top_in[14]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(chany_top_in[15]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(chany_top_in[16]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(chany_bottom_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(chany_top_in[17]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(chany_top_in[18]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(chany_top_in[19]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(chany_top_in[1]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(chany_top_in[2]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(chany_top_in[3]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(chany_top_in[4]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(chany_top_in[5]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(chany_top_in[6]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(chany_top_in[7]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(chany_bottom_in[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(chany_top_in[8]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(chany_top_in[9]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input42 (.I(pReset),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(chany_bottom_in[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(chany_bottom_in[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(chany_bottom_in[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(chany_bottom_in[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(chany_bottom_in[16]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output43 (.I(net43),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output44 (.I(net44),
    .Z(chany_bottom_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output45 (.I(net45),
    .Z(chany_bottom_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output46 (.I(net46),
    .Z(chany_bottom_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output47 (.I(net47),
    .Z(chany_bottom_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output48 (.I(net48),
    .Z(chany_bottom_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(chany_bottom_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output50 (.I(net50),
    .Z(chany_bottom_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output51 (.I(net51),
    .Z(chany_bottom_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output52 (.I(net52),
    .Z(chany_bottom_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output53 (.I(net53),
    .Z(chany_bottom_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output54 (.I(net54),
    .Z(chany_bottom_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output55 (.I(net55),
    .Z(chany_bottom_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output56 (.I(net56),
    .Z(chany_bottom_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output57 (.I(net57),
    .Z(chany_bottom_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output58 (.I(net58),
    .Z(chany_bottom_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output59 (.I(net59),
    .Z(chany_bottom_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output60 (.I(net60),
    .Z(chany_bottom_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output61 (.I(net61),
    .Z(chany_bottom_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output62 (.I(net62),
    .Z(chany_bottom_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output63 (.I(net63),
    .Z(chany_bottom_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output64 (.I(net64),
    .Z(chany_top_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output65 (.I(net65),
    .Z(chany_top_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output66 (.I(net66),
    .Z(chany_top_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(chany_top_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(chany_top_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output69 (.I(net69),
    .Z(chany_top_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output70 (.I(net70),
    .Z(chany_top_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(chany_top_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output72 (.I(net72),
    .Z(chany_top_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output73 (.I(net73),
    .Z(chany_top_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output74 (.I(net74),
    .Z(chany_top_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output75 (.I(net75),
    .Z(chany_top_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output76 (.I(net76),
    .Z(chany_top_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output77 (.I(net77),
    .Z(chany_top_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output78 (.I(net78),
    .Z(chany_top_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output79 (.I(net79),
    .Z(chany_top_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output80 (.I(net80),
    .Z(chany_top_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output81 (.I(net81),
    .Z(chany_top_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output82 (.I(net82),
    .Z(chany_top_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(chany_top_out[9]));
 assign left_grid_right_width_0_height_0_subtile_0__pin_I_1_ = net86;
 assign left_grid_right_width_0_height_0_subtile_0__pin_I_5_ = net85;
 assign left_grid_right_width_0_height_0_subtile_0__pin_I_9_ = net84;
 assign right_grid_left_width_0_height_0_subtile_0__pin_I_11_ = net87;
 assign right_grid_left_width_0_height_0_subtile_0__pin_I_3_ = net88;
 assign right_grid_left_width_0_height_0_subtile_0__pin_I_7_ = net89;
endmodule

