magic
tech gf180mcuD
magscale 1 10
timestamp 1702149169
<< metal1 >>
rect 13458 27806 13470 27858
rect 13522 27855 13534 27858
rect 14130 27855 14142 27858
rect 13522 27809 14142 27855
rect 13522 27806 13534 27809
rect 14130 27806 14142 27809
rect 14194 27806 14206 27858
rect 10098 26798 10110 26850
rect 10162 26847 10174 26850
rect 11106 26847 11118 26850
rect 10162 26801 11118 26847
rect 10162 26798 10174 26801
rect 11106 26798 11118 26801
rect 11170 26798 11182 26850
rect 16818 26798 16830 26850
rect 16882 26847 16894 26850
rect 17490 26847 17502 26850
rect 16882 26801 17502 26847
rect 16882 26798 16894 26801
rect 17490 26798 17502 26801
rect 17554 26798 17566 26850
rect 18834 26798 18846 26850
rect 18898 26847 18910 26850
rect 19618 26847 19630 26850
rect 18898 26801 19630 26847
rect 18898 26798 18910 26801
rect 19618 26798 19630 26801
rect 19682 26798 19694 26850
rect 22194 26798 22206 26850
rect 22258 26847 22270 26850
rect 22978 26847 22990 26850
rect 22258 26801 22990 26847
rect 22258 26798 22270 26801
rect 22978 26798 22990 26801
rect 23042 26798 23054 26850
rect 1344 26682 28720 26716
rect 1344 26630 8018 26682
rect 8070 26630 8122 26682
rect 8174 26630 8226 26682
rect 8278 26630 14822 26682
rect 14874 26630 14926 26682
rect 14978 26630 15030 26682
rect 15082 26630 21626 26682
rect 21678 26630 21730 26682
rect 21782 26630 21834 26682
rect 21886 26630 28430 26682
rect 28482 26630 28534 26682
rect 28586 26630 28638 26682
rect 28690 26630 28720 26682
rect 1344 26596 28720 26630
rect 7646 26514 7698 26526
rect 7646 26450 7698 26462
rect 8206 26514 8258 26526
rect 8206 26450 8258 26462
rect 8766 26514 8818 26526
rect 8766 26450 8818 26462
rect 11118 26514 11170 26526
rect 11118 26450 11170 26462
rect 12014 26514 12066 26526
rect 12014 26450 12066 26462
rect 13358 26514 13410 26526
rect 13358 26450 13410 26462
rect 23886 26514 23938 26526
rect 23886 26450 23938 26462
rect 25118 26514 25170 26526
rect 25118 26450 25170 26462
rect 9662 26402 9714 26414
rect 9662 26338 9714 26350
rect 12238 26402 12290 26414
rect 12238 26338 12290 26350
rect 12574 26402 12626 26414
rect 12574 26338 12626 26350
rect 15374 26402 15426 26414
rect 15374 26338 15426 26350
rect 16046 26402 16098 26414
rect 16046 26338 16098 26350
rect 26238 26402 26290 26414
rect 26238 26338 26290 26350
rect 10334 26290 10386 26302
rect 9874 26238 9886 26290
rect 9938 26238 9950 26290
rect 10334 26226 10386 26238
rect 13694 26290 13746 26302
rect 17054 26290 17106 26302
rect 20750 26290 20802 26302
rect 15586 26238 15598 26290
rect 15650 26238 15662 26290
rect 16258 26238 16270 26290
rect 16322 26238 16334 26290
rect 18722 26238 18734 26290
rect 18786 26238 18798 26290
rect 13694 26226 13746 26238
rect 17054 26226 17106 26238
rect 20750 26226 20802 26238
rect 22318 26290 22370 26302
rect 26786 26238 26798 26290
rect 26850 26238 26862 26290
rect 22318 26226 22370 26238
rect 14130 26126 14142 26178
rect 14194 26126 14206 26178
rect 17490 26126 17502 26178
rect 17554 26126 17566 26178
rect 19058 26126 19070 26178
rect 19122 26126 19134 26178
rect 21186 26126 21198 26178
rect 21250 26126 21262 26178
rect 22754 26126 22766 26178
rect 22818 26126 22830 26178
rect 27682 26126 27694 26178
rect 27746 26126 27758 26178
rect 1344 25898 28560 25932
rect 1344 25846 4616 25898
rect 4668 25846 4720 25898
rect 4772 25846 4824 25898
rect 4876 25846 11420 25898
rect 11472 25846 11524 25898
rect 11576 25846 11628 25898
rect 11680 25846 18224 25898
rect 18276 25846 18328 25898
rect 18380 25846 18432 25898
rect 18484 25846 25028 25898
rect 25080 25846 25132 25898
rect 25184 25846 25236 25898
rect 25288 25846 28560 25898
rect 1344 25812 28560 25846
rect 9438 25618 9490 25630
rect 9438 25554 9490 25566
rect 10782 25618 10834 25630
rect 15934 25618 15986 25630
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 10782 25554 10834 25566
rect 15934 25554 15986 25566
rect 17166 25618 17218 25630
rect 19630 25618 19682 25630
rect 18946 25566 18958 25618
rect 19010 25566 19022 25618
rect 17166 25554 17218 25566
rect 19630 25554 19682 25566
rect 11006 25506 11058 25518
rect 11006 25442 11058 25454
rect 12574 25506 12626 25518
rect 22990 25506 23042 25518
rect 16482 25454 16494 25506
rect 16546 25454 16558 25506
rect 18498 25454 18510 25506
rect 18562 25454 18574 25506
rect 20178 25454 20190 25506
rect 20242 25454 20254 25506
rect 21410 25454 21422 25506
rect 21474 25454 21486 25506
rect 22194 25454 22206 25506
rect 22258 25454 22270 25506
rect 12574 25442 12626 25454
rect 22990 25442 23042 25454
rect 27134 25506 27186 25518
rect 27134 25442 27186 25454
rect 28142 25506 28194 25518
rect 28142 25442 28194 25454
rect 11678 25394 11730 25406
rect 11678 25330 11730 25342
rect 12910 25394 12962 25406
rect 12910 25330 12962 25342
rect 15038 25394 15090 25406
rect 15038 25330 15090 25342
rect 16718 25394 16770 25406
rect 16718 25330 16770 25342
rect 20638 25394 20690 25406
rect 20638 25330 20690 25342
rect 21646 25394 21698 25406
rect 21646 25330 21698 25342
rect 22654 25394 22706 25406
rect 22654 25330 22706 25342
rect 1710 25282 1762 25294
rect 1710 25218 1762 25230
rect 11342 25282 11394 25294
rect 11342 25218 11394 25230
rect 13470 25282 13522 25294
rect 13470 25218 13522 25230
rect 19966 25282 20018 25294
rect 19966 25218 20018 25230
rect 21982 25282 22034 25294
rect 21982 25218 22034 25230
rect 27470 25282 27522 25294
rect 27470 25218 27522 25230
rect 27806 25282 27858 25294
rect 27806 25218 27858 25230
rect 1344 25114 28720 25148
rect 1344 25062 8018 25114
rect 8070 25062 8122 25114
rect 8174 25062 8226 25114
rect 8278 25062 14822 25114
rect 14874 25062 14926 25114
rect 14978 25062 15030 25114
rect 15082 25062 21626 25114
rect 21678 25062 21730 25114
rect 21782 25062 21834 25114
rect 21886 25062 28430 25114
rect 28482 25062 28534 25114
rect 28586 25062 28638 25114
rect 28690 25062 28720 25114
rect 1344 25028 28720 25062
rect 13134 24946 13186 24958
rect 13134 24882 13186 24894
rect 21758 24946 21810 24958
rect 21758 24882 21810 24894
rect 22430 24946 22482 24958
rect 22430 24882 22482 24894
rect 27022 24946 27074 24958
rect 27022 24882 27074 24894
rect 12798 24834 12850 24846
rect 12798 24770 12850 24782
rect 27358 24834 27410 24846
rect 27358 24770 27410 24782
rect 28142 24834 28194 24846
rect 28142 24770 28194 24782
rect 1344 24330 28560 24364
rect 1344 24278 4616 24330
rect 4668 24278 4720 24330
rect 4772 24278 4824 24330
rect 4876 24278 11420 24330
rect 11472 24278 11524 24330
rect 11576 24278 11628 24330
rect 11680 24278 18224 24330
rect 18276 24278 18328 24330
rect 18380 24278 18432 24330
rect 18484 24278 25028 24330
rect 25080 24278 25132 24330
rect 25184 24278 25236 24330
rect 25288 24278 28560 24330
rect 1344 24244 28560 24278
rect 9314 23886 9326 23938
rect 9378 23886 9390 23938
rect 18834 23886 18846 23938
rect 18898 23886 18910 23938
rect 9550 23826 9602 23838
rect 9550 23762 9602 23774
rect 19070 23826 19122 23838
rect 19070 23762 19122 23774
rect 27694 23714 27746 23726
rect 27694 23650 27746 23662
rect 28142 23714 28194 23726
rect 28142 23650 28194 23662
rect 1344 23546 28720 23580
rect 1344 23494 8018 23546
rect 8070 23494 8122 23546
rect 8174 23494 8226 23546
rect 8278 23494 14822 23546
rect 14874 23494 14926 23546
rect 14978 23494 15030 23546
rect 15082 23494 21626 23546
rect 21678 23494 21730 23546
rect 21782 23494 21834 23546
rect 21886 23494 28430 23546
rect 28482 23494 28534 23546
rect 28586 23494 28638 23546
rect 28690 23494 28720 23546
rect 1344 23460 28720 23494
rect 27134 23266 27186 23278
rect 27134 23202 27186 23214
rect 27470 23266 27522 23278
rect 27470 23202 27522 23214
rect 27806 23266 27858 23278
rect 27806 23202 27858 23214
rect 28142 23154 28194 23166
rect 28142 23090 28194 23102
rect 26910 23042 26962 23054
rect 26910 22978 26962 22990
rect 1344 22762 28560 22796
rect 1344 22710 4616 22762
rect 4668 22710 4720 22762
rect 4772 22710 4824 22762
rect 4876 22710 11420 22762
rect 11472 22710 11524 22762
rect 11576 22710 11628 22762
rect 11680 22710 18224 22762
rect 18276 22710 18328 22762
rect 18380 22710 18432 22762
rect 18484 22710 25028 22762
rect 25080 22710 25132 22762
rect 25184 22710 25236 22762
rect 25288 22710 28560 22762
rect 1344 22676 28560 22710
rect 27122 22318 27134 22370
rect 27186 22318 27198 22370
rect 28018 22206 28030 22258
rect 28082 22206 28094 22258
rect 1344 21978 28720 22012
rect 1344 21926 8018 21978
rect 8070 21926 8122 21978
rect 8174 21926 8226 21978
rect 8278 21926 14822 21978
rect 14874 21926 14926 21978
rect 14978 21926 15030 21978
rect 15082 21926 21626 21978
rect 21678 21926 21730 21978
rect 21782 21926 21834 21978
rect 21886 21926 28430 21978
rect 28482 21926 28534 21978
rect 28586 21926 28638 21978
rect 28690 21926 28720 21978
rect 1344 21892 28720 21926
rect 15710 21810 15762 21822
rect 15710 21746 15762 21758
rect 15374 21698 15426 21710
rect 15374 21634 15426 21646
rect 16046 21698 16098 21710
rect 16046 21634 16098 21646
rect 16382 21698 16434 21710
rect 27234 21646 27246 21698
rect 27298 21646 27310 21698
rect 16382 21634 16434 21646
rect 26014 21474 26066 21486
rect 26226 21422 26238 21474
rect 26290 21422 26302 21474
rect 26014 21410 26066 21422
rect 1344 21194 28560 21228
rect 1344 21142 4616 21194
rect 4668 21142 4720 21194
rect 4772 21142 4824 21194
rect 4876 21142 11420 21194
rect 11472 21142 11524 21194
rect 11576 21142 11628 21194
rect 11680 21142 18224 21194
rect 18276 21142 18328 21194
rect 18380 21142 18432 21194
rect 18484 21142 25028 21194
rect 25080 21142 25132 21194
rect 25184 21142 25236 21194
rect 25288 21142 28560 21194
rect 1344 21108 28560 21142
rect 22990 20802 23042 20814
rect 23650 20750 23662 20802
rect 23714 20750 23726 20802
rect 27794 20750 27806 20802
rect 27858 20750 27870 20802
rect 22990 20738 23042 20750
rect 27246 20690 27298 20702
rect 26898 20638 26910 20690
rect 26962 20638 26974 20690
rect 27570 20638 27582 20690
rect 27634 20638 27646 20690
rect 27246 20626 27298 20638
rect 17278 20578 17330 20590
rect 26686 20578 26738 20590
rect 26114 20526 26126 20578
rect 26178 20526 26190 20578
rect 17278 20514 17330 20526
rect 26686 20514 26738 20526
rect 1344 20410 28720 20444
rect 1344 20358 8018 20410
rect 8070 20358 8122 20410
rect 8174 20358 8226 20410
rect 8278 20358 14822 20410
rect 14874 20358 14926 20410
rect 14978 20358 15030 20410
rect 15082 20358 21626 20410
rect 21678 20358 21730 20410
rect 21782 20358 21834 20410
rect 21886 20358 28430 20410
rect 28482 20358 28534 20410
rect 28586 20358 28638 20410
rect 28690 20358 28720 20410
rect 1344 20324 28720 20358
rect 22766 20242 22818 20254
rect 22766 20178 22818 20190
rect 28142 20242 28194 20254
rect 28142 20178 28194 20190
rect 21646 20130 21698 20142
rect 11778 20078 11790 20130
rect 11842 20078 11854 20130
rect 14018 20078 14030 20130
rect 14082 20078 14094 20130
rect 16258 20078 16270 20130
rect 16322 20078 16334 20130
rect 13918 20018 13970 20030
rect 14033 20015 14079 20078
rect 21646 20066 21698 20078
rect 22430 20130 22482 20142
rect 27234 20078 27246 20130
rect 27298 20078 27310 20130
rect 22430 20066 22482 20078
rect 18958 20018 19010 20030
rect 25902 20018 25954 20030
rect 14242 20015 14254 20018
rect 14033 19969 14254 20015
rect 14242 19966 14254 19969
rect 14306 19966 14318 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 13918 19954 13970 19966
rect 18958 19954 19010 19966
rect 25902 19954 25954 19966
rect 14366 19906 14418 19918
rect 17614 19906 17666 19918
rect 10658 19854 10670 19906
rect 10722 19854 10734 19906
rect 13570 19854 13582 19906
rect 13634 19854 13646 19906
rect 15250 19854 15262 19906
rect 15314 19854 15326 19906
rect 17826 19854 17838 19906
rect 17890 19854 17902 19906
rect 26226 19854 26238 19906
rect 26290 19854 26302 19906
rect 14366 19842 14418 19854
rect 17614 19842 17666 19854
rect 1344 19626 28560 19660
rect 1344 19574 4616 19626
rect 4668 19574 4720 19626
rect 4772 19574 4824 19626
rect 4876 19574 11420 19626
rect 11472 19574 11524 19626
rect 11576 19574 11628 19626
rect 11680 19574 18224 19626
rect 18276 19574 18328 19626
rect 18380 19574 18432 19626
rect 18484 19574 25028 19626
rect 25080 19574 25132 19626
rect 25184 19574 25236 19626
rect 25288 19574 28560 19626
rect 1344 19540 28560 19574
rect 24894 19458 24946 19470
rect 24894 19394 24946 19406
rect 8642 19294 8654 19346
rect 8706 19294 8718 19346
rect 11442 19294 11454 19346
rect 11506 19294 11518 19346
rect 18274 19294 18286 19346
rect 18338 19294 18350 19346
rect 26674 19294 26686 19346
rect 26738 19294 26750 19346
rect 21422 19234 21474 19246
rect 13458 19182 13470 19234
rect 13522 19182 13534 19234
rect 14018 19182 14030 19234
rect 14082 19182 14094 19234
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 21422 19170 21474 19182
rect 17054 19122 17106 19134
rect 9650 19070 9662 19122
rect 9714 19070 9726 19122
rect 12450 19070 12462 19122
rect 12514 19070 12526 19122
rect 19282 19070 19294 19122
rect 19346 19070 19358 19122
rect 27682 19070 27694 19122
rect 27746 19070 27758 19122
rect 17054 19058 17106 19070
rect 25230 19010 25282 19022
rect 16258 18958 16270 19010
rect 16322 18958 16334 19010
rect 24098 18958 24110 19010
rect 24162 18958 24174 19010
rect 25230 18946 25282 18958
rect 1344 18842 28720 18876
rect 1344 18790 8018 18842
rect 8070 18790 8122 18842
rect 8174 18790 8226 18842
rect 8278 18790 14822 18842
rect 14874 18790 14926 18842
rect 14978 18790 15030 18842
rect 15082 18790 21626 18842
rect 21678 18790 21730 18842
rect 21782 18790 21834 18842
rect 21886 18790 28430 18842
rect 28482 18790 28534 18842
rect 28586 18790 28638 18842
rect 28690 18790 28720 18842
rect 1344 18756 28720 18790
rect 21310 18674 21362 18686
rect 5394 18622 5406 18674
rect 5458 18622 5470 18674
rect 13570 18622 13582 18674
rect 13634 18622 13646 18674
rect 21310 18610 21362 18622
rect 24110 18674 24162 18686
rect 24110 18610 24162 18622
rect 5966 18562 6018 18574
rect 20190 18562 20242 18574
rect 8418 18510 8430 18562
rect 8482 18510 8494 18562
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 23202 18510 23214 18562
rect 23266 18510 23278 18562
rect 28018 18510 28030 18562
rect 28082 18510 28094 18562
rect 5966 18498 6018 18510
rect 20190 18498 20242 18510
rect 2494 18450 2546 18462
rect 10670 18450 10722 18462
rect 14142 18450 14194 18462
rect 17502 18450 17554 18462
rect 2930 18398 2942 18450
rect 2994 18398 3006 18450
rect 11106 18398 11118 18450
rect 11170 18398 11182 18450
rect 14354 18398 14366 18450
rect 14418 18398 14430 18450
rect 16034 18398 16046 18450
rect 16098 18398 16110 18450
rect 17826 18398 17838 18450
rect 17890 18398 17902 18450
rect 24098 18398 24110 18450
rect 24162 18398 24174 18450
rect 2494 18386 2546 18398
rect 10670 18386 10722 18398
rect 14142 18386 14194 18398
rect 17502 18386 17554 18398
rect 1822 18338 1874 18350
rect 15374 18338 15426 18350
rect 7186 18286 7198 18338
rect 7250 18286 7262 18338
rect 1822 18274 1874 18286
rect 15374 18274 15426 18286
rect 16718 18338 16770 18350
rect 22194 18286 22206 18338
rect 22258 18286 22270 18338
rect 26674 18286 26686 18338
rect 26738 18286 26750 18338
rect 16718 18274 16770 18286
rect 20974 18226 21026 18238
rect 20974 18162 21026 18174
rect 1344 18058 28560 18092
rect 1344 18006 4616 18058
rect 4668 18006 4720 18058
rect 4772 18006 4824 18058
rect 4876 18006 11420 18058
rect 11472 18006 11524 18058
rect 11576 18006 11628 18058
rect 11680 18006 18224 18058
rect 18276 18006 18328 18058
rect 18380 18006 18432 18058
rect 18484 18006 25028 18058
rect 25080 18006 25132 18058
rect 25184 18006 25236 18058
rect 25288 18006 28560 18058
rect 1344 17972 28560 18006
rect 11790 17890 11842 17902
rect 11790 17826 11842 17838
rect 18510 17890 18562 17902
rect 18510 17826 18562 17838
rect 28254 17890 28306 17902
rect 28254 17826 28306 17838
rect 24222 17778 24274 17790
rect 19842 17726 19854 17778
rect 19906 17726 19918 17778
rect 20738 17726 20750 17778
rect 20802 17726 20814 17778
rect 22306 17726 22318 17778
rect 22370 17726 22382 17778
rect 24222 17714 24274 17726
rect 2270 17666 2322 17678
rect 2270 17602 2322 17614
rect 8094 17666 8146 17678
rect 15038 17666 15090 17678
rect 21422 17666 21474 17678
rect 8754 17614 8766 17666
rect 8818 17614 8830 17666
rect 15474 17614 15486 17666
rect 15538 17614 15550 17666
rect 18946 17614 18958 17666
rect 19010 17614 19022 17666
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 20514 17614 20526 17666
rect 20578 17614 20590 17666
rect 8094 17602 8146 17614
rect 15038 17602 15090 17614
rect 21422 17602 21474 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 24782 17666 24834 17678
rect 25218 17614 25230 17666
rect 25282 17614 25294 17666
rect 24782 17602 24834 17614
rect 7422 17554 7474 17566
rect 12350 17554 12402 17566
rect 12002 17502 12014 17554
rect 12066 17502 12078 17554
rect 7422 17490 7474 17502
rect 12350 17490 12402 17502
rect 17726 17554 17778 17566
rect 18722 17502 18734 17554
rect 18786 17502 18798 17554
rect 23538 17502 23550 17554
rect 23602 17502 23614 17554
rect 17726 17490 17778 17502
rect 1710 17442 1762 17454
rect 1710 17378 1762 17390
rect 7534 17442 7586 17454
rect 11218 17390 11230 17442
rect 11282 17390 11294 17442
rect 27570 17390 27582 17442
rect 27634 17390 27646 17442
rect 7534 17378 7586 17390
rect 1344 17274 28720 17308
rect 1344 17222 8018 17274
rect 8070 17222 8122 17274
rect 8174 17222 8226 17274
rect 8278 17222 14822 17274
rect 14874 17222 14926 17274
rect 14978 17222 15030 17274
rect 15082 17222 21626 17274
rect 21678 17222 21730 17274
rect 21782 17222 21834 17274
rect 21886 17222 28430 17274
rect 28482 17222 28534 17274
rect 28586 17222 28638 17274
rect 28690 17222 28720 17274
rect 1344 17188 28720 17222
rect 8318 17106 8370 17118
rect 7522 17054 7534 17106
rect 7586 17054 7598 17106
rect 8318 17042 8370 17054
rect 17838 17106 17890 17118
rect 25342 17106 25394 17118
rect 23426 17054 23438 17106
rect 23490 17054 23502 17106
rect 17838 17042 17890 17054
rect 25342 17042 25394 17054
rect 13358 16994 13410 17006
rect 2034 16942 2046 16994
rect 2098 16942 2110 16994
rect 13358 16930 13410 16942
rect 14142 16994 14194 17006
rect 16370 16942 16382 16994
rect 16434 16942 16446 16994
rect 19954 16942 19966 16994
rect 20018 16942 20030 16994
rect 24210 16942 24222 16994
rect 24274 16942 24286 16994
rect 27234 16942 27246 16994
rect 27298 16942 27310 16994
rect 14142 16930 14194 16942
rect 4622 16882 4674 16894
rect 10670 16882 10722 16894
rect 18286 16882 18338 16894
rect 5282 16830 5294 16882
rect 5346 16830 5358 16882
rect 9762 16830 9774 16882
rect 9826 16830 9838 16882
rect 11106 16830 11118 16882
rect 11170 16830 11182 16882
rect 4622 16818 4674 16830
rect 10670 16818 10722 16830
rect 18286 16818 18338 16830
rect 20526 16882 20578 16894
rect 25790 16882 25842 16894
rect 20850 16830 20862 16882
rect 20914 16830 20926 16882
rect 24434 16830 24446 16882
rect 24498 16830 24510 16882
rect 20526 16818 20578 16830
rect 25790 16818 25842 16830
rect 28142 16882 28194 16894
rect 28142 16818 28194 16830
rect 3154 16718 3166 16770
rect 3218 16718 3230 16770
rect 9538 16718 9550 16770
rect 9602 16718 9614 16770
rect 15362 16718 15374 16770
rect 15426 16718 15438 16770
rect 18610 16718 18622 16770
rect 18674 16718 18686 16770
rect 26226 16718 26238 16770
rect 26290 16718 26302 16770
rect 23998 16658 24050 16670
rect 23998 16594 24050 16606
rect 1344 16490 28560 16524
rect 1344 16438 4616 16490
rect 4668 16438 4720 16490
rect 4772 16438 4824 16490
rect 4876 16438 11420 16490
rect 11472 16438 11524 16490
rect 11576 16438 11628 16490
rect 11680 16438 18224 16490
rect 18276 16438 18328 16490
rect 18380 16438 18432 16490
rect 18484 16438 25028 16490
rect 25080 16438 25132 16490
rect 25184 16438 25236 16490
rect 25288 16438 28560 16490
rect 1344 16404 28560 16438
rect 10334 16322 10386 16334
rect 10334 16258 10386 16270
rect 5618 16158 5630 16210
rect 5682 16158 5694 16210
rect 12898 16158 12910 16210
rect 12962 16158 12974 16210
rect 18274 16158 18286 16210
rect 18338 16158 18350 16210
rect 27682 16158 27694 16210
rect 27746 16158 27758 16210
rect 6638 16098 6690 16110
rect 7298 16046 7310 16098
rect 7362 16046 7374 16098
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 14018 16046 14030 16098
rect 14082 16046 14094 16098
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 22082 16046 22094 16098
rect 22146 16046 22158 16098
rect 6638 16034 6690 16046
rect 5070 15986 5122 15998
rect 4722 15934 4734 15986
rect 4786 15934 4798 15986
rect 5070 15922 5122 15934
rect 5966 15986 6018 15998
rect 5966 15922 6018 15934
rect 9550 15986 9602 15998
rect 9550 15922 9602 15934
rect 12350 15986 12402 15998
rect 12350 15922 12402 15934
rect 12574 15986 12626 15998
rect 12574 15922 12626 15934
rect 17054 15986 17106 15998
rect 19282 15934 19294 15986
rect 19346 15934 19358 15986
rect 24882 15934 24894 15986
rect 24946 15934 24958 15986
rect 17054 15922 17106 15934
rect 20302 15874 20354 15886
rect 16482 15822 16494 15874
rect 16546 15822 16558 15874
rect 20302 15810 20354 15822
rect 28142 15874 28194 15886
rect 28142 15810 28194 15822
rect 1344 15706 28720 15740
rect 1344 15654 8018 15706
rect 8070 15654 8122 15706
rect 8174 15654 8226 15706
rect 8278 15654 14822 15706
rect 14874 15654 14926 15706
rect 14978 15654 15030 15706
rect 15082 15654 21626 15706
rect 21678 15654 21730 15706
rect 21782 15654 21834 15706
rect 21886 15654 28430 15706
rect 28482 15654 28534 15706
rect 28586 15654 28638 15706
rect 28690 15654 28720 15706
rect 1344 15620 28720 15654
rect 2046 15538 2098 15550
rect 15710 15538 15762 15550
rect 21758 15538 21810 15550
rect 2818 15486 2830 15538
rect 2882 15486 2894 15538
rect 20850 15486 20862 15538
rect 20914 15486 20926 15538
rect 2046 15474 2098 15486
rect 15710 15474 15762 15486
rect 21758 15474 21810 15486
rect 27134 15538 27186 15550
rect 27134 15474 27186 15486
rect 6738 15374 6750 15426
rect 6802 15374 6814 15426
rect 12786 15374 12798 15426
rect 12850 15374 12862 15426
rect 15138 15374 15150 15426
rect 15202 15374 15214 15426
rect 23650 15374 23662 15426
rect 23714 15374 23726 15426
rect 25330 15374 25342 15426
rect 25394 15374 25406 15426
rect 5518 15314 5570 15326
rect 21422 15314 21474 15326
rect 5058 15262 5070 15314
rect 5122 15262 5134 15314
rect 14466 15262 14478 15314
rect 14530 15262 14542 15314
rect 17826 15262 17838 15314
rect 17890 15262 17902 15314
rect 18386 15262 18398 15314
rect 18450 15262 18462 15314
rect 5518 15250 5570 15262
rect 21422 15250 21474 15262
rect 22318 15202 22370 15214
rect 27582 15202 27634 15214
rect 7970 15150 7982 15202
rect 8034 15150 8046 15202
rect 22642 15150 22654 15202
rect 22706 15150 22718 15202
rect 26450 15150 26462 15202
rect 26514 15150 26526 15202
rect 22318 15138 22370 15150
rect 27582 15138 27634 15150
rect 28030 15202 28082 15214
rect 28030 15138 28082 15150
rect 1344 14922 28560 14956
rect 1344 14870 4616 14922
rect 4668 14870 4720 14922
rect 4772 14870 4824 14922
rect 4876 14870 11420 14922
rect 11472 14870 11524 14922
rect 11576 14870 11628 14922
rect 11680 14870 18224 14922
rect 18276 14870 18328 14922
rect 18380 14870 18432 14922
rect 18484 14870 25028 14922
rect 25080 14870 25132 14922
rect 25184 14870 25236 14922
rect 25288 14870 28560 14922
rect 1344 14836 28560 14870
rect 19294 14754 19346 14766
rect 19294 14690 19346 14702
rect 23214 14754 23266 14766
rect 23214 14690 23266 14702
rect 20190 14642 20242 14654
rect 27134 14642 27186 14654
rect 4050 14590 4062 14642
rect 4114 14590 4126 14642
rect 12562 14590 12574 14642
rect 12626 14590 12638 14642
rect 21634 14590 21646 14642
rect 21698 14590 21710 14642
rect 20190 14578 20242 14590
rect 27134 14578 27186 14590
rect 10334 14530 10386 14542
rect 15822 14530 15874 14542
rect 26686 14530 26738 14542
rect 9650 14478 9662 14530
rect 9714 14478 9726 14530
rect 12786 14478 12798 14530
rect 12850 14478 12862 14530
rect 14690 14478 14702 14530
rect 14754 14478 14766 14530
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 26338 14478 26350 14530
rect 26402 14478 26414 14530
rect 28018 14478 28030 14530
rect 28082 14478 28094 14530
rect 10334 14466 10386 14478
rect 15822 14466 15874 14478
rect 26686 14466 26738 14478
rect 6414 14418 6466 14430
rect 3042 14366 3054 14418
rect 3106 14366 3118 14418
rect 6066 14366 6078 14418
rect 6130 14366 6142 14418
rect 6414 14354 6466 14366
rect 11902 14418 11954 14430
rect 22654 14418 22706 14430
rect 13906 14366 13918 14418
rect 13970 14366 13982 14418
rect 22978 14366 22990 14418
rect 23042 14366 23054 14418
rect 27794 14366 27806 14418
rect 27858 14366 27870 14418
rect 11902 14354 11954 14366
rect 22654 14354 22706 14366
rect 6638 14306 6690 14318
rect 12014 14306 12066 14318
rect 19742 14306 19794 14318
rect 7410 14254 7422 14306
rect 7474 14254 7486 14306
rect 18722 14254 18734 14306
rect 18786 14254 18798 14306
rect 6638 14242 6690 14254
rect 12014 14242 12066 14254
rect 19742 14242 19794 14254
rect 20750 14306 20802 14318
rect 27246 14306 27298 14318
rect 23986 14254 23998 14306
rect 24050 14254 24062 14306
rect 20750 14242 20802 14254
rect 27246 14242 27298 14254
rect 1344 14138 28720 14172
rect 1344 14086 8018 14138
rect 8070 14086 8122 14138
rect 8174 14086 8226 14138
rect 8278 14086 14822 14138
rect 14874 14086 14926 14138
rect 14978 14086 15030 14138
rect 15082 14086 21626 14138
rect 21678 14086 21730 14138
rect 21782 14086 21834 14138
rect 21886 14086 28430 14138
rect 28482 14086 28534 14138
rect 28586 14086 28638 14138
rect 28690 14086 28720 14138
rect 1344 14052 28720 14086
rect 4174 13970 4226 13982
rect 15150 13970 15202 13982
rect 23774 13970 23826 13982
rect 4946 13918 4958 13970
rect 5010 13918 5022 13970
rect 11778 13918 11790 13970
rect 11842 13918 11854 13970
rect 22978 13918 22990 13970
rect 23042 13918 23054 13970
rect 4174 13906 4226 13918
rect 15150 13906 15202 13918
rect 23774 13906 23826 13918
rect 25902 13970 25954 13982
rect 25902 13906 25954 13918
rect 8990 13858 9042 13870
rect 8642 13806 8654 13858
rect 8706 13806 8718 13858
rect 19394 13806 19406 13858
rect 19458 13806 19470 13858
rect 27458 13806 27470 13858
rect 27522 13806 27534 13858
rect 8990 13794 9042 13806
rect 7870 13746 7922 13758
rect 14814 13746 14866 13758
rect 7298 13694 7310 13746
rect 7362 13694 7374 13746
rect 14242 13694 14254 13746
rect 14306 13694 14318 13746
rect 7870 13682 7922 13694
rect 14814 13682 14866 13694
rect 20302 13746 20354 13758
rect 20738 13694 20750 13746
rect 20802 13694 20814 13746
rect 20302 13682 20354 13694
rect 24222 13634 24274 13646
rect 18386 13582 18398 13634
rect 18450 13582 18462 13634
rect 26226 13582 26238 13634
rect 26290 13582 26302 13634
rect 24222 13570 24274 13582
rect 11118 13522 11170 13534
rect 11118 13458 11170 13470
rect 1344 13354 28560 13388
rect 1344 13302 4616 13354
rect 4668 13302 4720 13354
rect 4772 13302 4824 13354
rect 4876 13302 11420 13354
rect 11472 13302 11524 13354
rect 11576 13302 11628 13354
rect 11680 13302 18224 13354
rect 18276 13302 18328 13354
rect 18380 13302 18432 13354
rect 18484 13302 25028 13354
rect 25080 13302 25132 13354
rect 25184 13302 25236 13354
rect 25288 13302 28560 13354
rect 1344 13268 28560 13302
rect 12798 13186 12850 13198
rect 12798 13122 12850 13134
rect 14926 13074 14978 13086
rect 4050 13022 4062 13074
rect 4114 13022 4126 13074
rect 7410 13022 7422 13074
rect 7474 13022 7486 13074
rect 14926 13010 14978 13022
rect 21422 13074 21474 13086
rect 21422 13010 21474 13022
rect 27358 13074 27410 13086
rect 27358 13010 27410 13022
rect 28142 13074 28194 13086
rect 28142 13010 28194 13022
rect 9326 12962 9378 12974
rect 22766 12962 22818 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 5842 12910 5854 12962
rect 5906 12910 5918 12962
rect 9650 12910 9662 12962
rect 9714 12910 9726 12962
rect 15138 12910 15150 12962
rect 15202 12910 15214 12962
rect 23426 12910 23438 12962
rect 23490 12910 23502 12962
rect 26674 12910 26686 12962
rect 26738 12910 26750 12962
rect 26898 12910 26910 12962
rect 26962 12910 26974 12962
rect 9326 12898 9378 12910
rect 22766 12898 22818 12910
rect 12014 12850 12066 12862
rect 3042 12798 3054 12850
rect 3106 12798 3118 12850
rect 6066 12798 6078 12850
rect 6130 12798 6142 12850
rect 8754 12798 8766 12850
rect 8818 12798 8830 12850
rect 20066 12798 20078 12850
rect 20130 12798 20142 12850
rect 12014 12786 12066 12798
rect 2046 12738 2098 12750
rect 2046 12674 2098 12686
rect 6526 12738 6578 12750
rect 26462 12738 26514 12750
rect 25890 12686 25902 12738
rect 25954 12686 25966 12738
rect 6526 12674 6578 12686
rect 26462 12674 26514 12686
rect 27470 12738 27522 12750
rect 27470 12674 27522 12686
rect 1344 12570 28720 12604
rect 1344 12518 8018 12570
rect 8070 12518 8122 12570
rect 8174 12518 8226 12570
rect 8278 12518 14822 12570
rect 14874 12518 14926 12570
rect 14978 12518 15030 12570
rect 15082 12518 21626 12570
rect 21678 12518 21730 12570
rect 21782 12518 21834 12570
rect 21886 12518 28430 12570
rect 28482 12518 28534 12570
rect 28586 12518 28638 12570
rect 28690 12518 28720 12570
rect 1344 12484 28720 12518
rect 7074 12350 7086 12402
rect 7138 12350 7150 12402
rect 8654 12290 8706 12302
rect 8654 12226 8706 12238
rect 18062 12290 18114 12302
rect 18062 12226 18114 12238
rect 23998 12290 24050 12302
rect 27234 12238 27246 12290
rect 27298 12238 27310 12290
rect 23998 12226 24050 12238
rect 1822 12178 1874 12190
rect 1822 12114 1874 12126
rect 3390 12178 3442 12190
rect 4398 12178 4450 12190
rect 20974 12178 21026 12190
rect 3714 12126 3726 12178
rect 3778 12126 3790 12178
rect 4722 12126 4734 12178
rect 4786 12126 4798 12178
rect 14466 12126 14478 12178
rect 14530 12126 14542 12178
rect 20402 12126 20414 12178
rect 20466 12126 20478 12178
rect 3390 12114 3442 12126
rect 4398 12114 4450 12126
rect 20974 12114 21026 12126
rect 21086 12178 21138 12190
rect 21634 12126 21646 12178
rect 21698 12126 21710 12178
rect 21086 12114 21138 12126
rect 25342 12066 25394 12078
rect 3938 12014 3950 12066
rect 4002 12014 4014 12066
rect 8866 12014 8878 12066
rect 8930 12014 8942 12066
rect 10098 12014 10110 12066
rect 10162 12014 10174 12066
rect 25342 12002 25394 12014
rect 25902 12066 25954 12078
rect 26226 12014 26238 12066
rect 26290 12014 26302 12066
rect 25902 12002 25954 12014
rect 7870 11954 7922 11966
rect 7870 11890 7922 11902
rect 17278 11954 17330 11966
rect 17278 11890 17330 11902
rect 24782 11954 24834 11966
rect 24782 11890 24834 11902
rect 1344 11786 28560 11820
rect 1344 11734 4616 11786
rect 4668 11734 4720 11786
rect 4772 11734 4824 11786
rect 4876 11734 11420 11786
rect 11472 11734 11524 11786
rect 11576 11734 11628 11786
rect 11680 11734 18224 11786
rect 18276 11734 18328 11786
rect 18380 11734 18432 11786
rect 18484 11734 25028 11786
rect 25080 11734 25132 11786
rect 25184 11734 25236 11786
rect 25288 11734 28560 11786
rect 1344 11700 28560 11734
rect 7198 11618 7250 11630
rect 7198 11554 7250 11566
rect 3826 11454 3838 11506
rect 3890 11454 3902 11506
rect 23538 11454 23550 11506
rect 23602 11454 23614 11506
rect 27010 11454 27022 11506
rect 27074 11454 27086 11506
rect 10670 11394 10722 11406
rect 10322 11342 10334 11394
rect 10386 11342 10398 11394
rect 10670 11330 10722 11342
rect 15710 11394 15762 11406
rect 19182 11394 19234 11406
rect 16146 11342 16158 11394
rect 16210 11342 16222 11394
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 15710 11330 15762 11342
rect 19182 11330 19234 11342
rect 7982 11282 8034 11294
rect 11454 11282 11506 11294
rect 12238 11282 12290 11294
rect 19742 11282 19794 11294
rect 4946 11230 4958 11282
rect 5010 11230 5022 11282
rect 11106 11230 11118 11282
rect 11170 11230 11182 11282
rect 11890 11230 11902 11282
rect 11954 11230 11966 11282
rect 19394 11230 19406 11282
rect 19458 11230 19470 11282
rect 7982 11218 8034 11230
rect 11454 11218 11506 11230
rect 12238 11218 12290 11230
rect 19742 11218 19794 11230
rect 20078 11282 20130 11294
rect 20078 11218 20130 11230
rect 27246 11282 27298 11294
rect 27246 11218 27298 11230
rect 27582 11282 27634 11294
rect 27582 11218 27634 11230
rect 12686 11170 12738 11182
rect 20190 11170 20242 11182
rect 18610 11118 18622 11170
rect 18674 11118 18686 11170
rect 12686 11106 12738 11118
rect 20190 11106 20242 11118
rect 27694 11170 27746 11182
rect 27694 11106 27746 11118
rect 1344 11002 28720 11036
rect 1344 10950 8018 11002
rect 8070 10950 8122 11002
rect 8174 10950 8226 11002
rect 8278 10950 14822 11002
rect 14874 10950 14926 11002
rect 14978 10950 15030 11002
rect 15082 10950 21626 11002
rect 21678 10950 21730 11002
rect 21782 10950 21834 11002
rect 21886 10950 28430 11002
rect 28482 10950 28534 11002
rect 28586 10950 28638 11002
rect 28690 10950 28720 11002
rect 1344 10916 28720 10950
rect 5294 10834 5346 10846
rect 11678 10834 11730 10846
rect 23998 10834 24050 10846
rect 4498 10782 4510 10834
rect 4562 10782 4574 10834
rect 8306 10782 8318 10834
rect 8370 10782 8382 10834
rect 15586 10782 15598 10834
rect 15650 10782 15662 10834
rect 23090 10782 23102 10834
rect 23154 10782 23166 10834
rect 5294 10770 5346 10782
rect 11678 10770 11730 10782
rect 23998 10770 24050 10782
rect 28142 10834 28194 10846
rect 28142 10770 28194 10782
rect 9874 10670 9886 10722
rect 9938 10670 9950 10722
rect 16370 10670 16382 10722
rect 16434 10670 16446 10722
rect 27570 10670 27582 10722
rect 27634 10670 27646 10722
rect 1822 10610 1874 10622
rect 5630 10610 5682 10622
rect 12462 10610 12514 10622
rect 19966 10610 20018 10622
rect 2146 10558 2158 10610
rect 2210 10558 2222 10610
rect 6066 10558 6078 10610
rect 6130 10558 6142 10610
rect 13010 10558 13022 10610
rect 13074 10558 13086 10610
rect 20626 10558 20638 10610
rect 20690 10558 20702 10610
rect 24546 10558 24558 10610
rect 24610 10558 24622 10610
rect 1822 10546 1874 10558
rect 5630 10546 5682 10558
rect 12462 10546 12514 10558
rect 19966 10546 20018 10558
rect 16718 10498 16770 10510
rect 11218 10446 11230 10498
rect 11282 10446 11294 10498
rect 16718 10434 16770 10446
rect 17502 10498 17554 10510
rect 17502 10434 17554 10446
rect 19294 10498 19346 10510
rect 19294 10434 19346 10446
rect 19742 10498 19794 10510
rect 24322 10446 24334 10498
rect 24386 10446 24398 10498
rect 26226 10446 26238 10498
rect 26290 10446 26302 10498
rect 19742 10434 19794 10446
rect 9102 10386 9154 10398
rect 9102 10322 9154 10334
rect 16158 10386 16210 10398
rect 16158 10322 16210 10334
rect 23662 10386 23714 10398
rect 23662 10322 23714 10334
rect 1344 10218 28560 10252
rect 1344 10166 4616 10218
rect 4668 10166 4720 10218
rect 4772 10166 4824 10218
rect 4876 10166 11420 10218
rect 11472 10166 11524 10218
rect 11576 10166 11628 10218
rect 11680 10166 18224 10218
rect 18276 10166 18328 10218
rect 18380 10166 18432 10218
rect 18484 10166 25028 10218
rect 25080 10166 25132 10218
rect 25184 10166 25236 10218
rect 25288 10166 28560 10218
rect 1344 10132 28560 10166
rect 9326 10050 9378 10062
rect 9326 9986 9378 9998
rect 28254 10050 28306 10062
rect 28254 9986 28306 9998
rect 19742 9938 19794 9950
rect 23538 9886 23550 9938
rect 23602 9886 23614 9938
rect 19742 9874 19794 9886
rect 12798 9826 12850 9838
rect 5618 9774 5630 9826
rect 5682 9774 5694 9826
rect 6178 9774 6190 9826
rect 6242 9774 6254 9826
rect 12338 9774 12350 9826
rect 12402 9774 12414 9826
rect 12798 9762 12850 9774
rect 15710 9826 15762 9838
rect 24782 9826 24834 9838
rect 16146 9774 16158 9826
rect 16210 9774 16222 9826
rect 20290 9774 20302 9826
rect 20354 9774 20366 9826
rect 21522 9774 21534 9826
rect 21586 9774 21598 9826
rect 25218 9774 25230 9826
rect 25282 9774 25294 9826
rect 15710 9762 15762 9774
rect 24782 9762 24834 9774
rect 4622 9714 4674 9726
rect 4274 9662 4286 9714
rect 4338 9662 4350 9714
rect 4622 9650 4674 9662
rect 10110 9714 10162 9726
rect 27470 9714 27522 9726
rect 19394 9662 19406 9714
rect 19458 9662 19470 9714
rect 20514 9662 20526 9714
rect 20578 9662 20590 9714
rect 10110 9650 10162 9662
rect 27470 9650 27522 9662
rect 5070 9602 5122 9614
rect 9214 9602 9266 9614
rect 19182 9602 19234 9614
rect 8530 9550 8542 9602
rect 8594 9550 8606 9602
rect 18610 9550 18622 9602
rect 18674 9550 18686 9602
rect 5070 9538 5122 9550
rect 9214 9538 9266 9550
rect 19182 9538 19234 9550
rect 1344 9434 28720 9468
rect 1344 9382 8018 9434
rect 8070 9382 8122 9434
rect 8174 9382 8226 9434
rect 8278 9382 14822 9434
rect 14874 9382 14926 9434
rect 14978 9382 15030 9434
rect 15082 9382 21626 9434
rect 21678 9382 21730 9434
rect 21782 9382 21834 9434
rect 21886 9382 28430 9434
rect 28482 9382 28534 9434
rect 28586 9382 28638 9434
rect 28690 9382 28720 9434
rect 1344 9348 28720 9382
rect 21982 9266 22034 9278
rect 5394 9214 5406 9266
rect 5458 9214 5470 9266
rect 20514 9214 20526 9266
rect 20578 9214 20590 9266
rect 21982 9202 22034 9214
rect 28142 9266 28194 9278
rect 28142 9202 28194 9214
rect 15598 9154 15650 9166
rect 8866 9102 8878 9154
rect 8930 9102 8942 9154
rect 10098 9102 10110 9154
rect 10162 9102 10174 9154
rect 23538 9102 23550 9154
rect 23602 9102 23614 9154
rect 24210 9102 24222 9154
rect 24274 9102 24286 9154
rect 27458 9102 27470 9154
rect 27522 9102 27534 9154
rect 15598 9090 15650 9102
rect 2494 9042 2546 9054
rect 17502 9042 17554 9054
rect 2818 8990 2830 9042
rect 2882 8990 2894 9042
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 13234 8990 13246 9042
rect 13298 8990 13310 9042
rect 18162 8990 18174 9042
rect 18226 8990 18238 9042
rect 24434 8990 24446 9042
rect 24498 8990 24510 9042
rect 2494 8978 2546 8990
rect 17502 8978 17554 8990
rect 21534 8930 21586 8942
rect 7522 8878 7534 8930
rect 7586 8878 7598 8930
rect 11442 8878 11454 8930
rect 11506 8878 11518 8930
rect 22418 8878 22430 8930
rect 22482 8878 22494 8930
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 21534 8866 21586 8878
rect 5966 8818 6018 8830
rect 5966 8754 6018 8766
rect 16382 8818 16434 8830
rect 16382 8754 16434 8766
rect 21198 8818 21250 8830
rect 21198 8754 21250 8766
rect 1344 8650 28560 8684
rect 1344 8598 4616 8650
rect 4668 8598 4720 8650
rect 4772 8598 4824 8650
rect 4876 8598 11420 8650
rect 11472 8598 11524 8650
rect 11576 8598 11628 8650
rect 11680 8598 18224 8650
rect 18276 8598 18328 8650
rect 18380 8598 18432 8650
rect 18484 8598 25028 8650
rect 25080 8598 25132 8650
rect 25184 8598 25236 8650
rect 25288 8598 28560 8650
rect 1344 8564 28560 8598
rect 6078 8370 6130 8382
rect 9326 8370 9378 8382
rect 28254 8370 28306 8382
rect 3602 8318 3614 8370
rect 3666 8318 3678 8370
rect 5730 8318 5742 8370
rect 5794 8318 5806 8370
rect 7410 8318 7422 8370
rect 7474 8318 7486 8370
rect 15138 8318 15150 8370
rect 15202 8318 15214 8370
rect 17602 8318 17614 8370
rect 17666 8318 17678 8370
rect 22306 8318 22318 8370
rect 22370 8318 22382 8370
rect 6078 8306 6130 8318
rect 9326 8306 9378 8318
rect 28254 8306 28306 8318
rect 12798 8258 12850 8270
rect 24558 8258 24610 8270
rect 12450 8206 12462 8258
rect 12514 8206 12526 8258
rect 14130 8206 14142 8258
rect 14194 8206 14206 8258
rect 25218 8206 25230 8258
rect 25282 8206 25294 8258
rect 12798 8194 12850 8206
rect 24558 8194 24610 8206
rect 2482 8094 2494 8146
rect 2546 8094 2558 8146
rect 8642 8094 8654 8146
rect 8706 8094 8718 8146
rect 18610 8094 18622 8146
rect 18674 8094 18686 8146
rect 23538 8094 23550 8146
rect 23602 8094 23614 8146
rect 6526 8034 6578 8046
rect 16830 8034 16882 8046
rect 10098 7982 10110 8034
rect 10162 7982 10174 8034
rect 27682 7982 27694 8034
rect 27746 7982 27758 8034
rect 6526 7970 6578 7982
rect 16830 7970 16882 7982
rect 1344 7866 28720 7900
rect 1344 7814 8018 7866
rect 8070 7814 8122 7866
rect 8174 7814 8226 7866
rect 8278 7814 14822 7866
rect 14874 7814 14926 7866
rect 14978 7814 15030 7866
rect 15082 7814 21626 7866
rect 21678 7814 21730 7866
rect 21782 7814 21834 7866
rect 21886 7814 28430 7866
rect 28482 7814 28534 7866
rect 28586 7814 28638 7866
rect 28690 7814 28720 7866
rect 1344 7780 28720 7814
rect 1598 7698 1650 7710
rect 25342 7698 25394 7710
rect 2370 7646 2382 7698
rect 2434 7646 2446 7698
rect 21858 7646 21870 7698
rect 21922 7646 21934 7698
rect 1598 7634 1650 7646
rect 25342 7634 25394 7646
rect 28142 7586 28194 7598
rect 7186 7534 7198 7586
rect 7250 7534 7262 7586
rect 9762 7534 9774 7586
rect 9826 7534 9838 7586
rect 12450 7534 12462 7586
rect 12514 7534 12526 7586
rect 16258 7534 16270 7586
rect 16322 7534 16334 7586
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 28142 7522 28194 7534
rect 5294 7474 5346 7486
rect 24558 7474 24610 7486
rect 4722 7422 4734 7474
rect 4786 7422 4798 7474
rect 12674 7422 12686 7474
rect 12738 7422 12750 7474
rect 24210 7422 24222 7474
rect 24274 7422 24286 7474
rect 5294 7410 5346 7422
rect 24558 7410 24610 7422
rect 13246 7362 13298 7374
rect 6178 7310 6190 7362
rect 6242 7310 6254 7362
rect 11106 7310 11118 7362
rect 11170 7310 11182 7362
rect 14914 7310 14926 7362
rect 14978 7310 14990 7362
rect 26226 7310 26238 7362
rect 26290 7310 26302 7362
rect 13246 7298 13298 7310
rect 21086 7250 21138 7262
rect 21086 7186 21138 7198
rect 1344 7082 28560 7116
rect 1344 7030 4616 7082
rect 4668 7030 4720 7082
rect 4772 7030 4824 7082
rect 4876 7030 11420 7082
rect 11472 7030 11524 7082
rect 11576 7030 11628 7082
rect 11680 7030 18224 7082
rect 18276 7030 18328 7082
rect 18380 7030 18432 7082
rect 18484 7030 25028 7082
rect 25080 7030 25132 7082
rect 25184 7030 25236 7082
rect 25288 7030 28560 7082
rect 1344 6996 28560 7030
rect 14466 6750 14478 6802
rect 14530 6750 14542 6802
rect 8654 6690 8706 6702
rect 7970 6638 7982 6690
rect 8034 6638 8046 6690
rect 8194 6638 8206 6690
rect 8258 6638 8270 6690
rect 8654 6626 8706 6638
rect 23998 6690 24050 6702
rect 27470 6690 27522 6702
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 23998 6626 24050 6638
rect 27470 6626 27522 6638
rect 27694 6690 27746 6702
rect 27694 6626 27746 6638
rect 21646 6578 21698 6590
rect 15810 6526 15822 6578
rect 15874 6526 15886 6578
rect 21646 6514 21698 6526
rect 21982 6578 22034 6590
rect 21982 6514 22034 6526
rect 22318 6466 22370 6478
rect 22318 6402 22370 6414
rect 23102 6466 23154 6478
rect 27806 6466 27858 6478
rect 26786 6414 26798 6466
rect 26850 6414 26862 6466
rect 23102 6402 23154 6414
rect 27806 6402 27858 6414
rect 1344 6298 28720 6332
rect 1344 6246 8018 6298
rect 8070 6246 8122 6298
rect 8174 6246 8226 6298
rect 8278 6246 14822 6298
rect 14874 6246 14926 6298
rect 14978 6246 15030 6298
rect 15082 6246 21626 6298
rect 21678 6246 21730 6298
rect 21782 6246 21834 6298
rect 21886 6246 28430 6298
rect 28482 6246 28534 6298
rect 28586 6246 28638 6298
rect 28690 6246 28720 6298
rect 1344 6212 28720 6246
rect 14814 6130 14866 6142
rect 14814 6066 14866 6078
rect 26350 6130 26402 6142
rect 26350 6066 26402 6078
rect 13806 6018 13858 6030
rect 13806 5954 13858 5966
rect 15150 6018 15202 6030
rect 20862 6018 20914 6030
rect 24670 6018 24722 6030
rect 15474 5966 15486 6018
rect 15538 5966 15550 6018
rect 22530 5966 22542 6018
rect 22594 5966 22606 6018
rect 27682 5966 27694 6018
rect 27746 5966 27758 6018
rect 15150 5954 15202 5966
rect 20862 5954 20914 5966
rect 24670 5954 24722 5966
rect 13470 5906 13522 5918
rect 13470 5842 13522 5854
rect 21198 5906 21250 5918
rect 21198 5842 21250 5854
rect 20638 5794 20690 5806
rect 21522 5742 21534 5794
rect 21586 5742 21598 5794
rect 24322 5742 24334 5794
rect 24386 5742 24398 5794
rect 26674 5742 26686 5794
rect 26738 5742 26750 5794
rect 20638 5730 20690 5742
rect 1344 5514 28560 5548
rect 1344 5462 4616 5514
rect 4668 5462 4720 5514
rect 4772 5462 4824 5514
rect 4876 5462 11420 5514
rect 11472 5462 11524 5514
rect 11576 5462 11628 5514
rect 11680 5462 18224 5514
rect 18276 5462 18328 5514
rect 18380 5462 18432 5514
rect 18484 5462 25028 5514
rect 25080 5462 25132 5514
rect 25184 5462 25236 5514
rect 25288 5462 28560 5514
rect 1344 5428 28560 5462
rect 23314 5182 23326 5234
rect 23378 5182 23390 5234
rect 24558 5122 24610 5134
rect 19394 5070 19406 5122
rect 19458 5070 19470 5122
rect 25218 5070 25230 5122
rect 25282 5070 25294 5122
rect 24558 5058 24610 5070
rect 19630 5010 19682 5022
rect 19630 4946 19682 4958
rect 19966 5010 20018 5022
rect 22306 4958 22318 5010
rect 22370 4958 22382 5010
rect 19966 4946 20018 4958
rect 20302 4898 20354 4910
rect 20302 4834 20354 4846
rect 21534 4898 21586 4910
rect 28254 4898 28306 4910
rect 27682 4846 27694 4898
rect 27746 4846 27758 4898
rect 21534 4834 21586 4846
rect 28254 4834 28306 4846
rect 1344 4730 28720 4764
rect 1344 4678 8018 4730
rect 8070 4678 8122 4730
rect 8174 4678 8226 4730
rect 8278 4678 14822 4730
rect 14874 4678 14926 4730
rect 14978 4678 15030 4730
rect 15082 4678 21626 4730
rect 21678 4678 21730 4730
rect 21782 4678 21834 4730
rect 21886 4678 28430 4730
rect 28482 4678 28534 4730
rect 28586 4678 28638 4730
rect 28690 4678 28720 4730
rect 1344 4644 28720 4678
rect 24782 4562 24834 4574
rect 24210 4510 24222 4562
rect 24274 4510 24286 4562
rect 24782 4498 24834 4510
rect 25342 4562 25394 4574
rect 25342 4498 25394 4510
rect 25902 4562 25954 4574
rect 25902 4498 25954 4510
rect 14142 4450 14194 4462
rect 14142 4386 14194 4398
rect 14926 4450 14978 4462
rect 14926 4386 14978 4398
rect 15262 4450 15314 4462
rect 15262 4386 15314 4398
rect 18062 4450 18114 4462
rect 18062 4386 18114 4398
rect 19294 4450 19346 4462
rect 28142 4450 28194 4462
rect 27234 4398 27246 4450
rect 27298 4398 27310 4450
rect 19294 4386 19346 4398
rect 28142 4386 28194 4398
rect 21310 4338 21362 4350
rect 14690 4286 14702 4338
rect 14754 4286 14766 4338
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 20738 4286 20750 4338
rect 20802 4286 20814 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 21310 4274 21362 4286
rect 12798 4226 12850 4238
rect 12798 4162 12850 4174
rect 18734 4226 18786 4238
rect 18734 4162 18786 4174
rect 19742 4226 19794 4238
rect 20402 4174 20414 4226
rect 20466 4174 20478 4226
rect 26226 4174 26238 4226
rect 26290 4174 26302 4226
rect 19742 4162 19794 4174
rect 1344 3946 28560 3980
rect 1344 3894 4616 3946
rect 4668 3894 4720 3946
rect 4772 3894 4824 3946
rect 4876 3894 11420 3946
rect 11472 3894 11524 3946
rect 11576 3894 11628 3946
rect 11680 3894 18224 3946
rect 18276 3894 18328 3946
rect 18380 3894 18432 3946
rect 18484 3894 25028 3946
rect 25080 3894 25132 3946
rect 25184 3894 25236 3946
rect 25288 3894 28560 3946
rect 1344 3860 28560 3894
rect 15586 3614 15598 3666
rect 15650 3614 15662 3666
rect 21522 3614 21534 3666
rect 21586 3614 21598 3666
rect 23090 3614 23102 3666
rect 23154 3614 23166 3666
rect 26114 3614 26126 3666
rect 26178 3614 26190 3666
rect 15150 3554 15202 3566
rect 19406 3554 19458 3566
rect 22318 3554 22370 3566
rect 14242 3502 14254 3554
rect 14306 3502 14318 3554
rect 17154 3502 17166 3554
rect 17218 3502 17230 3554
rect 18498 3502 18510 3554
rect 18562 3502 18574 3554
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 15150 3490 15202 3502
rect 19406 3490 19458 3502
rect 22318 3490 22370 3502
rect 22654 3554 22706 3566
rect 22654 3490 22706 3502
rect 12238 3442 12290 3454
rect 12238 3378 12290 3390
rect 12574 3442 12626 3454
rect 12574 3378 12626 3390
rect 16494 3442 16546 3454
rect 16494 3378 16546 3390
rect 16942 3442 16994 3454
rect 16942 3378 16994 3390
rect 19070 3442 19122 3454
rect 19070 3378 19122 3390
rect 19854 3442 19906 3454
rect 19854 3378 19906 3390
rect 21086 3442 21138 3454
rect 27458 3390 27470 3442
rect 27522 3390 27534 3442
rect 21086 3378 21138 3390
rect 13134 3330 13186 3342
rect 13134 3266 13186 3278
rect 13582 3330 13634 3342
rect 13582 3266 13634 3278
rect 17614 3330 17666 3342
rect 17614 3266 17666 3278
rect 18734 3330 18786 3342
rect 18734 3266 18786 3278
rect 24782 3330 24834 3342
rect 24782 3266 24834 3278
rect 1344 3162 28720 3196
rect 1344 3110 8018 3162
rect 8070 3110 8122 3162
rect 8174 3110 8226 3162
rect 8278 3110 14822 3162
rect 14874 3110 14926 3162
rect 14978 3110 15030 3162
rect 15082 3110 21626 3162
rect 21678 3110 21730 3162
rect 21782 3110 21834 3162
rect 21886 3110 28430 3162
rect 28482 3110 28534 3162
rect 28586 3110 28638 3162
rect 28690 3110 28720 3162
rect 1344 3076 28720 3110
rect 16818 1710 16830 1762
rect 16882 1759 16894 1762
rect 17602 1759 17614 1762
rect 16882 1713 17614 1759
rect 16882 1710 16894 1713
rect 17602 1710 17614 1713
rect 17666 1710 17678 1762
<< via1 >>
rect 13470 27806 13522 27858
rect 14142 27806 14194 27858
rect 10110 26798 10162 26850
rect 11118 26798 11170 26850
rect 16830 26798 16882 26850
rect 17502 26798 17554 26850
rect 18846 26798 18898 26850
rect 19630 26798 19682 26850
rect 22206 26798 22258 26850
rect 22990 26798 23042 26850
rect 8018 26630 8070 26682
rect 8122 26630 8174 26682
rect 8226 26630 8278 26682
rect 14822 26630 14874 26682
rect 14926 26630 14978 26682
rect 15030 26630 15082 26682
rect 21626 26630 21678 26682
rect 21730 26630 21782 26682
rect 21834 26630 21886 26682
rect 28430 26630 28482 26682
rect 28534 26630 28586 26682
rect 28638 26630 28690 26682
rect 7646 26462 7698 26514
rect 8206 26462 8258 26514
rect 8766 26462 8818 26514
rect 11118 26462 11170 26514
rect 12014 26462 12066 26514
rect 13358 26462 13410 26514
rect 23886 26462 23938 26514
rect 25118 26462 25170 26514
rect 9662 26350 9714 26402
rect 12238 26350 12290 26402
rect 12574 26350 12626 26402
rect 15374 26350 15426 26402
rect 16046 26350 16098 26402
rect 26238 26350 26290 26402
rect 9886 26238 9938 26290
rect 10334 26238 10386 26290
rect 13694 26238 13746 26290
rect 15598 26238 15650 26290
rect 16270 26238 16322 26290
rect 17054 26238 17106 26290
rect 18734 26238 18786 26290
rect 20750 26238 20802 26290
rect 22318 26238 22370 26290
rect 26798 26238 26850 26290
rect 14142 26126 14194 26178
rect 17502 26126 17554 26178
rect 19070 26126 19122 26178
rect 21198 26126 21250 26178
rect 22766 26126 22818 26178
rect 27694 26126 27746 26178
rect 4616 25846 4668 25898
rect 4720 25846 4772 25898
rect 4824 25846 4876 25898
rect 11420 25846 11472 25898
rect 11524 25846 11576 25898
rect 11628 25846 11680 25898
rect 18224 25846 18276 25898
rect 18328 25846 18380 25898
rect 18432 25846 18484 25898
rect 25028 25846 25080 25898
rect 25132 25846 25184 25898
rect 25236 25846 25288 25898
rect 9438 25566 9490 25618
rect 10782 25566 10834 25618
rect 13918 25566 13970 25618
rect 15934 25566 15986 25618
rect 17166 25566 17218 25618
rect 18958 25566 19010 25618
rect 19630 25566 19682 25618
rect 11006 25454 11058 25506
rect 12574 25454 12626 25506
rect 16494 25454 16546 25506
rect 18510 25454 18562 25506
rect 20190 25454 20242 25506
rect 21422 25454 21474 25506
rect 22206 25454 22258 25506
rect 22990 25454 23042 25506
rect 27134 25454 27186 25506
rect 28142 25454 28194 25506
rect 11678 25342 11730 25394
rect 12910 25342 12962 25394
rect 15038 25342 15090 25394
rect 16718 25342 16770 25394
rect 20638 25342 20690 25394
rect 21646 25342 21698 25394
rect 22654 25342 22706 25394
rect 1710 25230 1762 25282
rect 11342 25230 11394 25282
rect 13470 25230 13522 25282
rect 19966 25230 20018 25282
rect 21982 25230 22034 25282
rect 27470 25230 27522 25282
rect 27806 25230 27858 25282
rect 8018 25062 8070 25114
rect 8122 25062 8174 25114
rect 8226 25062 8278 25114
rect 14822 25062 14874 25114
rect 14926 25062 14978 25114
rect 15030 25062 15082 25114
rect 21626 25062 21678 25114
rect 21730 25062 21782 25114
rect 21834 25062 21886 25114
rect 28430 25062 28482 25114
rect 28534 25062 28586 25114
rect 28638 25062 28690 25114
rect 13134 24894 13186 24946
rect 21758 24894 21810 24946
rect 22430 24894 22482 24946
rect 27022 24894 27074 24946
rect 12798 24782 12850 24834
rect 27358 24782 27410 24834
rect 28142 24782 28194 24834
rect 4616 24278 4668 24330
rect 4720 24278 4772 24330
rect 4824 24278 4876 24330
rect 11420 24278 11472 24330
rect 11524 24278 11576 24330
rect 11628 24278 11680 24330
rect 18224 24278 18276 24330
rect 18328 24278 18380 24330
rect 18432 24278 18484 24330
rect 25028 24278 25080 24330
rect 25132 24278 25184 24330
rect 25236 24278 25288 24330
rect 9326 23886 9378 23938
rect 18846 23886 18898 23938
rect 9550 23774 9602 23826
rect 19070 23774 19122 23826
rect 27694 23662 27746 23714
rect 28142 23662 28194 23714
rect 8018 23494 8070 23546
rect 8122 23494 8174 23546
rect 8226 23494 8278 23546
rect 14822 23494 14874 23546
rect 14926 23494 14978 23546
rect 15030 23494 15082 23546
rect 21626 23494 21678 23546
rect 21730 23494 21782 23546
rect 21834 23494 21886 23546
rect 28430 23494 28482 23546
rect 28534 23494 28586 23546
rect 28638 23494 28690 23546
rect 27134 23214 27186 23266
rect 27470 23214 27522 23266
rect 27806 23214 27858 23266
rect 28142 23102 28194 23154
rect 26910 22990 26962 23042
rect 4616 22710 4668 22762
rect 4720 22710 4772 22762
rect 4824 22710 4876 22762
rect 11420 22710 11472 22762
rect 11524 22710 11576 22762
rect 11628 22710 11680 22762
rect 18224 22710 18276 22762
rect 18328 22710 18380 22762
rect 18432 22710 18484 22762
rect 25028 22710 25080 22762
rect 25132 22710 25184 22762
rect 25236 22710 25288 22762
rect 27134 22318 27186 22370
rect 28030 22206 28082 22258
rect 8018 21926 8070 21978
rect 8122 21926 8174 21978
rect 8226 21926 8278 21978
rect 14822 21926 14874 21978
rect 14926 21926 14978 21978
rect 15030 21926 15082 21978
rect 21626 21926 21678 21978
rect 21730 21926 21782 21978
rect 21834 21926 21886 21978
rect 28430 21926 28482 21978
rect 28534 21926 28586 21978
rect 28638 21926 28690 21978
rect 15710 21758 15762 21810
rect 15374 21646 15426 21698
rect 16046 21646 16098 21698
rect 16382 21646 16434 21698
rect 27246 21646 27298 21698
rect 26014 21422 26066 21474
rect 26238 21422 26290 21474
rect 4616 21142 4668 21194
rect 4720 21142 4772 21194
rect 4824 21142 4876 21194
rect 11420 21142 11472 21194
rect 11524 21142 11576 21194
rect 11628 21142 11680 21194
rect 18224 21142 18276 21194
rect 18328 21142 18380 21194
rect 18432 21142 18484 21194
rect 25028 21142 25080 21194
rect 25132 21142 25184 21194
rect 25236 21142 25288 21194
rect 22990 20750 23042 20802
rect 23662 20750 23714 20802
rect 27806 20750 27858 20802
rect 26910 20638 26962 20690
rect 27246 20638 27298 20690
rect 27582 20638 27634 20690
rect 17278 20526 17330 20578
rect 26126 20526 26178 20578
rect 26686 20526 26738 20578
rect 8018 20358 8070 20410
rect 8122 20358 8174 20410
rect 8226 20358 8278 20410
rect 14822 20358 14874 20410
rect 14926 20358 14978 20410
rect 15030 20358 15082 20410
rect 21626 20358 21678 20410
rect 21730 20358 21782 20410
rect 21834 20358 21886 20410
rect 28430 20358 28482 20410
rect 28534 20358 28586 20410
rect 28638 20358 28690 20410
rect 22766 20190 22818 20242
rect 28142 20190 28194 20242
rect 11790 20078 11842 20130
rect 14030 20078 14082 20130
rect 16270 20078 16322 20130
rect 21646 20078 21698 20130
rect 13918 19966 13970 20018
rect 22430 20078 22482 20130
rect 27246 20078 27298 20130
rect 14254 19966 14306 20018
rect 18958 19966 19010 20018
rect 19406 19966 19458 20018
rect 25902 19966 25954 20018
rect 10670 19854 10722 19906
rect 13582 19854 13634 19906
rect 14366 19854 14418 19906
rect 15262 19854 15314 19906
rect 17614 19854 17666 19906
rect 17838 19854 17890 19906
rect 26238 19854 26290 19906
rect 4616 19574 4668 19626
rect 4720 19574 4772 19626
rect 4824 19574 4876 19626
rect 11420 19574 11472 19626
rect 11524 19574 11576 19626
rect 11628 19574 11680 19626
rect 18224 19574 18276 19626
rect 18328 19574 18380 19626
rect 18432 19574 18484 19626
rect 25028 19574 25080 19626
rect 25132 19574 25184 19626
rect 25236 19574 25288 19626
rect 24894 19406 24946 19458
rect 8654 19294 8706 19346
rect 11454 19294 11506 19346
rect 18286 19294 18338 19346
rect 26686 19294 26738 19346
rect 13470 19182 13522 19234
rect 14030 19182 14082 19234
rect 21422 19182 21474 19234
rect 21870 19182 21922 19234
rect 9662 19070 9714 19122
rect 12462 19070 12514 19122
rect 17054 19070 17106 19122
rect 19294 19070 19346 19122
rect 27694 19070 27746 19122
rect 16270 18958 16322 19010
rect 24110 18958 24162 19010
rect 25230 18958 25282 19010
rect 8018 18790 8070 18842
rect 8122 18790 8174 18842
rect 8226 18790 8278 18842
rect 14822 18790 14874 18842
rect 14926 18790 14978 18842
rect 15030 18790 15082 18842
rect 21626 18790 21678 18842
rect 21730 18790 21782 18842
rect 21834 18790 21886 18842
rect 28430 18790 28482 18842
rect 28534 18790 28586 18842
rect 28638 18790 28690 18842
rect 5406 18622 5458 18674
rect 13582 18622 13634 18674
rect 21310 18622 21362 18674
rect 24110 18622 24162 18674
rect 5966 18510 6018 18562
rect 8430 18510 8482 18562
rect 16270 18510 16322 18562
rect 20190 18510 20242 18562
rect 23214 18510 23266 18562
rect 28030 18510 28082 18562
rect 2494 18398 2546 18450
rect 2942 18398 2994 18450
rect 10670 18398 10722 18450
rect 11118 18398 11170 18450
rect 14142 18398 14194 18450
rect 14366 18398 14418 18450
rect 16046 18398 16098 18450
rect 17502 18398 17554 18450
rect 17838 18398 17890 18450
rect 24110 18398 24162 18450
rect 1822 18286 1874 18338
rect 7198 18286 7250 18338
rect 15374 18286 15426 18338
rect 16718 18286 16770 18338
rect 22206 18286 22258 18338
rect 26686 18286 26738 18338
rect 20974 18174 21026 18226
rect 4616 18006 4668 18058
rect 4720 18006 4772 18058
rect 4824 18006 4876 18058
rect 11420 18006 11472 18058
rect 11524 18006 11576 18058
rect 11628 18006 11680 18058
rect 18224 18006 18276 18058
rect 18328 18006 18380 18058
rect 18432 18006 18484 18058
rect 25028 18006 25080 18058
rect 25132 18006 25184 18058
rect 25236 18006 25288 18058
rect 11790 17838 11842 17890
rect 18510 17838 18562 17890
rect 28254 17838 28306 17890
rect 19854 17726 19906 17778
rect 20750 17726 20802 17778
rect 22318 17726 22370 17778
rect 24222 17726 24274 17778
rect 2270 17614 2322 17666
rect 8094 17614 8146 17666
rect 8766 17614 8818 17666
rect 15038 17614 15090 17666
rect 15486 17614 15538 17666
rect 18958 17614 19010 17666
rect 19630 17614 19682 17666
rect 20526 17614 20578 17666
rect 21422 17614 21474 17666
rect 21870 17614 21922 17666
rect 24782 17614 24834 17666
rect 25230 17614 25282 17666
rect 7422 17502 7474 17554
rect 12014 17502 12066 17554
rect 12350 17502 12402 17554
rect 17726 17502 17778 17554
rect 18734 17502 18786 17554
rect 23550 17502 23602 17554
rect 1710 17390 1762 17442
rect 7534 17390 7586 17442
rect 11230 17390 11282 17442
rect 27582 17390 27634 17442
rect 8018 17222 8070 17274
rect 8122 17222 8174 17274
rect 8226 17222 8278 17274
rect 14822 17222 14874 17274
rect 14926 17222 14978 17274
rect 15030 17222 15082 17274
rect 21626 17222 21678 17274
rect 21730 17222 21782 17274
rect 21834 17222 21886 17274
rect 28430 17222 28482 17274
rect 28534 17222 28586 17274
rect 28638 17222 28690 17274
rect 7534 17054 7586 17106
rect 8318 17054 8370 17106
rect 17838 17054 17890 17106
rect 23438 17054 23490 17106
rect 25342 17054 25394 17106
rect 2046 16942 2098 16994
rect 13358 16942 13410 16994
rect 14142 16942 14194 16994
rect 16382 16942 16434 16994
rect 19966 16942 20018 16994
rect 24222 16942 24274 16994
rect 27246 16942 27298 16994
rect 4622 16830 4674 16882
rect 5294 16830 5346 16882
rect 9774 16830 9826 16882
rect 10670 16830 10722 16882
rect 11118 16830 11170 16882
rect 18286 16830 18338 16882
rect 20526 16830 20578 16882
rect 20862 16830 20914 16882
rect 24446 16830 24498 16882
rect 25790 16830 25842 16882
rect 28142 16830 28194 16882
rect 3166 16718 3218 16770
rect 9550 16718 9602 16770
rect 15374 16718 15426 16770
rect 18622 16718 18674 16770
rect 26238 16718 26290 16770
rect 23998 16606 24050 16658
rect 4616 16438 4668 16490
rect 4720 16438 4772 16490
rect 4824 16438 4876 16490
rect 11420 16438 11472 16490
rect 11524 16438 11576 16490
rect 11628 16438 11680 16490
rect 18224 16438 18276 16490
rect 18328 16438 18380 16490
rect 18432 16438 18484 16490
rect 25028 16438 25080 16490
rect 25132 16438 25184 16490
rect 25236 16438 25288 16490
rect 10334 16270 10386 16322
rect 5630 16158 5682 16210
rect 12910 16158 12962 16210
rect 18286 16158 18338 16210
rect 27694 16158 27746 16210
rect 6638 16046 6690 16098
rect 7310 16046 7362 16098
rect 13470 16046 13522 16098
rect 14030 16046 14082 16098
rect 20302 16046 20354 16098
rect 22094 16046 22146 16098
rect 4734 15934 4786 15986
rect 5070 15934 5122 15986
rect 5966 15934 6018 15986
rect 9550 15934 9602 15986
rect 12350 15934 12402 15986
rect 12574 15934 12626 15986
rect 17054 15934 17106 15986
rect 19294 15934 19346 15986
rect 24894 15934 24946 15986
rect 16494 15822 16546 15874
rect 20302 15822 20354 15874
rect 28142 15822 28194 15874
rect 8018 15654 8070 15706
rect 8122 15654 8174 15706
rect 8226 15654 8278 15706
rect 14822 15654 14874 15706
rect 14926 15654 14978 15706
rect 15030 15654 15082 15706
rect 21626 15654 21678 15706
rect 21730 15654 21782 15706
rect 21834 15654 21886 15706
rect 28430 15654 28482 15706
rect 28534 15654 28586 15706
rect 28638 15654 28690 15706
rect 2046 15486 2098 15538
rect 2830 15486 2882 15538
rect 15710 15486 15762 15538
rect 20862 15486 20914 15538
rect 21758 15486 21810 15538
rect 27134 15486 27186 15538
rect 6750 15374 6802 15426
rect 12798 15374 12850 15426
rect 15150 15374 15202 15426
rect 23662 15374 23714 15426
rect 25342 15374 25394 15426
rect 5070 15262 5122 15314
rect 5518 15262 5570 15314
rect 14478 15262 14530 15314
rect 17838 15262 17890 15314
rect 18398 15262 18450 15314
rect 21422 15262 21474 15314
rect 7982 15150 8034 15202
rect 22318 15150 22370 15202
rect 22654 15150 22706 15202
rect 26462 15150 26514 15202
rect 27582 15150 27634 15202
rect 28030 15150 28082 15202
rect 4616 14870 4668 14922
rect 4720 14870 4772 14922
rect 4824 14870 4876 14922
rect 11420 14870 11472 14922
rect 11524 14870 11576 14922
rect 11628 14870 11680 14922
rect 18224 14870 18276 14922
rect 18328 14870 18380 14922
rect 18432 14870 18484 14922
rect 25028 14870 25080 14922
rect 25132 14870 25184 14922
rect 25236 14870 25288 14922
rect 19294 14702 19346 14754
rect 23214 14702 23266 14754
rect 4062 14590 4114 14642
rect 12574 14590 12626 14642
rect 20190 14590 20242 14642
rect 21646 14590 21698 14642
rect 27134 14590 27186 14642
rect 9662 14478 9714 14530
rect 10334 14478 10386 14530
rect 12798 14478 12850 14530
rect 14702 14478 14754 14530
rect 15822 14478 15874 14530
rect 16270 14478 16322 14530
rect 21870 14478 21922 14530
rect 26350 14478 26402 14530
rect 26686 14478 26738 14530
rect 28030 14478 28082 14530
rect 3054 14366 3106 14418
rect 6078 14366 6130 14418
rect 6414 14366 6466 14418
rect 11902 14366 11954 14418
rect 13918 14366 13970 14418
rect 22654 14366 22706 14418
rect 22990 14366 23042 14418
rect 27806 14366 27858 14418
rect 6638 14254 6690 14306
rect 7422 14254 7474 14306
rect 12014 14254 12066 14306
rect 18734 14254 18786 14306
rect 19742 14254 19794 14306
rect 20750 14254 20802 14306
rect 23998 14254 24050 14306
rect 27246 14254 27298 14306
rect 8018 14086 8070 14138
rect 8122 14086 8174 14138
rect 8226 14086 8278 14138
rect 14822 14086 14874 14138
rect 14926 14086 14978 14138
rect 15030 14086 15082 14138
rect 21626 14086 21678 14138
rect 21730 14086 21782 14138
rect 21834 14086 21886 14138
rect 28430 14086 28482 14138
rect 28534 14086 28586 14138
rect 28638 14086 28690 14138
rect 4174 13918 4226 13970
rect 4958 13918 5010 13970
rect 11790 13918 11842 13970
rect 15150 13918 15202 13970
rect 22990 13918 23042 13970
rect 23774 13918 23826 13970
rect 25902 13918 25954 13970
rect 8654 13806 8706 13858
rect 8990 13806 9042 13858
rect 19406 13806 19458 13858
rect 27470 13806 27522 13858
rect 7310 13694 7362 13746
rect 7870 13694 7922 13746
rect 14254 13694 14306 13746
rect 14814 13694 14866 13746
rect 20302 13694 20354 13746
rect 20750 13694 20802 13746
rect 18398 13582 18450 13634
rect 24222 13582 24274 13634
rect 26238 13582 26290 13634
rect 11118 13470 11170 13522
rect 4616 13302 4668 13354
rect 4720 13302 4772 13354
rect 4824 13302 4876 13354
rect 11420 13302 11472 13354
rect 11524 13302 11576 13354
rect 11628 13302 11680 13354
rect 18224 13302 18276 13354
rect 18328 13302 18380 13354
rect 18432 13302 18484 13354
rect 25028 13302 25080 13354
rect 25132 13302 25184 13354
rect 25236 13302 25288 13354
rect 12798 13134 12850 13186
rect 4062 13022 4114 13074
rect 7422 13022 7474 13074
rect 14926 13022 14978 13074
rect 21422 13022 21474 13074
rect 27358 13022 27410 13074
rect 28142 13022 28194 13074
rect 1822 12910 1874 12962
rect 5854 12910 5906 12962
rect 9326 12910 9378 12962
rect 9662 12910 9714 12962
rect 15150 12910 15202 12962
rect 22766 12910 22818 12962
rect 23438 12910 23490 12962
rect 26686 12910 26738 12962
rect 26910 12910 26962 12962
rect 3054 12798 3106 12850
rect 6078 12798 6130 12850
rect 8766 12798 8818 12850
rect 12014 12798 12066 12850
rect 20078 12798 20130 12850
rect 2046 12686 2098 12738
rect 6526 12686 6578 12738
rect 25902 12686 25954 12738
rect 26462 12686 26514 12738
rect 27470 12686 27522 12738
rect 8018 12518 8070 12570
rect 8122 12518 8174 12570
rect 8226 12518 8278 12570
rect 14822 12518 14874 12570
rect 14926 12518 14978 12570
rect 15030 12518 15082 12570
rect 21626 12518 21678 12570
rect 21730 12518 21782 12570
rect 21834 12518 21886 12570
rect 28430 12518 28482 12570
rect 28534 12518 28586 12570
rect 28638 12518 28690 12570
rect 7086 12350 7138 12402
rect 8654 12238 8706 12290
rect 18062 12238 18114 12290
rect 23998 12238 24050 12290
rect 27246 12238 27298 12290
rect 1822 12126 1874 12178
rect 3390 12126 3442 12178
rect 3726 12126 3778 12178
rect 4398 12126 4450 12178
rect 4734 12126 4786 12178
rect 14478 12126 14530 12178
rect 20414 12126 20466 12178
rect 20974 12126 21026 12178
rect 21086 12126 21138 12178
rect 21646 12126 21698 12178
rect 3950 12014 4002 12066
rect 8878 12014 8930 12066
rect 10110 12014 10162 12066
rect 25342 12014 25394 12066
rect 25902 12014 25954 12066
rect 26238 12014 26290 12066
rect 7870 11902 7922 11954
rect 17278 11902 17330 11954
rect 24782 11902 24834 11954
rect 4616 11734 4668 11786
rect 4720 11734 4772 11786
rect 4824 11734 4876 11786
rect 11420 11734 11472 11786
rect 11524 11734 11576 11786
rect 11628 11734 11680 11786
rect 18224 11734 18276 11786
rect 18328 11734 18380 11786
rect 18432 11734 18484 11786
rect 25028 11734 25080 11786
rect 25132 11734 25184 11786
rect 25236 11734 25288 11786
rect 7198 11566 7250 11618
rect 3838 11454 3890 11506
rect 23550 11454 23602 11506
rect 27022 11454 27074 11506
rect 10334 11342 10386 11394
rect 10670 11342 10722 11394
rect 15710 11342 15762 11394
rect 16158 11342 16210 11394
rect 19182 11342 19234 11394
rect 21870 11342 21922 11394
rect 4958 11230 5010 11282
rect 7982 11230 8034 11282
rect 11118 11230 11170 11282
rect 11454 11230 11506 11282
rect 11902 11230 11954 11282
rect 12238 11230 12290 11282
rect 19406 11230 19458 11282
rect 19742 11230 19794 11282
rect 20078 11230 20130 11282
rect 27246 11230 27298 11282
rect 27582 11230 27634 11282
rect 12686 11118 12738 11170
rect 18622 11118 18674 11170
rect 20190 11118 20242 11170
rect 27694 11118 27746 11170
rect 8018 10950 8070 11002
rect 8122 10950 8174 11002
rect 8226 10950 8278 11002
rect 14822 10950 14874 11002
rect 14926 10950 14978 11002
rect 15030 10950 15082 11002
rect 21626 10950 21678 11002
rect 21730 10950 21782 11002
rect 21834 10950 21886 11002
rect 28430 10950 28482 11002
rect 28534 10950 28586 11002
rect 28638 10950 28690 11002
rect 4510 10782 4562 10834
rect 5294 10782 5346 10834
rect 8318 10782 8370 10834
rect 11678 10782 11730 10834
rect 15598 10782 15650 10834
rect 23102 10782 23154 10834
rect 23998 10782 24050 10834
rect 28142 10782 28194 10834
rect 9886 10670 9938 10722
rect 16382 10670 16434 10722
rect 27582 10670 27634 10722
rect 1822 10558 1874 10610
rect 2158 10558 2210 10610
rect 5630 10558 5682 10610
rect 6078 10558 6130 10610
rect 12462 10558 12514 10610
rect 13022 10558 13074 10610
rect 19966 10558 20018 10610
rect 20638 10558 20690 10610
rect 24558 10558 24610 10610
rect 11230 10446 11282 10498
rect 16718 10446 16770 10498
rect 17502 10446 17554 10498
rect 19294 10446 19346 10498
rect 19742 10446 19794 10498
rect 24334 10446 24386 10498
rect 26238 10446 26290 10498
rect 9102 10334 9154 10386
rect 16158 10334 16210 10386
rect 23662 10334 23714 10386
rect 4616 10166 4668 10218
rect 4720 10166 4772 10218
rect 4824 10166 4876 10218
rect 11420 10166 11472 10218
rect 11524 10166 11576 10218
rect 11628 10166 11680 10218
rect 18224 10166 18276 10218
rect 18328 10166 18380 10218
rect 18432 10166 18484 10218
rect 25028 10166 25080 10218
rect 25132 10166 25184 10218
rect 25236 10166 25288 10218
rect 9326 9998 9378 10050
rect 28254 9998 28306 10050
rect 19742 9886 19794 9938
rect 23550 9886 23602 9938
rect 5630 9774 5682 9826
rect 6190 9774 6242 9826
rect 12350 9774 12402 9826
rect 12798 9774 12850 9826
rect 15710 9774 15762 9826
rect 16158 9774 16210 9826
rect 20302 9774 20354 9826
rect 21534 9774 21586 9826
rect 24782 9774 24834 9826
rect 25230 9774 25282 9826
rect 4286 9662 4338 9714
rect 4622 9662 4674 9714
rect 10110 9662 10162 9714
rect 19406 9662 19458 9714
rect 20526 9662 20578 9714
rect 27470 9662 27522 9714
rect 5070 9550 5122 9602
rect 8542 9550 8594 9602
rect 9214 9550 9266 9602
rect 18622 9550 18674 9602
rect 19182 9550 19234 9602
rect 8018 9382 8070 9434
rect 8122 9382 8174 9434
rect 8226 9382 8278 9434
rect 14822 9382 14874 9434
rect 14926 9382 14978 9434
rect 15030 9382 15082 9434
rect 21626 9382 21678 9434
rect 21730 9382 21782 9434
rect 21834 9382 21886 9434
rect 28430 9382 28482 9434
rect 28534 9382 28586 9434
rect 28638 9382 28690 9434
rect 5406 9214 5458 9266
rect 20526 9214 20578 9266
rect 21982 9214 22034 9266
rect 28142 9214 28194 9266
rect 8878 9102 8930 9154
rect 10110 9102 10162 9154
rect 15598 9102 15650 9154
rect 23550 9102 23602 9154
rect 24222 9102 24274 9154
rect 27470 9102 27522 9154
rect 2494 8990 2546 9042
rect 2830 8990 2882 9042
rect 12798 8990 12850 9042
rect 13246 8990 13298 9042
rect 17502 8990 17554 9042
rect 18174 8990 18226 9042
rect 24446 8990 24498 9042
rect 7534 8878 7586 8930
rect 11454 8878 11506 8930
rect 21534 8878 21586 8930
rect 22430 8878 22482 8930
rect 26238 8878 26290 8930
rect 5966 8766 6018 8818
rect 16382 8766 16434 8818
rect 21198 8766 21250 8818
rect 4616 8598 4668 8650
rect 4720 8598 4772 8650
rect 4824 8598 4876 8650
rect 11420 8598 11472 8650
rect 11524 8598 11576 8650
rect 11628 8598 11680 8650
rect 18224 8598 18276 8650
rect 18328 8598 18380 8650
rect 18432 8598 18484 8650
rect 25028 8598 25080 8650
rect 25132 8598 25184 8650
rect 25236 8598 25288 8650
rect 3614 8318 3666 8370
rect 5742 8318 5794 8370
rect 6078 8318 6130 8370
rect 7422 8318 7474 8370
rect 9326 8318 9378 8370
rect 15150 8318 15202 8370
rect 17614 8318 17666 8370
rect 22318 8318 22370 8370
rect 28254 8318 28306 8370
rect 12462 8206 12514 8258
rect 12798 8206 12850 8258
rect 14142 8206 14194 8258
rect 24558 8206 24610 8258
rect 25230 8206 25282 8258
rect 2494 8094 2546 8146
rect 8654 8094 8706 8146
rect 18622 8094 18674 8146
rect 23550 8094 23602 8146
rect 6526 7982 6578 8034
rect 10110 7982 10162 8034
rect 16830 7982 16882 8034
rect 27694 7982 27746 8034
rect 8018 7814 8070 7866
rect 8122 7814 8174 7866
rect 8226 7814 8278 7866
rect 14822 7814 14874 7866
rect 14926 7814 14978 7866
rect 15030 7814 15082 7866
rect 21626 7814 21678 7866
rect 21730 7814 21782 7866
rect 21834 7814 21886 7866
rect 28430 7814 28482 7866
rect 28534 7814 28586 7866
rect 28638 7814 28690 7866
rect 1598 7646 1650 7698
rect 2382 7646 2434 7698
rect 21870 7646 21922 7698
rect 25342 7646 25394 7698
rect 7198 7534 7250 7586
rect 9774 7534 9826 7586
rect 12462 7534 12514 7586
rect 16270 7534 16322 7586
rect 27246 7534 27298 7586
rect 28142 7534 28194 7586
rect 4734 7422 4786 7474
rect 5294 7422 5346 7474
rect 12686 7422 12738 7474
rect 24222 7422 24274 7474
rect 24558 7422 24610 7474
rect 6190 7310 6242 7362
rect 11118 7310 11170 7362
rect 13246 7310 13298 7362
rect 14926 7310 14978 7362
rect 26238 7310 26290 7362
rect 21086 7198 21138 7250
rect 4616 7030 4668 7082
rect 4720 7030 4772 7082
rect 4824 7030 4876 7082
rect 11420 7030 11472 7082
rect 11524 7030 11576 7082
rect 11628 7030 11680 7082
rect 18224 7030 18276 7082
rect 18328 7030 18380 7082
rect 18432 7030 18484 7082
rect 25028 7030 25080 7082
rect 25132 7030 25184 7082
rect 25236 7030 25288 7082
rect 14478 6750 14530 6802
rect 7982 6638 8034 6690
rect 8206 6638 8258 6690
rect 8654 6638 8706 6690
rect 23998 6638 24050 6690
rect 24446 6638 24498 6690
rect 27470 6638 27522 6690
rect 27694 6638 27746 6690
rect 15822 6526 15874 6578
rect 21646 6526 21698 6578
rect 21982 6526 22034 6578
rect 22318 6414 22370 6466
rect 23102 6414 23154 6466
rect 26798 6414 26850 6466
rect 27806 6414 27858 6466
rect 8018 6246 8070 6298
rect 8122 6246 8174 6298
rect 8226 6246 8278 6298
rect 14822 6246 14874 6298
rect 14926 6246 14978 6298
rect 15030 6246 15082 6298
rect 21626 6246 21678 6298
rect 21730 6246 21782 6298
rect 21834 6246 21886 6298
rect 28430 6246 28482 6298
rect 28534 6246 28586 6298
rect 28638 6246 28690 6298
rect 14814 6078 14866 6130
rect 26350 6078 26402 6130
rect 13806 5966 13858 6018
rect 15150 5966 15202 6018
rect 15486 5966 15538 6018
rect 20862 5966 20914 6018
rect 22542 5966 22594 6018
rect 24670 5966 24722 6018
rect 27694 5966 27746 6018
rect 13470 5854 13522 5906
rect 21198 5854 21250 5906
rect 20638 5742 20690 5794
rect 21534 5742 21586 5794
rect 24334 5742 24386 5794
rect 26686 5742 26738 5794
rect 4616 5462 4668 5514
rect 4720 5462 4772 5514
rect 4824 5462 4876 5514
rect 11420 5462 11472 5514
rect 11524 5462 11576 5514
rect 11628 5462 11680 5514
rect 18224 5462 18276 5514
rect 18328 5462 18380 5514
rect 18432 5462 18484 5514
rect 25028 5462 25080 5514
rect 25132 5462 25184 5514
rect 25236 5462 25288 5514
rect 23326 5182 23378 5234
rect 19406 5070 19458 5122
rect 24558 5070 24610 5122
rect 25230 5070 25282 5122
rect 19630 4958 19682 5010
rect 19966 4958 20018 5010
rect 22318 4958 22370 5010
rect 20302 4846 20354 4898
rect 21534 4846 21586 4898
rect 27694 4846 27746 4898
rect 28254 4846 28306 4898
rect 8018 4678 8070 4730
rect 8122 4678 8174 4730
rect 8226 4678 8278 4730
rect 14822 4678 14874 4730
rect 14926 4678 14978 4730
rect 15030 4678 15082 4730
rect 21626 4678 21678 4730
rect 21730 4678 21782 4730
rect 21834 4678 21886 4730
rect 28430 4678 28482 4730
rect 28534 4678 28586 4730
rect 28638 4678 28690 4730
rect 24222 4510 24274 4562
rect 24782 4510 24834 4562
rect 25342 4510 25394 4562
rect 25902 4510 25954 4562
rect 14142 4398 14194 4450
rect 14926 4398 14978 4450
rect 15262 4398 15314 4450
rect 18062 4398 18114 4450
rect 19294 4398 19346 4450
rect 27246 4398 27298 4450
rect 28142 4398 28194 4450
rect 14702 4286 14754 4338
rect 19070 4286 19122 4338
rect 20750 4286 20802 4338
rect 21310 4286 21362 4338
rect 21646 4286 21698 4338
rect 12798 4174 12850 4226
rect 18734 4174 18786 4226
rect 19742 4174 19794 4226
rect 20414 4174 20466 4226
rect 26238 4174 26290 4226
rect 4616 3894 4668 3946
rect 4720 3894 4772 3946
rect 4824 3894 4876 3946
rect 11420 3894 11472 3946
rect 11524 3894 11576 3946
rect 11628 3894 11680 3946
rect 18224 3894 18276 3946
rect 18328 3894 18380 3946
rect 18432 3894 18484 3946
rect 25028 3894 25080 3946
rect 25132 3894 25184 3946
rect 25236 3894 25288 3946
rect 15598 3614 15650 3666
rect 21534 3614 21586 3666
rect 23102 3614 23154 3666
rect 26126 3614 26178 3666
rect 14254 3502 14306 3554
rect 15150 3502 15202 3554
rect 17166 3502 17218 3554
rect 18510 3502 18562 3554
rect 19406 3502 19458 3554
rect 20078 3502 20130 3554
rect 22318 3502 22370 3554
rect 22654 3502 22706 3554
rect 12238 3390 12290 3442
rect 12574 3390 12626 3442
rect 16494 3390 16546 3442
rect 16942 3390 16994 3442
rect 19070 3390 19122 3442
rect 19854 3390 19906 3442
rect 21086 3390 21138 3442
rect 27470 3390 27522 3442
rect 13134 3278 13186 3330
rect 13582 3278 13634 3330
rect 17614 3278 17666 3330
rect 18734 3278 18786 3330
rect 24782 3278 24834 3330
rect 8018 3110 8070 3162
rect 8122 3110 8174 3162
rect 8226 3110 8278 3162
rect 14822 3110 14874 3162
rect 14926 3110 14978 3162
rect 15030 3110 15082 3162
rect 21626 3110 21678 3162
rect 21730 3110 21782 3162
rect 21834 3110 21886 3162
rect 28430 3110 28482 3162
rect 28534 3110 28586 3162
rect 28638 3110 28690 3162
rect 16830 1710 16882 1762
rect 17614 1710 17666 1762
<< metal2 >>
rect 7392 29200 7504 30000
rect 8064 29200 8176 30000
rect 8736 29200 8848 30000
rect 9408 29200 9520 30000
rect 10080 29200 10192 30000
rect 10752 29200 10864 30000
rect 11424 29200 11536 30000
rect 12096 29200 12208 30000
rect 12768 29200 12880 30000
rect 13440 29200 13552 30000
rect 14112 29200 14224 30000
rect 14784 29200 14896 30000
rect 15456 29200 15568 30000
rect 16128 29200 16240 30000
rect 16800 29200 16912 30000
rect 17472 29200 17584 30000
rect 18144 29200 18256 30000
rect 18816 29200 18928 30000
rect 19488 29200 19600 30000
rect 20160 29200 20272 30000
rect 20832 29200 20944 30000
rect 21504 29200 21616 30000
rect 22176 29200 22288 30000
rect 22848 29200 22960 30000
rect 24864 29200 24976 30000
rect 7420 26516 7476 29200
rect 8092 27412 8148 29200
rect 7868 27356 8148 27412
rect 7644 26516 7700 26526
rect 7420 26514 7700 26516
rect 7420 26462 7646 26514
rect 7698 26462 7700 26514
rect 7420 26460 7700 26462
rect 7868 26516 7924 27356
rect 8016 26684 8280 26694
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8016 26618 8280 26628
rect 8204 26516 8260 26526
rect 7868 26514 8260 26516
rect 7868 26462 8206 26514
rect 8258 26462 8260 26514
rect 7868 26460 8260 26462
rect 7644 26450 7700 26460
rect 8204 26450 8260 26460
rect 8764 26514 8820 29200
rect 9436 26964 9492 29200
rect 9436 26908 9940 26964
rect 8764 26462 8766 26514
rect 8818 26462 8820 26514
rect 8764 26450 8820 26462
rect 9660 26404 9716 26414
rect 9324 26402 9716 26404
rect 9324 26350 9662 26402
rect 9714 26350 9716 26402
rect 9324 26348 9716 26350
rect 4614 25900 4878 25910
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4614 25834 4878 25844
rect 1708 25284 1764 25294
rect 1708 25190 1764 25228
rect 8016 25116 8280 25126
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8016 25050 8280 25060
rect 4614 24332 4878 24342
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4614 24266 4878 24276
rect 9324 23938 9380 26348
rect 9660 26338 9716 26348
rect 9884 26292 9940 26908
rect 10108 26850 10164 29200
rect 10108 26798 10110 26850
rect 10162 26798 10164 26850
rect 10108 26786 10164 26798
rect 9772 26290 9940 26292
rect 9772 26238 9886 26290
rect 9938 26238 9940 26290
rect 9772 26236 9940 26238
rect 9772 26180 9828 26236
rect 9884 26226 9940 26236
rect 10332 26290 10388 26302
rect 10332 26238 10334 26290
rect 10386 26238 10388 26290
rect 9436 26124 9828 26180
rect 9436 25618 9492 26124
rect 9436 25566 9438 25618
rect 9490 25566 9492 25618
rect 9436 25554 9492 25566
rect 9324 23886 9326 23938
rect 9378 23886 9380 23938
rect 9324 23874 9380 23886
rect 9548 25284 9604 25294
rect 9548 23826 9604 25228
rect 10332 25284 10388 26238
rect 10780 25620 10836 29200
rect 11116 26850 11172 26862
rect 11116 26798 11118 26850
rect 11170 26798 11172 26850
rect 11116 26514 11172 26798
rect 11452 26628 11508 29200
rect 11452 26572 11732 26628
rect 11116 26462 11118 26514
rect 11170 26462 11172 26514
rect 11116 26450 11172 26462
rect 11676 26068 11732 26572
rect 12012 26516 12068 26526
rect 12124 26516 12180 29200
rect 12012 26514 12292 26516
rect 12012 26462 12014 26514
rect 12066 26462 12292 26514
rect 12012 26460 12292 26462
rect 12012 26450 12068 26460
rect 12236 26402 12292 26460
rect 12236 26350 12238 26402
rect 12290 26350 12292 26402
rect 12236 26338 12292 26350
rect 12572 26402 12628 26414
rect 12572 26350 12574 26402
rect 12626 26350 12628 26402
rect 11676 26012 11844 26068
rect 11418 25900 11682 25910
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11418 25834 11682 25844
rect 11788 25732 11844 26012
rect 11676 25676 11844 25732
rect 10780 25618 11060 25620
rect 10780 25566 10782 25618
rect 10834 25566 11060 25618
rect 10780 25564 11060 25566
rect 10780 25554 10836 25564
rect 11004 25506 11060 25564
rect 11004 25454 11006 25506
rect 11058 25454 11060 25506
rect 11004 25442 11060 25454
rect 11676 25394 11732 25676
rect 12572 25506 12628 26350
rect 12796 25732 12852 29200
rect 13468 27858 13524 29200
rect 14140 28084 14196 29200
rect 13468 27806 13470 27858
rect 13522 27806 13524 27858
rect 13468 27794 13524 27806
rect 14028 28028 14196 28084
rect 13356 26516 13412 26526
rect 13356 26422 13412 26460
rect 14028 26516 14084 28028
rect 14028 26450 14084 26460
rect 14140 27858 14196 27870
rect 14140 27806 14142 27858
rect 14194 27806 14196 27858
rect 12796 25666 12852 25676
rect 12908 26292 12964 26302
rect 12572 25454 12574 25506
rect 12626 25454 12628 25506
rect 12572 25442 12628 25454
rect 11676 25342 11678 25394
rect 11730 25342 11732 25394
rect 11676 25330 11732 25342
rect 12908 25394 12964 26236
rect 13692 26292 13748 26302
rect 13692 26198 13748 26236
rect 14140 26178 14196 27806
rect 14812 27076 14868 29200
rect 14700 27020 14868 27076
rect 14700 26516 14756 27020
rect 14820 26684 15084 26694
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 14820 26618 15084 26628
rect 14700 26460 15092 26516
rect 14140 26126 14142 26178
rect 14194 26126 14196 26178
rect 14140 26114 14196 26126
rect 13916 25732 13972 25742
rect 13916 25618 13972 25676
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 13916 25554 13972 25566
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12908 25330 12964 25342
rect 15036 25394 15092 26460
rect 15036 25342 15038 25394
rect 15090 25342 15092 25394
rect 15036 25330 15092 25342
rect 15372 26402 15428 26414
rect 15372 26350 15374 26402
rect 15426 26350 15428 26402
rect 10332 25218 10388 25228
rect 11340 25284 11396 25294
rect 11340 25190 11396 25228
rect 12796 25284 12852 25294
rect 13468 25284 13524 25294
rect 12796 24834 12852 25228
rect 13132 25282 13524 25284
rect 13132 25230 13470 25282
rect 13522 25230 13524 25282
rect 13132 25228 13524 25230
rect 13132 24946 13188 25228
rect 13468 25218 13524 25228
rect 14820 25116 15084 25126
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 14820 25050 15084 25060
rect 13132 24894 13134 24946
rect 13186 24894 13188 24946
rect 13132 24882 13188 24894
rect 12796 24782 12798 24834
rect 12850 24782 12852 24834
rect 12796 24770 12852 24782
rect 11418 24332 11682 24342
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11418 24266 11682 24276
rect 9548 23774 9550 23826
rect 9602 23774 9604 23826
rect 9548 23762 9604 23774
rect 8016 23548 8280 23558
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8016 23482 8280 23492
rect 14820 23548 15084 23558
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 14820 23482 15084 23492
rect 4614 22764 4878 22774
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4614 22698 4878 22708
rect 11418 22764 11682 22774
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11418 22698 11682 22708
rect 8016 21980 8280 21990
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8016 21914 8280 21924
rect 14820 21980 15084 21990
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 14820 21914 15084 21924
rect 15372 21698 15428 26350
rect 15484 26292 15540 29200
rect 16044 26402 16100 26414
rect 16044 26350 16046 26402
rect 16098 26350 16100 26402
rect 15596 26292 15652 26302
rect 15484 26290 15988 26292
rect 15484 26238 15598 26290
rect 15650 26238 15988 26290
rect 15484 26236 15988 26238
rect 15596 26226 15652 26236
rect 15932 25618 15988 26236
rect 15932 25566 15934 25618
rect 15986 25566 15988 25618
rect 15932 25554 15988 25566
rect 15708 21812 15764 21822
rect 15708 21718 15764 21756
rect 15372 21646 15374 21698
rect 15426 21646 15428 21698
rect 15372 21634 15428 21646
rect 16044 21698 16100 26350
rect 16156 26292 16212 29200
rect 16828 26850 16884 29200
rect 17500 27188 17556 29200
rect 17500 27132 17668 27188
rect 16828 26798 16830 26850
rect 16882 26798 16884 26850
rect 16828 26786 16884 26798
rect 17500 26850 17556 26862
rect 17500 26798 17502 26850
rect 17554 26798 17556 26850
rect 16268 26292 16324 26302
rect 17052 26292 17108 26302
rect 16156 26236 16268 26292
rect 16268 26198 16324 26236
rect 16716 26290 17108 26292
rect 16716 26238 17054 26290
rect 17106 26238 17108 26290
rect 16716 26236 17108 26238
rect 16492 25620 16548 25630
rect 16492 25506 16548 25564
rect 16492 25454 16494 25506
rect 16546 25454 16548 25506
rect 16492 25442 16548 25454
rect 16716 25394 16772 26236
rect 17052 26226 17108 26236
rect 17164 26292 17220 26302
rect 17164 25618 17220 26236
rect 17500 26178 17556 26798
rect 17612 26516 17668 27132
rect 18172 26852 18228 29200
rect 18172 26786 18228 26796
rect 18844 26850 18900 29200
rect 18844 26798 18846 26850
rect 18898 26798 18900 26850
rect 18844 26786 18900 26798
rect 18956 26852 19012 26862
rect 17612 26450 17668 26460
rect 17500 26126 17502 26178
rect 17554 26126 17556 26178
rect 17500 26114 17556 26126
rect 18732 26290 18788 26302
rect 18732 26238 18734 26290
rect 18786 26238 18788 26290
rect 18222 25900 18486 25910
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18222 25834 18486 25844
rect 17164 25566 17166 25618
rect 17218 25566 17220 25618
rect 17164 25554 17220 25566
rect 18508 25508 18564 25518
rect 18508 25506 18676 25508
rect 18508 25454 18510 25506
rect 18562 25454 18676 25506
rect 18508 25452 18676 25454
rect 18508 25442 18564 25452
rect 16716 25342 16718 25394
rect 16770 25342 16772 25394
rect 16716 25330 16772 25342
rect 18222 24332 18486 24342
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18222 24266 18486 24276
rect 18222 22764 18486 22774
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18222 22698 18486 22708
rect 18620 21812 18676 25452
rect 18620 21746 18676 21756
rect 16044 21646 16046 21698
rect 16098 21646 16100 21698
rect 16044 21634 16100 21646
rect 16380 21700 16436 21710
rect 16380 21606 16436 21644
rect 18732 21700 18788 26238
rect 18956 25618 19012 26796
rect 19068 26516 19124 26526
rect 19068 26178 19124 26460
rect 19516 26516 19572 29200
rect 20188 27300 20244 29200
rect 20188 27244 20692 27300
rect 19516 26450 19572 26460
rect 19628 26850 19684 26862
rect 19628 26798 19630 26850
rect 19682 26798 19684 26850
rect 19068 26126 19070 26178
rect 19122 26126 19124 26178
rect 19068 26114 19124 26126
rect 18956 25566 18958 25618
rect 19010 25566 19012 25618
rect 18956 25554 19012 25566
rect 19628 25618 19684 26798
rect 19628 25566 19630 25618
rect 19682 25566 19684 25618
rect 19628 25508 19684 25566
rect 19628 25442 19684 25452
rect 20188 25508 20244 25518
rect 20188 25414 20244 25452
rect 19068 25396 19124 25406
rect 18956 25284 19012 25294
rect 18844 23940 18900 23950
rect 18956 23940 19012 25228
rect 18844 23938 19012 23940
rect 18844 23886 18846 23938
rect 18898 23886 19012 23938
rect 18844 23884 19012 23886
rect 18844 23874 18900 23884
rect 19068 23826 19124 25340
rect 20636 25394 20692 27244
rect 20636 25342 20638 25394
rect 20690 25342 20692 25394
rect 20636 25330 20692 25342
rect 20748 26290 20804 26302
rect 20748 26238 20750 26290
rect 20802 26238 20804 26290
rect 20748 25396 20804 26238
rect 20860 25508 20916 29200
rect 21532 26852 21588 29200
rect 21532 26786 21588 26796
rect 22204 26850 22260 29200
rect 22204 26798 22206 26850
rect 22258 26798 22260 26850
rect 22204 26786 22260 26798
rect 22764 26852 22820 26862
rect 21624 26684 21888 26694
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21624 26618 21888 26628
rect 21196 26516 21252 26526
rect 21196 26178 21252 26460
rect 22316 26292 22372 26302
rect 21196 26126 21198 26178
rect 21250 26126 21252 26178
rect 21196 26114 21252 26126
rect 21644 26290 22372 26292
rect 21644 26238 22318 26290
rect 22370 26238 22372 26290
rect 21644 26236 22372 26238
rect 20860 25442 20916 25452
rect 21308 25508 21364 25518
rect 20748 25330 20804 25340
rect 19964 25284 20020 25294
rect 19964 25190 20020 25228
rect 21308 24948 21364 25452
rect 21420 25506 21476 25518
rect 21420 25454 21422 25506
rect 21474 25454 21476 25506
rect 21420 25284 21476 25454
rect 21644 25394 21700 26236
rect 22316 26226 22372 26236
rect 22764 26178 22820 26796
rect 22876 26516 22932 29200
rect 22876 26450 22932 26460
rect 22988 26850 23044 26862
rect 22988 26798 22990 26850
rect 23042 26798 23044 26850
rect 22764 26126 22766 26178
rect 22818 26126 22820 26178
rect 22764 26114 22820 26126
rect 22652 25620 22708 25630
rect 22204 25508 22260 25518
rect 22204 25414 22260 25452
rect 21644 25342 21646 25394
rect 21698 25342 21700 25394
rect 21644 25330 21700 25342
rect 22652 25394 22708 25564
rect 22988 25508 23044 26798
rect 23884 26516 23940 26526
rect 24892 26516 24948 29200
rect 28140 26852 28196 26862
rect 25116 26516 25172 26526
rect 24892 26514 25172 26516
rect 24892 26462 25118 26514
rect 25170 26462 25172 26514
rect 24892 26460 25172 26462
rect 23884 26422 23940 26460
rect 25116 26450 25172 26460
rect 26236 26402 26292 26414
rect 26236 26350 26238 26402
rect 26290 26350 26292 26402
rect 26236 26292 26292 26350
rect 26236 26226 26292 26236
rect 26796 26292 26852 26302
rect 26796 26290 27076 26292
rect 26796 26238 26798 26290
rect 26850 26238 27076 26290
rect 26796 26236 27076 26238
rect 26796 26226 26852 26236
rect 25026 25900 25290 25910
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25026 25834 25290 25844
rect 22652 25342 22654 25394
rect 22706 25342 22708 25394
rect 22652 25330 22708 25342
rect 22764 25506 23044 25508
rect 22764 25454 22990 25506
rect 23042 25454 23044 25506
rect 22764 25452 23044 25454
rect 21420 25218 21476 25228
rect 21980 25284 22036 25294
rect 21980 25190 22036 25228
rect 22764 25172 22820 25452
rect 22988 25442 23044 25452
rect 21624 25116 21888 25126
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21624 25050 21888 25060
rect 22428 25116 22820 25172
rect 21756 24948 21812 24958
rect 21308 24946 21812 24948
rect 21308 24894 21758 24946
rect 21810 24894 21812 24946
rect 21308 24892 21812 24894
rect 21756 24882 21812 24892
rect 22428 24946 22484 25116
rect 22428 24894 22430 24946
rect 22482 24894 22484 24946
rect 22428 24882 22484 24894
rect 27020 24946 27076 26236
rect 27692 26178 27748 26190
rect 27692 26126 27694 26178
rect 27746 26126 27748 26178
rect 27692 25620 27748 26126
rect 27692 25554 27748 25564
rect 27132 25508 27188 25518
rect 27132 25414 27188 25452
rect 28140 25508 28196 26796
rect 28428 26684 28692 26694
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28428 26618 28692 26628
rect 28140 25414 28196 25452
rect 27468 25284 27524 25294
rect 27804 25284 27860 25294
rect 27468 25190 27524 25228
rect 27580 25282 27860 25284
rect 27580 25230 27806 25282
rect 27858 25230 27860 25282
rect 27580 25228 27860 25230
rect 27020 24894 27022 24946
rect 27074 24894 27076 24946
rect 27020 24882 27076 24894
rect 27356 24836 27412 24846
rect 27580 24836 27636 25228
rect 27804 25218 27860 25228
rect 28428 25116 28692 25126
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28428 25050 28692 25060
rect 27356 24834 27636 24836
rect 27356 24782 27358 24834
rect 27410 24782 27636 24834
rect 27356 24780 27636 24782
rect 28140 24834 28196 24846
rect 28140 24782 28142 24834
rect 28194 24782 28196 24834
rect 27356 24770 27412 24780
rect 25026 24332 25290 24342
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25026 24266 25290 24276
rect 28140 24276 28196 24782
rect 28140 24210 28196 24220
rect 19068 23774 19070 23826
rect 19122 23774 19124 23826
rect 19068 23762 19124 23774
rect 27692 23716 27748 23726
rect 27692 23622 27748 23660
rect 28140 23716 28196 23726
rect 28140 23714 28308 23716
rect 28140 23662 28142 23714
rect 28194 23662 28308 23714
rect 28140 23660 28308 23662
rect 28140 23650 28196 23660
rect 21624 23548 21888 23558
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21624 23482 21888 23492
rect 27132 23266 27188 23278
rect 27132 23214 27134 23266
rect 27186 23214 27188 23266
rect 26908 23044 26964 23054
rect 26908 22950 26964 22988
rect 25026 22764 25290 22774
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25026 22698 25290 22708
rect 27132 22370 27188 23214
rect 27468 23268 27524 23278
rect 27804 23268 27860 23278
rect 27468 23266 27860 23268
rect 27468 23214 27470 23266
rect 27522 23214 27806 23266
rect 27858 23214 27860 23266
rect 27468 23212 27860 23214
rect 27468 23202 27524 23212
rect 27804 23202 27860 23212
rect 27132 22318 27134 22370
rect 27186 22318 27188 22370
rect 27132 22306 27188 22318
rect 28140 23154 28196 23166
rect 28140 23102 28142 23154
rect 28194 23102 28196 23154
rect 28140 23044 28196 23102
rect 28028 22260 28084 22270
rect 28028 22166 28084 22204
rect 21624 21980 21888 21990
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21624 21914 21888 21924
rect 18732 21634 18788 21644
rect 24892 21700 24948 21710
rect 23660 21476 23716 21486
rect 4614 21196 4878 21206
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4614 21130 4878 21140
rect 11418 21196 11682 21206
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11418 21130 11682 21140
rect 18222 21196 18486 21206
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18222 21130 18486 21140
rect 22988 20804 23044 20814
rect 22764 20802 23044 20804
rect 22764 20750 22990 20802
rect 23042 20750 23044 20802
rect 22764 20748 23044 20750
rect 17276 20578 17332 20590
rect 17276 20526 17278 20578
rect 17330 20526 17332 20578
rect 8016 20412 8280 20422
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8016 20346 8280 20356
rect 14820 20412 15084 20422
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 14820 20346 15084 20356
rect 11788 20130 11844 20142
rect 14028 20132 14084 20142
rect 11788 20078 11790 20130
rect 11842 20078 11844 20130
rect 8764 19908 8820 19918
rect 4614 19628 4878 19638
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4614 19562 4878 19572
rect 8652 19346 8708 19358
rect 8652 19294 8654 19346
rect 8706 19294 8708 19346
rect 8016 18844 8280 18854
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8016 18778 8280 18788
rect 5404 18676 5460 18686
rect 8316 18676 8372 18686
rect 5404 18674 5684 18676
rect 5404 18622 5406 18674
rect 5458 18622 5684 18674
rect 5404 18620 5684 18622
rect 5404 18610 5460 18620
rect 2492 18450 2548 18462
rect 2492 18398 2494 18450
rect 2546 18398 2548 18450
rect 1820 18340 1876 18350
rect 1708 18338 1876 18340
rect 1708 18286 1822 18338
rect 1874 18286 1876 18338
rect 1708 18284 1876 18286
rect 1708 17442 1764 18284
rect 1820 18274 1876 18284
rect 2268 17668 2324 17678
rect 2268 17574 2324 17612
rect 1708 17390 1710 17442
rect 1762 17390 1764 17442
rect 1708 16884 1764 17390
rect 1708 16818 1764 16828
rect 2044 16994 2100 17006
rect 2044 16942 2046 16994
rect 2098 16942 2100 16994
rect 2044 15538 2100 16942
rect 2492 16884 2548 18398
rect 2492 16818 2548 16828
rect 2940 18450 2996 18462
rect 2940 18398 2942 18450
rect 2994 18398 2996 18450
rect 2940 16772 2996 18398
rect 5292 18340 5348 18350
rect 4614 18060 4878 18070
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4614 17994 4878 18004
rect 4620 16884 4676 16894
rect 4620 16790 4676 16828
rect 5292 16882 5348 18284
rect 5292 16830 5294 16882
rect 5346 16830 5348 16882
rect 5292 16818 5348 16830
rect 3164 16772 3220 16782
rect 2940 16770 3220 16772
rect 2940 16718 3166 16770
rect 3218 16718 3220 16770
rect 2940 16716 3220 16718
rect 3164 16706 3220 16716
rect 5516 16772 5572 16782
rect 4614 16492 4878 16502
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4614 16426 4878 16436
rect 5516 16100 5572 16716
rect 5628 16210 5684 18620
rect 5964 18564 6020 18574
rect 5964 18470 6020 18508
rect 7196 18340 7252 18350
rect 7196 18246 7252 18284
rect 5628 16158 5630 16210
rect 5682 16158 5684 16210
rect 5628 16146 5684 16158
rect 7308 17780 7364 17790
rect 2044 15486 2046 15538
rect 2098 15486 2100 15538
rect 2044 15474 2100 15486
rect 2828 15988 2884 15998
rect 2828 15538 2884 15932
rect 4732 15988 4788 15998
rect 4732 15894 4788 15932
rect 5068 15988 5124 15998
rect 5068 15986 5236 15988
rect 5068 15934 5070 15986
rect 5122 15934 5236 15986
rect 5068 15932 5236 15934
rect 5068 15922 5124 15932
rect 2828 15486 2830 15538
rect 2882 15486 2884 15538
rect 2828 15474 2884 15486
rect 4172 15428 4228 15438
rect 4060 15316 4116 15326
rect 4060 14642 4116 15260
rect 4060 14590 4062 14642
rect 4114 14590 4116 14642
rect 4060 14578 4116 14590
rect 3052 14418 3108 14430
rect 3052 14366 3054 14418
rect 3106 14366 3108 14418
rect 3052 14308 3108 14366
rect 3052 14242 3108 14252
rect 4172 13970 4228 15372
rect 5068 15316 5124 15326
rect 5068 15222 5124 15260
rect 5180 15092 5236 15932
rect 5516 15314 5572 16044
rect 6636 16100 6692 16110
rect 6636 16006 6692 16044
rect 7308 16098 7364 17724
rect 8092 17668 8148 17678
rect 7868 17666 8148 17668
rect 7868 17614 8094 17666
rect 8146 17614 8148 17666
rect 7868 17612 8148 17614
rect 7420 17554 7476 17566
rect 7420 17502 7422 17554
rect 7474 17502 7476 17554
rect 7420 16884 7476 17502
rect 7532 17442 7588 17454
rect 7532 17390 7534 17442
rect 7586 17390 7588 17442
rect 7532 17106 7588 17390
rect 7532 17054 7534 17106
rect 7586 17054 7588 17106
rect 7532 17042 7588 17054
rect 7420 16818 7476 16828
rect 7308 16046 7310 16098
rect 7362 16046 7364 16098
rect 7308 16034 7364 16046
rect 7756 16100 7812 16110
rect 7868 16100 7924 17612
rect 8092 17602 8148 17612
rect 8316 17444 8372 18620
rect 8428 18564 8484 18574
rect 8428 18470 8484 18508
rect 8652 18004 8708 19294
rect 8652 17938 8708 17948
rect 8764 17666 8820 19852
rect 10668 19908 10724 19918
rect 10668 19814 10724 19852
rect 11418 19628 11682 19638
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11418 19562 11682 19572
rect 11452 19348 11508 19358
rect 11116 19346 11508 19348
rect 11116 19294 11454 19346
rect 11506 19294 11508 19346
rect 11116 19292 11508 19294
rect 9660 19122 9716 19134
rect 9660 19070 9662 19122
rect 9714 19070 9716 19122
rect 9660 18676 9716 19070
rect 9660 18610 9716 18620
rect 10668 18450 10724 18462
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 8764 17614 8766 17666
rect 8818 17614 8820 17666
rect 8764 17602 8820 17614
rect 10332 18228 10388 18238
rect 8316 17388 8484 17444
rect 8016 17276 8280 17286
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8016 17210 8280 17220
rect 8316 17108 8372 17118
rect 8428 17108 8484 17388
rect 8316 17106 8484 17108
rect 8316 17054 8318 17106
rect 8370 17054 8484 17106
rect 8316 17052 8484 17054
rect 8316 17042 8372 17052
rect 7812 16044 7924 16100
rect 7756 16034 7812 16044
rect 5964 15988 6020 15998
rect 5964 15986 6244 15988
rect 5964 15934 5966 15986
rect 6018 15934 6244 15986
rect 5964 15932 6244 15934
rect 5964 15922 6020 15932
rect 5516 15262 5518 15314
rect 5570 15262 5572 15314
rect 5516 15250 5572 15262
rect 5292 15092 5348 15102
rect 5180 15036 5292 15092
rect 5292 15026 5348 15036
rect 6188 15092 6244 15932
rect 6748 15428 6804 15438
rect 6748 15334 6804 15372
rect 7868 15428 7924 16044
rect 8988 16884 9044 16894
rect 8016 15708 8280 15718
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8016 15642 8280 15652
rect 4614 14924 4878 14934
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4614 14858 4878 14868
rect 4172 13918 4174 13970
rect 4226 13918 4228 13970
rect 4172 13906 4228 13918
rect 4956 14420 5012 14430
rect 4956 13970 5012 14364
rect 6076 14420 6132 14430
rect 6188 14420 6244 15036
rect 6412 14420 6468 14430
rect 6188 14418 6468 14420
rect 6188 14366 6414 14418
rect 6466 14366 6468 14418
rect 6188 14364 6468 14366
rect 6076 14326 6132 14364
rect 4956 13918 4958 13970
rect 5010 13918 5012 13970
rect 4956 13906 5012 13918
rect 6412 13636 6468 14364
rect 6636 14308 6692 14318
rect 6636 14214 6692 14252
rect 7420 14308 7476 14318
rect 7420 14214 7476 14252
rect 6412 13570 6468 13580
rect 7308 13746 7364 13758
rect 7308 13694 7310 13746
rect 7362 13694 7364 13746
rect 4614 13356 4878 13366
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4614 13290 4878 13300
rect 4060 13074 4116 13086
rect 4060 13022 4062 13074
rect 4114 13022 4116 13074
rect 1820 12962 1876 12974
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1820 12180 1876 12910
rect 4060 12964 4116 13022
rect 7308 13076 7364 13694
rect 7868 13746 7924 15372
rect 7980 15202 8036 15214
rect 7980 15150 7982 15202
rect 8034 15150 8036 15202
rect 7980 14868 8036 15150
rect 7980 14802 8036 14812
rect 8988 14420 9044 16828
rect 9772 16884 9828 16894
rect 9772 16790 9828 16828
rect 9548 16770 9604 16782
rect 9548 16718 9550 16770
rect 9602 16718 9604 16770
rect 9548 15986 9604 16718
rect 10332 16322 10388 18172
rect 10668 16882 10724 18398
rect 11116 18450 11172 19292
rect 11452 19282 11508 19292
rect 11788 19236 11844 20078
rect 13916 20130 14084 20132
rect 13916 20078 14030 20130
rect 14082 20078 14084 20130
rect 13916 20076 14084 20078
rect 13916 20018 13972 20076
rect 14028 20066 14084 20076
rect 14140 20132 14196 20142
rect 13916 19966 13918 20018
rect 13970 19966 13972 20018
rect 13916 19954 13972 19966
rect 13580 19906 13636 19918
rect 13580 19854 13582 19906
rect 13634 19854 13636 19906
rect 11116 18398 11118 18450
rect 11170 18398 11172 18450
rect 11116 18386 11172 18398
rect 11676 19180 11844 19236
rect 13468 19234 13524 19246
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 11676 18228 11732 19180
rect 12460 19124 12516 19134
rect 11676 18162 11732 18172
rect 11788 19122 12516 19124
rect 11788 19070 12462 19122
rect 12514 19070 12516 19122
rect 11788 19068 12516 19070
rect 11418 18060 11682 18070
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11418 17994 11682 18004
rect 11788 17890 11844 19068
rect 12460 19058 12516 19068
rect 11788 17838 11790 17890
rect 11842 17838 11844 17890
rect 11788 17826 11844 17838
rect 11228 17556 11284 17566
rect 11228 17442 11284 17500
rect 12012 17556 12068 17566
rect 12012 17462 12068 17500
rect 12348 17554 12404 17566
rect 12348 17502 12350 17554
rect 12402 17502 12404 17554
rect 11228 17390 11230 17442
rect 11282 17390 11284 17442
rect 11228 17378 11284 17390
rect 10668 16830 10670 16882
rect 10722 16830 10724 16882
rect 10668 16772 10724 16830
rect 10332 16270 10334 16322
rect 10386 16270 10388 16322
rect 10332 16258 10388 16270
rect 10444 16716 10668 16772
rect 9548 15934 9550 15986
rect 9602 15934 9604 15986
rect 9548 15922 9604 15934
rect 8652 14308 8708 14318
rect 8016 14140 8280 14150
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8016 14074 8280 14084
rect 8652 13858 8708 14252
rect 8652 13806 8654 13858
rect 8706 13806 8708 13858
rect 8652 13794 8708 13806
rect 8988 13858 9044 14364
rect 8988 13806 8990 13858
rect 9042 13806 9044 13858
rect 7868 13694 7870 13746
rect 7922 13694 7924 13746
rect 7868 13682 7924 13694
rect 8652 13636 8708 13646
rect 7420 13076 7476 13086
rect 7308 13074 7476 13076
rect 7308 13022 7422 13074
rect 7474 13022 7476 13074
rect 7308 13020 7476 13022
rect 7420 13010 7476 13020
rect 4060 12898 4116 12908
rect 5852 12962 5908 12974
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 3052 12850 3108 12862
rect 3052 12798 3054 12850
rect 3106 12798 3108 12850
rect 1820 12086 1876 12124
rect 2044 12738 2100 12750
rect 2044 12686 2046 12738
rect 2098 12686 2100 12738
rect 1820 10610 1876 10622
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 10388 1876 10558
rect 2044 10612 2100 12686
rect 3052 11956 3108 12798
rect 3724 12740 3780 12750
rect 3388 12180 3444 12190
rect 3724 12180 3780 12684
rect 5852 12740 5908 12910
rect 6076 12852 6132 12862
rect 6076 12758 6132 12796
rect 7084 12852 7140 12862
rect 5852 12674 5908 12684
rect 6524 12740 6580 12750
rect 3388 12178 3780 12180
rect 3388 12126 3390 12178
rect 3442 12126 3726 12178
rect 3778 12126 3780 12178
rect 3388 12124 3780 12126
rect 3388 12114 3444 12124
rect 3724 12114 3780 12124
rect 3836 12348 4788 12404
rect 3052 11890 3108 11900
rect 3836 11506 3892 12348
rect 4396 12178 4452 12190
rect 4396 12126 4398 12178
rect 4450 12126 4452 12178
rect 3948 12068 4004 12078
rect 3948 12066 4340 12068
rect 3948 12014 3950 12066
rect 4002 12014 4340 12066
rect 3948 12012 4340 12014
rect 3948 12002 4004 12012
rect 3836 11454 3838 11506
rect 3890 11454 3892 11506
rect 3836 11442 3892 11454
rect 4284 11396 4340 12012
rect 4396 11620 4452 12126
rect 4732 12178 4788 12348
rect 4732 12126 4734 12178
rect 4786 12126 4788 12178
rect 4732 12114 4788 12126
rect 4614 11788 4878 11798
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4614 11722 4878 11732
rect 4396 11554 4452 11564
rect 5628 11396 5684 11406
rect 4284 11340 4564 11396
rect 4508 10834 4564 11340
rect 4956 11284 5012 11294
rect 4956 11282 5348 11284
rect 4956 11230 4958 11282
rect 5010 11230 5348 11282
rect 4956 11228 5348 11230
rect 4956 11218 5012 11228
rect 4508 10782 4510 10834
rect 4562 10782 4564 10834
rect 4508 10770 4564 10782
rect 5292 10834 5348 11228
rect 5292 10782 5294 10834
rect 5346 10782 5348 10834
rect 5292 10770 5348 10782
rect 2156 10612 2212 10622
rect 2044 10610 2212 10612
rect 2044 10558 2158 10610
rect 2210 10558 2212 10610
rect 2044 10556 2212 10558
rect 2156 10546 2212 10556
rect 5628 10610 5684 11340
rect 5628 10558 5630 10610
rect 5682 10558 5684 10610
rect 1820 10322 1876 10332
rect 2492 10388 2548 10398
rect 2380 9716 2436 9726
rect 1596 8148 1652 8158
rect 1596 7698 1652 8092
rect 1596 7646 1598 7698
rect 1650 7646 1652 7698
rect 1596 7634 1652 7646
rect 2380 7698 2436 9660
rect 2492 9042 2548 10332
rect 5628 10388 5684 10558
rect 4614 10220 4878 10230
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4614 10154 4878 10164
rect 5628 9828 5684 10332
rect 5292 9826 5684 9828
rect 5292 9774 5630 9826
rect 5682 9774 5684 9826
rect 5292 9772 5684 9774
rect 4284 9716 4340 9726
rect 4284 9622 4340 9660
rect 4620 9714 4676 9726
rect 4620 9662 4622 9714
rect 4674 9662 4676 9714
rect 4620 9604 4676 9662
rect 5068 9604 5124 9614
rect 4620 9602 5124 9604
rect 4620 9550 5070 9602
rect 5122 9550 5124 9602
rect 4620 9548 5124 9550
rect 2492 8990 2494 9042
rect 2546 8990 2548 9042
rect 2492 8978 2548 8990
rect 2828 9042 2884 9054
rect 2828 8990 2830 9042
rect 2882 8990 2884 9042
rect 2828 8372 2884 8990
rect 4614 8652 4878 8662
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4614 8586 4878 8596
rect 5068 8484 5124 9548
rect 5068 8418 5124 8428
rect 2828 8306 2884 8316
rect 3612 8372 3668 8382
rect 3612 8278 3668 8316
rect 4732 8372 4788 8382
rect 2492 8148 2548 8158
rect 2492 8054 2548 8092
rect 2380 7646 2382 7698
rect 2434 7646 2436 7698
rect 2380 7634 2436 7646
rect 4732 7474 4788 8316
rect 4732 7422 4734 7474
rect 4786 7422 4788 7474
rect 4732 7410 4788 7422
rect 5292 7474 5348 9772
rect 5628 9762 5684 9772
rect 6076 10610 6132 10622
rect 6076 10558 6078 10610
rect 6130 10558 6132 10610
rect 5404 9268 5460 9278
rect 5404 9266 5796 9268
rect 5404 9214 5406 9266
rect 5458 9214 5796 9266
rect 5404 9212 5796 9214
rect 5404 9202 5460 9212
rect 5740 8370 5796 9212
rect 6076 8932 6132 10558
rect 6076 8866 6132 8876
rect 6188 9826 6244 9838
rect 6188 9774 6190 9826
rect 6242 9774 6244 9826
rect 5740 8318 5742 8370
rect 5794 8318 5796 8370
rect 5740 8306 5796 8318
rect 5964 8818 6020 8830
rect 5964 8766 5966 8818
rect 6018 8766 6020 8818
rect 5964 7588 6020 8766
rect 6076 8484 6132 8494
rect 6076 8370 6132 8428
rect 6076 8318 6078 8370
rect 6130 8318 6132 8370
rect 6076 8306 6132 8318
rect 5964 7522 6020 7532
rect 5292 7422 5294 7474
rect 5346 7422 5348 7474
rect 5292 7410 5348 7422
rect 6188 7362 6244 9774
rect 6188 7310 6190 7362
rect 6242 7310 6244 7362
rect 6188 7298 6244 7310
rect 6524 8484 6580 12684
rect 7084 12402 7140 12796
rect 8016 12572 8280 12582
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8016 12506 8280 12516
rect 7084 12350 7086 12402
rect 7138 12350 7140 12402
rect 7084 12338 7140 12350
rect 8652 12290 8708 13580
rect 8988 13636 9044 13806
rect 8988 13570 9044 13580
rect 9324 15428 9380 15438
rect 8764 13524 8820 13534
rect 8764 12850 8820 13468
rect 9324 12962 9380 15372
rect 10444 15428 10500 16716
rect 10668 16706 10724 16716
rect 11116 16882 11172 16894
rect 11116 16830 11118 16882
rect 11170 16830 11172 16882
rect 11116 16660 11172 16830
rect 11116 16594 11172 16604
rect 11418 16492 11682 16502
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11418 16426 11682 16436
rect 12348 16212 12404 17502
rect 13356 16996 13412 17006
rect 12908 16994 13412 16996
rect 12908 16942 13358 16994
rect 13410 16942 13412 16994
rect 12908 16940 13412 16942
rect 12348 16156 12740 16212
rect 12348 15988 12404 15998
rect 12572 15988 12628 15998
rect 12348 15986 12572 15988
rect 12348 15934 12350 15986
rect 12402 15934 12572 15986
rect 12348 15932 12572 15934
rect 12348 15922 12404 15932
rect 12572 15894 12628 15932
rect 9660 14868 9716 14878
rect 9660 14530 9716 14812
rect 9660 14478 9662 14530
rect 9714 14478 9716 14530
rect 9660 14466 9716 14478
rect 10332 14532 10388 14542
rect 10444 14532 10500 15372
rect 11418 14924 11682 14934
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11418 14858 11682 14868
rect 12572 14644 12628 14654
rect 10332 14530 10500 14532
rect 10332 14478 10334 14530
rect 10386 14478 10500 14530
rect 10332 14476 10500 14478
rect 11788 14642 12628 14644
rect 11788 14590 12574 14642
rect 12626 14590 12628 14642
rect 11788 14588 12628 14590
rect 10332 14466 10388 14476
rect 11788 13970 11844 14588
rect 12572 14578 12628 14588
rect 12684 14532 12740 16156
rect 12908 16210 12964 16940
rect 13356 16930 13412 16940
rect 12908 16158 12910 16210
rect 12962 16158 12964 16210
rect 12908 16146 12964 16158
rect 13468 16772 13524 19182
rect 13580 18674 13636 19854
rect 14028 19908 14084 19918
rect 14028 19234 14084 19852
rect 14028 19182 14030 19234
rect 14082 19182 14084 19234
rect 14028 19170 14084 19182
rect 13580 18622 13582 18674
rect 13634 18622 13636 18674
rect 13580 18610 13636 18622
rect 14140 18450 14196 20076
rect 16268 20132 16324 20142
rect 16268 20038 16324 20076
rect 14252 20018 14308 20030
rect 14252 19966 14254 20018
rect 14306 19966 14308 20018
rect 14252 19908 14308 19966
rect 14364 19908 14420 19918
rect 15260 19908 15316 19918
rect 14252 19906 14532 19908
rect 14252 19854 14366 19906
rect 14418 19854 14532 19906
rect 14252 19852 14532 19854
rect 14364 19842 14420 19852
rect 14140 18398 14142 18450
rect 14194 18398 14196 18450
rect 14140 18386 14196 18398
rect 14364 18450 14420 18462
rect 14364 18398 14366 18450
rect 14418 18398 14420 18450
rect 14364 17668 14420 18398
rect 14476 18340 14532 19852
rect 17276 19908 17332 20526
rect 21624 20412 21888 20422
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21624 20346 21888 20356
rect 22764 20242 22820 20748
rect 22988 20738 23044 20748
rect 23660 20802 23716 21420
rect 23660 20750 23662 20802
rect 23714 20750 23716 20802
rect 23660 20738 23716 20750
rect 22764 20190 22766 20242
rect 22818 20190 22820 20242
rect 21644 20132 21700 20142
rect 20748 20130 21700 20132
rect 20748 20078 21646 20130
rect 21698 20078 21700 20130
rect 20748 20076 21700 20078
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 17612 19908 17668 19918
rect 17836 19908 17892 19918
rect 17276 19906 17668 19908
rect 17276 19854 17614 19906
rect 17666 19854 17668 19906
rect 17276 19852 17668 19854
rect 15260 19814 15316 19852
rect 14476 18274 14532 18284
rect 14588 19460 14644 19470
rect 14140 16996 14196 17006
rect 14140 16902 14196 16940
rect 13468 16098 13524 16716
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 12796 15428 12852 15438
rect 12796 15334 12852 15372
rect 13468 15428 13524 16046
rect 14028 16772 14084 16782
rect 14028 16098 14084 16716
rect 14028 16046 14030 16098
rect 14082 16046 14084 16098
rect 14028 16034 14084 16046
rect 13468 15362 13524 15372
rect 14364 15428 14420 17612
rect 14364 15362 14420 15372
rect 14476 15314 14532 15326
rect 14476 15262 14478 15314
rect 14530 15262 14532 15314
rect 12796 14532 12852 14542
rect 12684 14530 12852 14532
rect 12684 14478 12798 14530
rect 12850 14478 12852 14530
rect 12684 14476 12852 14478
rect 11900 14420 11956 14430
rect 11900 14326 11956 14364
rect 12796 14420 12852 14476
rect 12796 14354 12852 14364
rect 13916 14420 13972 14430
rect 13916 14326 13972 14364
rect 11788 13918 11790 13970
rect 11842 13918 11844 13970
rect 11788 13906 11844 13918
rect 12012 14306 12068 14318
rect 12012 14254 12014 14306
rect 12066 14254 12068 14306
rect 11116 13524 11172 13534
rect 11116 13430 11172 13468
rect 11418 13356 11682 13366
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11418 13290 11682 13300
rect 9324 12910 9326 12962
rect 9378 12910 9380 12962
rect 9324 12898 9380 12910
rect 9660 12964 9716 12974
rect 9660 12870 9716 12908
rect 8764 12798 8766 12850
rect 8818 12798 8820 12850
rect 8764 12786 8820 12798
rect 12012 12850 12068 14254
rect 14252 13746 14308 13758
rect 14252 13694 14254 13746
rect 14306 13694 14308 13746
rect 14252 13636 14308 13694
rect 14252 13570 14308 13580
rect 12796 13188 12852 13198
rect 12796 13094 12852 13132
rect 12012 12798 12014 12850
rect 12066 12798 12068 12850
rect 12012 12786 12068 12798
rect 14476 13076 14532 15262
rect 14588 13524 14644 19404
rect 15484 19348 15540 19358
rect 14820 18844 15084 18854
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 14820 18778 15084 18788
rect 15036 18452 15092 18462
rect 15036 17666 15092 18396
rect 15372 18340 15428 18350
rect 15372 18246 15428 18284
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 17602 15092 17614
rect 15484 17666 15540 19292
rect 17052 19124 17108 19134
rect 17052 19030 17108 19068
rect 16268 19010 16324 19022
rect 16268 18958 16270 19010
rect 16322 18958 16324 19010
rect 16268 18562 16324 18958
rect 16268 18510 16270 18562
rect 16322 18510 16324 18562
rect 16268 18498 16324 18510
rect 16044 18450 16100 18462
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18340 16100 18398
rect 17500 18452 17556 18462
rect 17500 18358 17556 18396
rect 16044 18274 16100 18284
rect 16716 18340 16772 18350
rect 15484 17614 15486 17666
rect 15538 17614 15540 17666
rect 15484 17602 15540 17614
rect 16716 17668 16772 18284
rect 16716 17602 16772 17612
rect 17612 17668 17668 19852
rect 17612 17602 17668 17612
rect 17724 19906 17892 19908
rect 17724 19854 17838 19906
rect 17890 19854 17892 19906
rect 17724 19852 17892 19854
rect 17724 17554 17780 19852
rect 17836 19842 17892 19852
rect 18222 19628 18486 19638
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18222 19562 18486 19572
rect 18284 19348 18340 19358
rect 18284 19254 18340 19292
rect 18956 19236 19012 19966
rect 18620 18676 18676 18686
rect 17836 18450 17892 18462
rect 17836 18398 17838 18450
rect 17890 18398 17892 18450
rect 17836 18340 17892 18398
rect 17836 18274 17892 18284
rect 17948 18452 18004 18462
rect 17724 17502 17726 17554
rect 17778 17502 17780 17554
rect 17724 17490 17780 17502
rect 14820 17276 15084 17286
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 14820 17210 15084 17220
rect 17836 17108 17892 17118
rect 17948 17108 18004 18396
rect 18222 18060 18486 18070
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18222 17994 18486 18004
rect 18508 17892 18564 17902
rect 18620 17892 18676 18620
rect 18956 18564 19012 19180
rect 19404 20018 19460 20030
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19292 19124 19348 19134
rect 19292 19030 19348 19068
rect 18956 18498 19012 18508
rect 18508 17890 18676 17892
rect 18508 17838 18510 17890
rect 18562 17838 18676 17890
rect 18508 17836 18676 17838
rect 18508 17826 18564 17836
rect 19404 17780 19460 19966
rect 20188 18564 20244 18574
rect 19404 17714 19460 17724
rect 19852 18562 20244 18564
rect 19852 18510 20190 18562
rect 20242 18510 20244 18562
rect 19852 18508 20244 18510
rect 19852 17778 19908 18508
rect 20188 18498 20244 18508
rect 19852 17726 19854 17778
rect 19906 17726 19908 17778
rect 19852 17714 19908 17726
rect 20748 17778 20804 20076
rect 21644 20066 21700 20076
rect 22428 20132 22484 20142
rect 22428 20038 22484 20076
rect 21868 19908 21924 19918
rect 21420 19236 21476 19246
rect 21308 19180 21420 19236
rect 21308 18674 21364 19180
rect 21420 19142 21476 19180
rect 21868 19234 21924 19852
rect 21868 19182 21870 19234
rect 21922 19182 21924 19234
rect 21868 19170 21924 19182
rect 22764 19236 22820 20190
rect 24892 19458 24948 21644
rect 27244 21700 27300 21710
rect 27244 21606 27300 21644
rect 28140 21588 28196 22988
rect 28252 22932 28308 23660
rect 28428 23548 28692 23558
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28428 23482 28692 23492
rect 28252 22866 28308 22876
rect 28428 21980 28692 21990
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28428 21914 28692 21924
rect 28140 21522 28196 21532
rect 26012 21474 26068 21486
rect 26012 21422 26014 21474
rect 26066 21422 26068 21474
rect 25026 21196 25290 21206
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25026 21130 25290 21140
rect 26012 20188 26068 21422
rect 26236 21476 26292 21486
rect 26236 21382 26292 21420
rect 27468 20860 27860 20916
rect 26124 20692 26180 20702
rect 26124 20578 26180 20636
rect 26908 20692 26964 20702
rect 26908 20598 26964 20636
rect 27244 20690 27300 20702
rect 27244 20638 27246 20690
rect 27298 20638 27300 20690
rect 26124 20526 26126 20578
rect 26178 20526 26180 20578
rect 26124 20514 26180 20526
rect 26684 20578 26740 20590
rect 26684 20526 26686 20578
rect 26738 20526 26740 20578
rect 25564 20132 26068 20188
rect 26684 20188 26740 20526
rect 27244 20468 27300 20638
rect 27468 20468 27524 20860
rect 27804 20804 27860 20860
rect 27804 20802 28196 20804
rect 27804 20750 27806 20802
rect 27858 20750 28196 20802
rect 27804 20748 28196 20750
rect 27804 20738 27860 20748
rect 27244 20412 27524 20468
rect 27580 20690 27636 20702
rect 27580 20638 27582 20690
rect 27634 20638 27636 20690
rect 26684 20132 26964 20188
rect 25026 19628 25290 19638
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25026 19562 25290 19572
rect 24892 19406 24894 19458
rect 24946 19406 24948 19458
rect 24892 19394 24948 19406
rect 21624 18844 21888 18854
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21624 18778 21888 18788
rect 21308 18622 21310 18674
rect 21362 18622 21364 18674
rect 21308 18610 21364 18622
rect 22764 18564 22820 19180
rect 24108 19010 24164 19022
rect 24108 18958 24110 19010
rect 24162 18958 24164 19010
rect 22764 18498 22820 18508
rect 23212 18676 23268 18686
rect 23212 18562 23268 18620
rect 24108 18674 24164 18958
rect 24108 18622 24110 18674
rect 24162 18622 24164 18674
rect 24108 18610 24164 18622
rect 25228 19012 25284 19022
rect 25564 19012 25620 20132
rect 25228 19010 25620 19012
rect 25228 18958 25230 19010
rect 25282 18958 25620 19010
rect 25228 18956 25620 18958
rect 25900 20020 25956 20030
rect 23212 18510 23214 18562
rect 23266 18510 23268 18562
rect 23212 18498 23268 18510
rect 24108 18450 24164 18462
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 22204 18340 22260 18350
rect 22204 18246 22260 18284
rect 24108 18340 24164 18398
rect 24892 18452 24948 18462
rect 24164 18284 24276 18340
rect 24108 18274 24164 18284
rect 20972 18228 21028 18238
rect 20972 18134 21028 18172
rect 23548 18228 23604 18238
rect 20748 17726 20750 17778
rect 20802 17726 20804 17778
rect 20748 17714 20804 17726
rect 22316 17780 22372 17790
rect 22316 17686 22372 17724
rect 18956 17666 19012 17678
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 17836 17106 18004 17108
rect 17836 17054 17838 17106
rect 17890 17054 18004 17106
rect 17836 17052 18004 17054
rect 18732 17554 18788 17566
rect 18732 17502 18734 17554
rect 18786 17502 18788 17554
rect 16380 16996 16436 17006
rect 16380 16902 16436 16940
rect 15372 16772 15428 16782
rect 15372 16678 15428 16716
rect 15708 16772 15764 16782
rect 15708 15988 15764 16716
rect 14820 15708 15084 15718
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 14820 15642 15084 15652
rect 15708 15538 15764 15932
rect 15708 15486 15710 15538
rect 15762 15486 15764 15538
rect 15708 15474 15764 15486
rect 16268 16212 16324 16222
rect 14700 15428 14756 15438
rect 14700 14530 14756 15372
rect 15148 15428 15204 15438
rect 15148 15334 15204 15372
rect 14700 14478 14702 14530
rect 14754 14478 14756 14530
rect 14700 14466 14756 14478
rect 15148 14532 15204 14542
rect 14820 14140 15084 14150
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 14820 14074 15084 14084
rect 15148 13972 15204 14476
rect 15820 14532 15876 14542
rect 15820 14438 15876 14476
rect 16268 14530 16324 16156
rect 17052 15988 17108 15998
rect 17052 15894 17108 15932
rect 16492 15876 16548 15886
rect 16492 15782 16548 15820
rect 16268 14478 16270 14530
rect 16322 14478 16324 14530
rect 16268 14466 16324 14478
rect 17836 15314 17892 17052
rect 18284 16882 18340 16894
rect 18284 16830 18286 16882
rect 18338 16830 18340 16882
rect 18284 16772 18340 16830
rect 18284 16706 18340 16716
rect 18620 16770 18676 16782
rect 18620 16718 18622 16770
rect 18674 16718 18676 16770
rect 18620 16660 18676 16718
rect 18620 16594 18676 16604
rect 18222 16492 18486 16502
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18222 16426 18486 16436
rect 18284 16212 18340 16222
rect 18284 16118 18340 16156
rect 17836 15262 17838 15314
rect 17890 15262 17892 15314
rect 17836 14532 17892 15262
rect 18396 15316 18452 15326
rect 18396 15222 18452 15260
rect 18222 14924 18486 14934
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18222 14858 18486 14868
rect 17836 14466 17892 14476
rect 18732 14306 18788 17502
rect 18956 16884 19012 17614
rect 19628 17668 19684 17678
rect 19628 17574 19684 17612
rect 20524 17668 20580 17678
rect 20524 17574 20580 17612
rect 21420 17668 21476 17678
rect 21420 17574 21476 17612
rect 21868 17668 21924 17678
rect 21868 17574 21924 17612
rect 23548 17554 23604 18172
rect 24220 17780 24276 18284
rect 24892 18228 24948 18396
rect 25228 18228 25284 18956
rect 25900 18340 25956 19964
rect 26236 19908 26292 19918
rect 26236 19814 26292 19852
rect 26684 19348 26740 19358
rect 25900 18274 25956 18284
rect 26124 19346 26740 19348
rect 26124 19294 26686 19346
rect 26738 19294 26740 19346
rect 26124 19292 26740 19294
rect 24892 18172 25284 18228
rect 24220 17778 24500 17780
rect 24220 17726 24222 17778
rect 24274 17726 24500 17778
rect 24220 17724 24500 17726
rect 24220 17668 24276 17724
rect 24220 17602 24276 17612
rect 23548 17502 23550 17554
rect 23602 17502 23604 17554
rect 23548 17490 23604 17502
rect 21624 17276 21888 17286
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21624 17210 21888 17220
rect 23436 17106 23492 17118
rect 23436 17054 23438 17106
rect 23490 17054 23492 17106
rect 19964 16994 20020 17006
rect 19964 16942 19966 16994
rect 20018 16942 20020 16994
rect 18956 16818 19012 16828
rect 19740 16884 19796 16894
rect 19292 15988 19348 15998
rect 19292 15894 19348 15932
rect 19292 15428 19348 15438
rect 19292 14754 19348 15372
rect 19292 14702 19294 14754
rect 19346 14702 19348 14754
rect 19292 14690 19348 14702
rect 18732 14254 18734 14306
rect 18786 14254 18788 14306
rect 18732 14242 18788 14254
rect 19740 14308 19796 16828
rect 19964 15988 20020 16942
rect 23436 16996 23492 17054
rect 24444 17108 24500 17724
rect 23436 16930 23492 16940
rect 24220 16996 24276 17006
rect 24220 16902 24276 16940
rect 20524 16882 20580 16894
rect 20860 16884 20916 16894
rect 20524 16830 20526 16882
rect 20578 16830 20580 16882
rect 20300 16772 20356 16782
rect 20300 16098 20356 16716
rect 20300 16046 20302 16098
rect 20354 16046 20356 16098
rect 20300 16034 20356 16046
rect 19964 15922 20020 15932
rect 20300 15876 20356 15886
rect 20300 15782 20356 15820
rect 20524 15540 20580 16830
rect 20188 15484 20524 15540
rect 20188 14642 20244 15484
rect 20524 15474 20580 15484
rect 20748 16882 20916 16884
rect 20748 16830 20862 16882
rect 20914 16830 20916 16882
rect 20748 16828 20916 16830
rect 20748 15316 20804 16828
rect 20860 16818 20916 16828
rect 24444 16882 24500 17052
rect 24444 16830 24446 16882
rect 24498 16830 24500 16882
rect 24444 16818 24500 16830
rect 24780 17668 24836 17678
rect 24892 17668 24948 18172
rect 25026 18060 25290 18070
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25026 17994 25290 18004
rect 24780 17666 24948 17668
rect 24780 17614 24782 17666
rect 24834 17614 24948 17666
rect 24780 17612 24948 17614
rect 25228 17668 25284 17678
rect 26124 17668 26180 19292
rect 26684 19282 26740 19292
rect 26908 19124 26964 20132
rect 27244 20132 27300 20142
rect 27244 20038 27300 20076
rect 27356 20020 27412 20412
rect 27356 19954 27412 19964
rect 26908 19058 26964 19068
rect 26684 18340 26740 18350
rect 25228 17666 26180 17668
rect 25228 17614 25230 17666
rect 25282 17614 26180 17666
rect 25228 17612 26180 17614
rect 26236 18338 26740 18340
rect 26236 18286 26686 18338
rect 26738 18286 26740 18338
rect 26236 18284 26740 18286
rect 24780 16884 24836 17612
rect 25228 17602 25284 17612
rect 25340 17108 25396 17118
rect 26236 17108 26292 18284
rect 26684 18274 26740 18284
rect 27580 17442 27636 20638
rect 28140 20242 28196 20748
rect 28428 20412 28692 20422
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28428 20346 28692 20356
rect 28140 20190 28142 20242
rect 28194 20190 28196 20242
rect 28140 20178 28196 20190
rect 27692 19124 27748 19134
rect 27692 19030 27748 19068
rect 28428 18844 28692 18854
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28428 18778 28692 18788
rect 28028 18564 28084 18574
rect 28028 18562 28308 18564
rect 28028 18510 28030 18562
rect 28082 18510 28308 18562
rect 28028 18508 28308 18510
rect 28028 18498 28084 18508
rect 28252 17890 28308 18508
rect 28252 17838 28254 17890
rect 28306 17838 28308 17890
rect 28252 17826 28308 17838
rect 27580 17390 27582 17442
rect 27634 17390 27636 17442
rect 27580 17378 27636 17390
rect 28428 17276 28692 17286
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28428 17210 28692 17220
rect 25340 17014 25396 17052
rect 25452 17052 26292 17108
rect 27132 17108 27188 17118
rect 24892 16884 24948 16894
rect 24780 16828 24892 16884
rect 23996 16658 24052 16670
rect 23996 16606 23998 16658
rect 24050 16606 24052 16658
rect 22092 16098 22148 16110
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 21624 15708 21888 15718
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21624 15642 21888 15652
rect 20860 15540 20916 15550
rect 21756 15540 21812 15550
rect 20860 15538 21700 15540
rect 20860 15486 20862 15538
rect 20914 15486 21700 15538
rect 20860 15484 21700 15486
rect 20860 15474 20916 15484
rect 21420 15316 21476 15326
rect 20748 15260 20916 15316
rect 20188 14590 20190 14642
rect 20242 14590 20244 14642
rect 20188 14578 20244 14590
rect 19740 14214 19796 14252
rect 20636 14308 20692 14318
rect 20748 14308 20804 14318
rect 20692 14306 20804 14308
rect 20692 14254 20750 14306
rect 20802 14254 20804 14306
rect 20692 14252 20804 14254
rect 14812 13970 15204 13972
rect 14812 13918 15150 13970
rect 15202 13918 15204 13970
rect 14812 13916 15204 13918
rect 14812 13746 14868 13916
rect 15148 13878 15204 13916
rect 14812 13694 14814 13746
rect 14866 13694 14868 13746
rect 14812 13682 14868 13694
rect 19404 13858 19460 13870
rect 19404 13806 19406 13858
rect 19458 13806 19460 13858
rect 18396 13636 18452 13646
rect 18396 13542 18452 13580
rect 14588 13468 14980 13524
rect 8652 12238 8654 12290
rect 8706 12238 8708 12290
rect 8652 12226 8708 12238
rect 14476 12178 14532 13020
rect 14924 13076 14980 13468
rect 18222 13356 18486 13366
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18222 13290 18486 13300
rect 19404 13188 19460 13806
rect 19404 13122 19460 13132
rect 20300 13746 20356 13758
rect 20300 13694 20302 13746
rect 20354 13694 20356 13746
rect 20076 13076 20132 13086
rect 14924 13074 15204 13076
rect 14924 13022 14926 13074
rect 14978 13022 15204 13074
rect 14924 13020 15204 13022
rect 14924 13010 14980 13020
rect 15148 12962 15204 13020
rect 15148 12910 15150 12962
rect 15202 12910 15204 12962
rect 15148 12898 15204 12910
rect 20076 12850 20132 13020
rect 20076 12798 20078 12850
rect 20130 12798 20132 12850
rect 14820 12572 15084 12582
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 14820 12506 15084 12516
rect 20076 12404 20132 12798
rect 20076 12338 20132 12348
rect 14476 12126 14478 12178
rect 14530 12126 14532 12178
rect 14476 12114 14532 12126
rect 18060 12290 18116 12302
rect 18060 12238 18062 12290
rect 18114 12238 18116 12290
rect 8876 12068 8932 12078
rect 8876 11974 8932 12012
rect 10108 12066 10164 12078
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 7196 11956 7252 11966
rect 7196 11618 7252 11900
rect 7868 11956 7924 11966
rect 7868 11954 8484 11956
rect 7868 11902 7870 11954
rect 7922 11902 8484 11954
rect 7868 11900 8484 11902
rect 7868 11890 7924 11900
rect 8428 11844 8484 11900
rect 8428 11788 8708 11844
rect 7196 11566 7198 11618
rect 7250 11566 7252 11618
rect 7196 11554 7252 11566
rect 7980 11732 8036 11742
rect 7980 11282 8036 11676
rect 7980 11230 7982 11282
rect 8034 11230 8036 11282
rect 7980 11218 8036 11230
rect 8016 11004 8280 11014
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8016 10938 8280 10948
rect 8316 10836 8372 10846
rect 8316 10742 8372 10780
rect 8540 9602 8596 9614
rect 8540 9550 8542 9602
rect 8594 9550 8596 9602
rect 8016 9436 8280 9446
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8016 9370 8280 9380
rect 7532 8932 7588 8942
rect 7532 8838 7588 8876
rect 6524 8034 6580 8428
rect 7420 8372 7476 8382
rect 7420 8278 7476 8316
rect 6524 7982 6526 8034
rect 6578 7982 6580 8034
rect 4614 7084 4878 7094
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4614 7018 4878 7028
rect 6524 6692 6580 7982
rect 8016 7868 8280 7878
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8016 7802 8280 7812
rect 8540 7700 8596 9550
rect 8652 8146 8708 11788
rect 10108 11732 10164 12014
rect 17276 11954 17332 11966
rect 17276 11902 17278 11954
rect 17330 11902 17332 11954
rect 11418 11788 11682 11798
rect 10108 11666 10164 11676
rect 10668 11732 10724 11742
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11418 11722 11682 11732
rect 10332 11396 10388 11406
rect 10332 11302 10388 11340
rect 10668 11394 10724 11676
rect 10668 11342 10670 11394
rect 10722 11342 10724 11394
rect 10108 11172 10164 11182
rect 9884 10724 9940 10734
rect 9324 10722 9940 10724
rect 9324 10670 9886 10722
rect 9938 10670 9940 10722
rect 9324 10668 9940 10670
rect 9100 10388 9156 10398
rect 9100 10386 9268 10388
rect 9100 10334 9102 10386
rect 9154 10334 9268 10386
rect 9100 10332 9268 10334
rect 9100 10322 9156 10332
rect 9212 9828 9268 10332
rect 9324 10050 9380 10668
rect 9884 10658 9940 10668
rect 9324 9998 9326 10050
rect 9378 9998 9380 10050
rect 9324 9986 9380 9998
rect 9212 9772 9828 9828
rect 9212 9604 9268 9614
rect 8876 9602 9268 9604
rect 8876 9550 9214 9602
rect 9266 9550 9268 9602
rect 8876 9548 9268 9550
rect 8876 9154 8932 9548
rect 9212 9538 9268 9548
rect 8876 9102 8878 9154
rect 8930 9102 8932 9154
rect 8876 9090 8932 9102
rect 9324 9156 9380 9166
rect 9324 8370 9380 9100
rect 9324 8318 9326 8370
rect 9378 8318 9380 8370
rect 9324 8306 9380 8318
rect 8652 8094 8654 8146
rect 8706 8094 8708 8146
rect 8652 8082 8708 8094
rect 8204 7644 8596 7700
rect 7196 7588 7252 7598
rect 7196 7494 7252 7532
rect 6524 6626 6580 6636
rect 7980 6692 8036 6702
rect 7980 6598 8036 6636
rect 8204 6690 8260 7644
rect 9772 7586 9828 9772
rect 10108 9714 10164 11116
rect 10668 10612 10724 11342
rect 14588 11396 14644 11406
rect 11116 11282 11172 11294
rect 11116 11230 11118 11282
rect 11170 11230 11172 11282
rect 11116 10836 11172 11230
rect 11452 11282 11508 11294
rect 11452 11230 11454 11282
rect 11506 11230 11508 11282
rect 11452 10948 11508 11230
rect 11900 11282 11956 11294
rect 11900 11230 11902 11282
rect 11954 11230 11956 11282
rect 11900 11172 11956 11230
rect 12236 11282 12292 11294
rect 12236 11230 12238 11282
rect 12290 11230 12292 11282
rect 12236 11172 12292 11230
rect 12684 11172 12740 11182
rect 11900 11106 11956 11116
rect 12012 11170 12964 11172
rect 12012 11118 12686 11170
rect 12738 11118 12964 11170
rect 12012 11116 12964 11118
rect 12012 10948 12068 11116
rect 12684 11106 12740 11116
rect 11452 10892 12068 10948
rect 11116 10770 11172 10780
rect 11676 10834 11732 10892
rect 11676 10782 11678 10834
rect 11730 10782 11732 10834
rect 11676 10770 11732 10782
rect 10668 10546 10724 10556
rect 12460 10612 12516 10622
rect 12516 10556 12852 10612
rect 12460 10518 12516 10556
rect 11228 10500 11284 10510
rect 11228 10406 11284 10444
rect 11418 10220 11682 10230
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11418 10154 11682 10164
rect 10108 9662 10110 9714
rect 10162 9662 10164 9714
rect 10108 9650 10164 9662
rect 11116 9828 11172 9838
rect 10108 9156 10164 9166
rect 10108 9062 10164 9100
rect 10108 8036 10164 8046
rect 10108 7942 10164 7980
rect 9772 7534 9774 7586
rect 9826 7534 9828 7586
rect 9772 7522 9828 7534
rect 11116 7362 11172 9772
rect 12348 9828 12404 9838
rect 12348 9734 12404 9772
rect 12796 9826 12852 10556
rect 12908 10164 12964 11116
rect 13020 10610 13076 10622
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 13020 10500 13076 10558
rect 13020 10434 13076 10444
rect 12908 10098 12964 10108
rect 12796 9774 12798 9826
rect 12850 9774 12852 9826
rect 11452 9044 11508 9054
rect 11452 8930 11508 8988
rect 11452 8878 11454 8930
rect 11506 8878 11508 8930
rect 11452 8866 11508 8878
rect 12796 9042 12852 9774
rect 12796 8990 12798 9042
rect 12850 8990 12852 9042
rect 11418 8652 11682 8662
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11418 8586 11682 8596
rect 12460 8260 12516 8298
rect 12460 8194 12516 8204
rect 12796 8258 12852 8990
rect 13244 9044 13300 9054
rect 13244 8950 13300 8988
rect 12796 8206 12798 8258
rect 12850 8206 12852 8258
rect 12796 8194 12852 8206
rect 14140 8258 14196 8270
rect 14140 8206 14142 8258
rect 14194 8206 14196 8258
rect 12460 8036 12516 8046
rect 12460 7586 12516 7980
rect 14140 8036 14196 8206
rect 14140 7970 14196 7980
rect 14476 8260 14532 8270
rect 12460 7534 12462 7586
rect 12514 7534 12516 7586
rect 12460 7522 12516 7534
rect 11116 7310 11118 7362
rect 11170 7310 11172 7362
rect 11116 7298 11172 7310
rect 12684 7474 12740 7486
rect 12684 7422 12686 7474
rect 12738 7422 12740 7474
rect 12684 7364 12740 7422
rect 13244 7364 13300 7374
rect 12684 7308 13244 7364
rect 11418 7084 11682 7094
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11418 7018 11682 7028
rect 12684 6804 12740 7308
rect 13244 7270 13300 7308
rect 12684 6738 12740 6748
rect 14476 6802 14532 8204
rect 14588 7364 14644 11340
rect 15708 11394 15764 11406
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 14820 11004 15084 11014
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 14820 10938 15084 10948
rect 15596 10836 15652 10846
rect 15596 10742 15652 10780
rect 15148 10164 15204 10174
rect 14820 9436 15084 9446
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 14820 9370 15084 9380
rect 15148 8370 15204 10108
rect 15708 9826 15764 11342
rect 16156 11396 16212 11406
rect 16156 11394 16324 11396
rect 16156 11342 16158 11394
rect 16210 11342 16324 11394
rect 16156 11340 16324 11342
rect 16156 11330 16212 11340
rect 16156 10388 16212 10398
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15148 8318 15150 8370
rect 15202 8318 15204 8370
rect 14820 7868 15084 7878
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 14820 7802 15084 7812
rect 14924 7364 14980 7374
rect 14588 7362 14980 7364
rect 14588 7310 14926 7362
rect 14978 7310 14980 7362
rect 14588 7308 14980 7310
rect 14924 7298 14980 7308
rect 15148 7364 15204 8318
rect 14476 6750 14478 6802
rect 14530 6750 14532 6802
rect 14476 6738 14532 6750
rect 8204 6638 8206 6690
rect 8258 6638 8260 6690
rect 8204 6626 8260 6638
rect 8652 6692 8708 6702
rect 8652 6598 8708 6636
rect 8016 6300 8280 6310
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8016 6234 8280 6244
rect 14820 6300 15084 6310
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 14820 6234 15084 6244
rect 14812 6132 14868 6142
rect 15148 6132 15204 7308
rect 14812 6130 15204 6132
rect 14812 6078 14814 6130
rect 14866 6078 15204 6130
rect 14812 6076 15204 6078
rect 14812 6066 14868 6076
rect 13804 6020 13860 6030
rect 13804 6018 14308 6020
rect 13804 5966 13806 6018
rect 13858 5966 14308 6018
rect 13804 5964 14308 5966
rect 13804 5954 13860 5964
rect 12572 5908 12628 5918
rect 4614 5516 4878 5526
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4614 5450 4878 5460
rect 11418 5516 11682 5526
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11418 5450 11682 5460
rect 8016 4732 8280 4742
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8016 4666 8280 4676
rect 4614 3948 4878 3958
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4614 3882 4878 3892
rect 11418 3948 11682 3958
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11418 3882 11682 3892
rect 12236 3444 12292 3454
rect 12124 3442 12516 3444
rect 12124 3390 12238 3442
rect 12290 3390 12516 3442
rect 12124 3388 12516 3390
rect 8016 3164 8280 3174
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8016 3098 8280 3108
rect 12124 800 12180 3388
rect 12236 3378 12292 3388
rect 12460 3220 12516 3388
rect 12572 3442 12628 5852
rect 13468 5908 13524 5918
rect 13468 5814 13524 5852
rect 14140 4450 14196 4462
rect 14140 4398 14142 4450
rect 14194 4398 14196 4450
rect 12572 3390 12574 3442
rect 12626 3390 12628 3442
rect 12572 3378 12628 3390
rect 12796 4226 12852 4238
rect 12796 4174 12798 4226
rect 12850 4174 12852 4226
rect 12796 3220 12852 4174
rect 13132 3332 13188 3342
rect 13580 3332 13636 3342
rect 12460 3164 12852 3220
rect 12908 3330 13188 3332
rect 12908 3278 13134 3330
rect 13186 3278 13188 3330
rect 12908 3276 13188 3278
rect 12908 1652 12964 3276
rect 13132 3266 13188 3276
rect 13468 3330 13636 3332
rect 13468 3278 13582 3330
rect 13634 3278 13636 3330
rect 13468 3276 13636 3278
rect 12796 1596 12964 1652
rect 12796 800 12852 1596
rect 13468 800 13524 3276
rect 13580 3266 13636 3276
rect 14140 800 14196 4398
rect 14252 3554 14308 5964
rect 15148 6018 15204 6076
rect 15596 9154 15652 9166
rect 15596 9102 15598 9154
rect 15650 9102 15652 9154
rect 15148 5966 15150 6018
rect 15202 5966 15204 6018
rect 15148 5954 15204 5966
rect 15484 6020 15540 6030
rect 15596 6020 15652 9102
rect 15708 9044 15764 9774
rect 15708 8978 15764 8988
rect 15820 10386 16212 10388
rect 15820 10334 16158 10386
rect 16210 10334 16212 10386
rect 15820 10332 16212 10334
rect 15820 6578 15876 10332
rect 16156 10322 16212 10332
rect 16268 10052 16324 11340
rect 16380 10836 16436 10846
rect 16380 10722 16436 10780
rect 16380 10670 16382 10722
rect 16434 10670 16436 10722
rect 16380 10658 16436 10670
rect 16716 10500 16772 10510
rect 16716 10406 16772 10444
rect 16268 9986 16324 9996
rect 16156 9826 16212 9838
rect 16156 9774 16158 9826
rect 16210 9774 16212 9826
rect 16156 8372 16212 9774
rect 16156 8306 16212 8316
rect 16380 8818 16436 8830
rect 16380 8766 16382 8818
rect 16434 8766 16436 8818
rect 16380 8148 16436 8766
rect 16380 8082 16436 8092
rect 16828 8036 16884 8046
rect 16828 7942 16884 7980
rect 16268 7588 16324 7598
rect 16268 7494 16324 7532
rect 17276 7588 17332 11902
rect 18060 11508 18116 12238
rect 19628 12180 19684 12190
rect 18222 11788 18486 11798
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18222 11722 18486 11732
rect 18060 11442 18116 11452
rect 19180 11396 19236 11406
rect 19180 11302 19236 11340
rect 18620 11284 18676 11294
rect 18620 11170 18676 11228
rect 19404 11284 19460 11294
rect 19404 11190 19460 11228
rect 18620 11118 18622 11170
rect 18674 11118 18676 11170
rect 18620 11106 18676 11118
rect 17500 10500 17556 10510
rect 17500 10406 17556 10444
rect 19292 10500 19348 10510
rect 19628 10500 19684 12124
rect 20300 12180 20356 13694
rect 20300 12114 20356 12124
rect 20412 12292 20468 12302
rect 20412 12178 20468 12236
rect 20412 12126 20414 12178
rect 20466 12126 20468 12178
rect 20412 12114 20468 12126
rect 20636 11956 20692 14252
rect 20748 14242 20804 14252
rect 20748 13746 20804 13758
rect 20748 13694 20750 13746
rect 20802 13694 20804 13746
rect 20748 13636 20804 13694
rect 20748 13570 20804 13580
rect 20412 11900 20692 11956
rect 20188 11508 20244 11518
rect 19740 11284 19796 11294
rect 20076 11284 20132 11294
rect 19740 11282 20132 11284
rect 19740 11230 19742 11282
rect 19794 11230 20078 11282
rect 20130 11230 20132 11282
rect 19740 11228 20132 11230
rect 19740 11218 19796 11228
rect 19964 10610 20020 10622
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19740 10500 19796 10510
rect 19964 10500 20020 10558
rect 19292 10498 20020 10500
rect 19292 10446 19294 10498
rect 19346 10446 19742 10498
rect 19794 10446 20020 10498
rect 19292 10444 20020 10446
rect 18222 10220 18486 10230
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18222 10154 18486 10164
rect 18620 9716 18676 9726
rect 18620 9602 18676 9660
rect 18620 9550 18622 9602
rect 18674 9550 18676 9602
rect 18620 9538 18676 9550
rect 19180 9604 19236 9614
rect 19180 9510 19236 9548
rect 17500 9044 17556 9054
rect 17500 8950 17556 8988
rect 18172 9042 18228 9054
rect 18172 8990 18174 9042
rect 18226 8990 18228 9042
rect 18172 8932 18228 8990
rect 19292 9044 19348 10444
rect 19740 10434 19796 10444
rect 19740 9940 19796 9950
rect 20076 9940 20132 11228
rect 20188 11170 20244 11452
rect 20188 11118 20190 11170
rect 20242 11118 20244 11170
rect 20188 11106 20244 11118
rect 20300 9940 20356 9950
rect 20076 9884 20300 9940
rect 19740 9846 19796 9884
rect 20300 9826 20356 9884
rect 20300 9774 20302 9826
rect 20354 9774 20356 9826
rect 20300 9762 20356 9774
rect 19404 9716 19460 9726
rect 19404 9622 19460 9660
rect 19292 8978 19348 8988
rect 18172 8866 18228 8876
rect 18222 8652 18486 8662
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18222 8586 18486 8596
rect 17612 8372 17668 8382
rect 17612 8278 17668 8316
rect 18620 8148 18676 8158
rect 18620 8054 18676 8092
rect 20412 8036 20468 11900
rect 20636 10610 20692 10622
rect 20636 10558 20638 10610
rect 20690 10558 20692 10610
rect 20524 9714 20580 9726
rect 20524 9662 20526 9714
rect 20578 9662 20580 9714
rect 20524 9266 20580 9662
rect 20524 9214 20526 9266
rect 20578 9214 20580 9266
rect 20524 9202 20580 9214
rect 20636 9268 20692 10558
rect 20860 10500 20916 15260
rect 21420 15222 21476 15260
rect 21644 14642 21700 15484
rect 21644 14590 21646 14642
rect 21698 14590 21700 14642
rect 21644 14578 21700 14590
rect 21756 14308 21812 15484
rect 21420 14252 21812 14308
rect 21868 14530 21924 14542
rect 21868 14478 21870 14530
rect 21922 14478 21924 14530
rect 21868 14308 21924 14478
rect 21420 13076 21476 14252
rect 21868 14242 21924 14252
rect 21624 14140 21888 14150
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21624 14074 21888 14084
rect 20972 13074 21476 13076
rect 20972 13022 21422 13074
rect 21474 13022 21476 13074
rect 20972 13020 21476 13022
rect 20972 12178 21028 13020
rect 21420 13010 21476 13020
rect 21624 12572 21888 12582
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21624 12506 21888 12516
rect 21868 12404 21924 12414
rect 22092 12404 22148 16046
rect 23212 15988 23268 15998
rect 22316 15202 22372 15214
rect 22316 15150 22318 15202
rect 22370 15150 22372 15202
rect 22316 14420 22372 15150
rect 22652 15204 22708 15214
rect 22652 15110 22708 15148
rect 23212 14754 23268 15932
rect 23660 15428 23716 15438
rect 23660 15334 23716 15372
rect 23996 15428 24052 16606
rect 23996 15362 24052 15372
rect 24892 15986 24948 16828
rect 25026 16492 25290 16502
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25026 16426 25290 16436
rect 24892 15934 24894 15986
rect 24946 15934 24948 15986
rect 24892 15540 24948 15934
rect 23212 14702 23214 14754
rect 23266 14702 23268 14754
rect 23212 14690 23268 14702
rect 23772 14756 23828 14766
rect 22652 14420 22708 14430
rect 22316 14418 22708 14420
rect 22316 14366 22654 14418
rect 22706 14366 22708 14418
rect 22316 14364 22708 14366
rect 22316 14308 22372 14364
rect 22316 14242 22372 14252
rect 22652 13972 22708 14364
rect 22652 13906 22708 13916
rect 22988 14418 23044 14430
rect 22988 14366 22990 14418
rect 23042 14366 23044 14418
rect 22988 13970 23044 14366
rect 22988 13918 22990 13970
rect 23042 13918 23044 13970
rect 22988 13906 23044 13918
rect 23772 13970 23828 14700
rect 24892 14532 24948 15484
rect 25340 15428 25396 15438
rect 25340 15334 25396 15372
rect 25026 14924 25290 14934
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25026 14858 25290 14868
rect 23996 14308 24052 14318
rect 23996 14214 24052 14252
rect 23772 13918 23774 13970
rect 23826 13918 23828 13970
rect 23772 13906 23828 13918
rect 24220 13634 24276 13646
rect 24220 13582 24222 13634
rect 24274 13582 24276 13634
rect 23436 13188 23492 13198
rect 21924 12348 22148 12404
rect 22764 12962 22820 12974
rect 22764 12910 22766 12962
rect 22818 12910 22820 12962
rect 20972 12126 20974 12178
rect 21026 12126 21028 12178
rect 20972 12114 21028 12126
rect 21084 12180 21140 12190
rect 21644 12180 21700 12190
rect 21084 12086 21140 12124
rect 21196 12178 21700 12180
rect 21196 12126 21646 12178
rect 21698 12126 21700 12178
rect 21196 12124 21700 12126
rect 20860 10434 20916 10444
rect 21196 9492 21252 12124
rect 21644 12114 21700 12124
rect 21868 11394 21924 12348
rect 21868 11342 21870 11394
rect 21922 11342 21924 11394
rect 21868 11330 21924 11342
rect 21980 12180 22036 12190
rect 21624 11004 21888 11014
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21624 10938 21888 10948
rect 21532 9826 21588 9838
rect 21532 9774 21534 9826
rect 21586 9774 21588 9826
rect 21532 9604 21588 9774
rect 21420 9548 21588 9604
rect 21196 9436 21364 9492
rect 20636 9202 20692 9212
rect 21196 8818 21252 8830
rect 21196 8766 21198 8818
rect 21250 8766 21252 8818
rect 21196 8148 21252 8766
rect 21196 8082 21252 8092
rect 20412 7970 20468 7980
rect 17276 7522 17332 7532
rect 21084 7250 21140 7262
rect 21084 7198 21086 7250
rect 21138 7198 21140 7250
rect 18222 7084 18486 7094
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18222 7018 18486 7028
rect 20524 6692 20580 6702
rect 15820 6526 15822 6578
rect 15874 6526 15876 6578
rect 15820 6514 15876 6526
rect 18844 6580 18900 6590
rect 15484 6018 15652 6020
rect 15484 5966 15486 6018
rect 15538 5966 15652 6018
rect 15484 5964 15652 5966
rect 15484 5954 15540 5964
rect 18222 5516 18486 5526
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18222 5450 18486 5460
rect 14820 4732 15084 4742
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 14820 4666 15084 4676
rect 14924 4452 14980 4462
rect 14924 4450 15204 4452
rect 14924 4398 14926 4450
rect 14978 4398 15204 4450
rect 14924 4396 15204 4398
rect 14924 4386 14980 4396
rect 14700 4340 14756 4350
rect 14700 4246 14756 4284
rect 14252 3502 14254 3554
rect 14306 3502 14308 3554
rect 14252 3490 14308 3502
rect 15148 3554 15204 4396
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3490 15204 3502
rect 15260 4450 15316 4462
rect 18060 4452 18116 4462
rect 15260 4398 15262 4450
rect 15314 4398 15316 4450
rect 15260 3332 15316 4398
rect 17500 4450 18116 4452
rect 17500 4398 18062 4450
rect 18114 4398 18116 4450
rect 17500 4396 18116 4398
rect 16940 4340 16996 4350
rect 15596 3666 15652 3678
rect 15596 3614 15598 3666
rect 15650 3614 15652 3666
rect 15596 3388 15652 3614
rect 15148 3276 15316 3332
rect 15484 3332 15652 3388
rect 16492 3556 16548 3566
rect 16492 3442 16548 3500
rect 16492 3390 16494 3442
rect 16546 3390 16548 3442
rect 14820 3164 15084 3174
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 14820 3098 15084 3108
rect 15148 2996 15204 3276
rect 14812 2940 15204 2996
rect 14812 800 14868 2940
rect 15484 800 15540 3332
rect 16492 2212 16548 3390
rect 16940 3442 16996 4284
rect 17164 3556 17220 3566
rect 17164 3462 17220 3500
rect 16940 3390 16942 3442
rect 16994 3390 16996 3442
rect 16940 3378 16996 3390
rect 16156 2156 16548 2212
rect 16156 800 16212 2156
rect 16828 1762 16884 1774
rect 16828 1710 16830 1762
rect 16882 1710 16884 1762
rect 16828 800 16884 1710
rect 17500 800 17556 4396
rect 18060 4386 18116 4396
rect 18732 4228 18788 4238
rect 18620 4226 18788 4228
rect 18620 4174 18734 4226
rect 18786 4174 18788 4226
rect 18620 4172 18788 4174
rect 18222 3948 18486 3958
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18222 3882 18486 3892
rect 18508 3556 18564 3566
rect 18620 3556 18676 4172
rect 18732 4162 18788 4172
rect 18508 3554 18676 3556
rect 18508 3502 18510 3554
rect 18562 3502 18676 3554
rect 18508 3500 18676 3502
rect 17612 3330 17668 3342
rect 17612 3278 17614 3330
rect 17666 3278 17668 3330
rect 17612 1762 17668 3278
rect 18508 2772 18564 3500
rect 18844 3388 18900 6524
rect 19628 6468 19684 6478
rect 19404 6020 19460 6030
rect 19404 5122 19460 5964
rect 19404 5070 19406 5122
rect 19458 5070 19460 5122
rect 19404 5058 19460 5070
rect 19628 5010 19684 6412
rect 19628 4958 19630 5010
rect 19682 4958 19684 5010
rect 19628 4946 19684 4958
rect 19964 5010 20020 5022
rect 19964 4958 19966 5010
rect 20018 4958 20020 5010
rect 19292 4452 19348 4462
rect 19292 4358 19348 4396
rect 18732 3332 18900 3388
rect 19068 4338 19124 4350
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 3442 19124 4286
rect 19740 4228 19796 4238
rect 19068 3390 19070 3442
rect 19122 3390 19124 3442
rect 19068 3378 19124 3390
rect 19404 4226 19796 4228
rect 19404 4174 19742 4226
rect 19794 4174 19796 4226
rect 19404 4172 19796 4174
rect 19404 3554 19460 4172
rect 19740 4162 19796 4172
rect 19404 3502 19406 3554
rect 19458 3502 19460 3554
rect 19404 3388 19460 3502
rect 19292 3332 19460 3388
rect 19516 3668 19572 3678
rect 18732 3330 18788 3332
rect 18732 3278 18734 3330
rect 18786 3278 18788 3330
rect 18732 3266 18788 3278
rect 18508 2706 18564 2716
rect 19292 2548 19348 3332
rect 17612 1710 17614 1762
rect 17666 1710 17668 1762
rect 17612 1698 17668 1710
rect 18844 2492 19348 2548
rect 18844 800 18900 2492
rect 19516 800 19572 3612
rect 19852 3444 19908 3454
rect 19964 3444 20020 4958
rect 20300 4898 20356 4910
rect 20300 4846 20302 4898
rect 20354 4846 20356 4898
rect 20076 3556 20132 3566
rect 20188 3556 20244 3566
rect 20076 3554 20188 3556
rect 20076 3502 20078 3554
rect 20130 3502 20188 3554
rect 20076 3500 20188 3502
rect 20076 3490 20132 3500
rect 19852 3442 20020 3444
rect 19852 3390 19854 3442
rect 19906 3390 20020 3442
rect 19852 3388 20020 3390
rect 19852 3378 19908 3388
rect 20188 800 20244 3500
rect 20300 3444 20356 4846
rect 20524 4340 20580 6636
rect 20860 6020 20916 6030
rect 20860 5926 20916 5964
rect 21084 6020 21140 7198
rect 21084 5954 21140 5964
rect 21196 5906 21252 5918
rect 21196 5854 21198 5906
rect 21250 5854 21252 5906
rect 20636 5796 20692 5806
rect 21196 5796 21252 5854
rect 20636 5794 21252 5796
rect 20636 5742 20638 5794
rect 20690 5742 21252 5794
rect 20636 5740 21252 5742
rect 20636 5730 20692 5740
rect 21084 5684 21140 5740
rect 21084 5618 21140 5628
rect 21308 5460 21364 9436
rect 21420 8932 21476 9548
rect 21624 9436 21888 9446
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21624 9370 21888 9380
rect 21980 9266 22036 12124
rect 22764 12180 22820 12910
rect 23436 12962 23492 13132
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12898 23492 12910
rect 23996 12290 24052 12302
rect 23996 12238 23998 12290
rect 24050 12238 24052 12290
rect 22764 12114 22820 12124
rect 23548 12180 23604 12190
rect 23548 11508 23604 12124
rect 23996 11732 24052 12238
rect 23996 11666 24052 11676
rect 24220 12068 24276 13582
rect 24220 11508 24276 12012
rect 23548 11506 24276 11508
rect 23548 11454 23550 11506
rect 23602 11454 24276 11506
rect 23548 11452 24276 11454
rect 24780 11954 24836 11966
rect 24780 11902 24782 11954
rect 24834 11902 24836 11954
rect 23548 11442 23604 11452
rect 23100 10834 23156 10846
rect 23100 10782 23102 10834
rect 23154 10782 23156 10834
rect 21980 9214 21982 9266
rect 22034 9214 22036 9266
rect 21980 9202 22036 9214
rect 22316 9268 22372 9278
rect 21980 9044 22036 9054
rect 21532 8932 21588 8942
rect 21420 8930 21588 8932
rect 21420 8878 21534 8930
rect 21586 8878 21588 8930
rect 21420 8876 21588 8878
rect 21532 8036 21588 8876
rect 21532 7970 21588 7980
rect 21624 7868 21888 7878
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21624 7802 21888 7812
rect 21868 7700 21924 7710
rect 21980 7700 22036 8988
rect 22316 8370 22372 9212
rect 23100 9268 23156 10782
rect 23996 10834 24052 11452
rect 23996 10782 23998 10834
rect 24050 10782 24052 10834
rect 23660 10388 23716 10398
rect 23660 10294 23716 10332
rect 23548 9940 23604 9950
rect 23548 9846 23604 9884
rect 23100 9202 23156 9212
rect 23548 9604 23604 9614
rect 23548 9154 23604 9548
rect 23548 9102 23550 9154
rect 23602 9102 23604 9154
rect 23548 9090 23604 9102
rect 22428 8932 22484 8942
rect 22428 8838 22484 8876
rect 22316 8318 22318 8370
rect 22370 8318 22372 8370
rect 22316 8306 22372 8318
rect 23996 8260 24052 10782
rect 24556 10612 24612 10622
rect 24444 10556 24556 10612
rect 24332 10498 24388 10510
rect 24332 10446 24334 10498
rect 24386 10446 24388 10498
rect 24220 9268 24276 9278
rect 24220 9154 24276 9212
rect 24220 9102 24222 9154
rect 24274 9102 24276 9154
rect 24220 9090 24276 9102
rect 24332 9044 24388 10446
rect 24332 8978 24388 8988
rect 24444 9940 24500 10556
rect 24556 10518 24612 10556
rect 24780 10052 24836 11902
rect 24444 9042 24500 9884
rect 24444 8990 24446 9042
rect 24498 8990 24500 9042
rect 24444 8820 24500 8990
rect 23548 8148 23604 8158
rect 23548 8054 23604 8092
rect 21868 7698 22036 7700
rect 21868 7646 21870 7698
rect 21922 7646 22036 7698
rect 21868 7644 22036 7646
rect 21868 7634 21924 7644
rect 21532 6692 21588 6702
rect 21588 6636 21700 6692
rect 21532 6626 21588 6636
rect 21644 6578 21700 6636
rect 23996 6690 24052 8204
rect 24332 8764 24500 8820
rect 24668 9996 24836 10052
rect 24220 7474 24276 7486
rect 24220 7422 24222 7474
rect 24274 7422 24276 7474
rect 24220 7364 24276 7422
rect 24220 7298 24276 7308
rect 23996 6638 23998 6690
rect 24050 6638 24052 6690
rect 23996 6626 24052 6638
rect 24332 6692 24388 8764
rect 24668 8428 24724 9996
rect 24780 9828 24836 9838
rect 24892 9828 24948 14476
rect 25026 13356 25290 13366
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25026 13290 25290 13300
rect 25340 12068 25396 12078
rect 25340 11974 25396 12012
rect 25026 11788 25290 11798
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25026 11722 25290 11732
rect 25026 10220 25290 10230
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25026 10154 25290 10164
rect 24780 9826 24948 9828
rect 24780 9774 24782 9826
rect 24834 9774 24948 9826
rect 24780 9772 24948 9774
rect 25228 9828 25284 9838
rect 25452 9828 25508 17052
rect 25788 16884 25844 16894
rect 25788 16790 25844 16828
rect 26236 16772 26292 16782
rect 26124 16770 26292 16772
rect 26124 16718 26238 16770
rect 26290 16718 26292 16770
rect 26124 16716 26292 16718
rect 25900 13972 25956 13982
rect 25900 13878 25956 13916
rect 26124 13188 26180 16716
rect 26236 16706 26292 16716
rect 27132 15538 27188 17052
rect 27132 15486 27134 15538
rect 27186 15486 27188 15538
rect 26460 15204 26516 15214
rect 26348 15202 26516 15204
rect 26348 15150 26462 15202
rect 26514 15150 26516 15202
rect 26348 15148 26516 15150
rect 26348 14530 26404 15148
rect 26460 15138 26516 15148
rect 27132 14642 27188 15486
rect 27244 16994 27300 17006
rect 27244 16942 27246 16994
rect 27298 16942 27300 16994
rect 27244 14756 27300 16942
rect 28140 16884 28196 16894
rect 28140 16790 28196 16828
rect 27692 16210 27748 16222
rect 27692 16158 27694 16210
rect 27746 16158 27748 16210
rect 27244 14690 27300 14700
rect 27468 15316 27524 15326
rect 27132 14590 27134 14642
rect 27186 14590 27188 14642
rect 27132 14578 27188 14590
rect 26348 14478 26350 14530
rect 26402 14478 26404 14530
rect 26348 14466 26404 14478
rect 26684 14532 26740 14542
rect 26684 14438 26740 14476
rect 27244 14306 27300 14318
rect 27244 14254 27246 14306
rect 27298 14254 27300 14306
rect 26908 14196 26964 14206
rect 26236 13636 26292 13646
rect 26236 13542 26292 13580
rect 26124 13122 26180 13132
rect 26908 13524 26964 14140
rect 27244 14084 27300 14254
rect 26684 12964 26740 12974
rect 25900 12962 26740 12964
rect 25900 12910 26686 12962
rect 26738 12910 26740 12962
rect 25900 12908 26740 12910
rect 25900 12738 25956 12908
rect 26684 12898 26740 12908
rect 26908 12962 26964 13468
rect 26908 12910 26910 12962
rect 26962 12910 26964 12962
rect 26908 12898 26964 12910
rect 27132 14028 27300 14084
rect 25900 12686 25902 12738
rect 25954 12686 25956 12738
rect 25900 12674 25956 12686
rect 26460 12740 26516 12750
rect 26460 12738 26628 12740
rect 26460 12686 26462 12738
rect 26514 12686 26628 12738
rect 26460 12684 26628 12686
rect 26460 12674 26516 12684
rect 26572 12628 26628 12684
rect 26796 12684 26964 12740
rect 26796 12628 26852 12684
rect 26572 12572 26852 12628
rect 26236 12292 26292 12302
rect 25900 12068 25956 12078
rect 25900 11974 25956 12012
rect 26236 12066 26292 12236
rect 26236 12014 26238 12066
rect 26290 12014 26292 12066
rect 26236 12002 26292 12014
rect 26796 11172 26852 11182
rect 26236 10500 26292 10510
rect 26236 10406 26292 10444
rect 25228 9826 25508 9828
rect 25228 9774 25230 9826
rect 25282 9774 25508 9826
rect 25228 9772 25508 9774
rect 26236 10052 26292 10062
rect 24780 9268 24836 9772
rect 25228 9762 25284 9772
rect 24780 9202 24836 9212
rect 26236 8930 26292 9996
rect 26236 8878 26238 8930
rect 26290 8878 26292 8930
rect 26236 8866 26292 8878
rect 25026 8652 25290 8662
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25026 8586 25290 8596
rect 24668 8372 24948 8428
rect 24556 8260 24612 8270
rect 24556 7700 24612 8204
rect 24556 7474 24612 7644
rect 24556 7422 24558 7474
rect 24610 7422 24612 7474
rect 24332 6626 24388 6636
rect 24444 6690 24500 6702
rect 24444 6638 24446 6690
rect 24498 6638 24500 6690
rect 21644 6526 21646 6578
rect 21698 6526 21700 6578
rect 21644 6514 21700 6526
rect 21980 6580 22036 6590
rect 21980 6486 22036 6524
rect 22316 6468 22372 6478
rect 22316 6374 22372 6412
rect 23100 6466 23156 6478
rect 23100 6414 23102 6466
rect 23154 6414 23156 6466
rect 21624 6300 21888 6310
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21624 6234 21888 6244
rect 23100 6132 23156 6414
rect 23100 6066 23156 6076
rect 22540 6020 22596 6030
rect 22540 5926 22596 5964
rect 21084 5404 21364 5460
rect 21532 5794 21588 5806
rect 21532 5742 21534 5794
rect 21586 5742 21588 5794
rect 21084 4564 21140 5404
rect 21532 5348 21588 5742
rect 21084 4498 21140 4508
rect 21196 5292 21588 5348
rect 24332 5794 24388 5806
rect 24332 5742 24334 5794
rect 24386 5742 24388 5794
rect 20748 4340 20804 4350
rect 20524 4338 20804 4340
rect 20524 4286 20750 4338
rect 20802 4286 20804 4338
rect 20524 4284 20804 4286
rect 20748 4274 20804 4284
rect 21196 4340 21252 5292
rect 23324 5236 23380 5246
rect 23324 5142 23380 5180
rect 21196 4274 21252 4284
rect 21308 5124 21364 5134
rect 21308 4338 21364 5068
rect 22316 5012 22372 5022
rect 22316 4918 22372 4956
rect 21532 4900 21588 4910
rect 21308 4286 21310 4338
rect 21362 4286 21364 4338
rect 21308 4274 21364 4286
rect 21420 4898 21588 4900
rect 21420 4846 21534 4898
rect 21586 4846 21588 4898
rect 21420 4844 21588 4846
rect 20412 4228 20468 4238
rect 20412 4134 20468 4172
rect 21420 4116 21476 4844
rect 21532 4834 21588 4844
rect 21624 4732 21888 4742
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21624 4666 21888 4676
rect 24220 4564 24276 4574
rect 24332 4564 24388 5742
rect 24444 4900 24500 6638
rect 24556 5124 24612 7422
rect 24668 6692 24724 6702
rect 24668 6018 24724 6636
rect 24668 5966 24670 6018
rect 24722 5966 24724 6018
rect 24668 5954 24724 5966
rect 24556 5030 24612 5068
rect 24444 4834 24500 4844
rect 24780 5012 24836 5022
rect 24220 4562 24388 4564
rect 24220 4510 24222 4562
rect 24274 4510 24388 4562
rect 24220 4508 24388 4510
rect 24780 4562 24836 4956
rect 24780 4510 24782 4562
rect 24834 4510 24836 4562
rect 24220 4498 24276 4508
rect 24780 4498 24836 4510
rect 22652 4452 22708 4462
rect 21644 4340 21700 4350
rect 21644 4246 21700 4284
rect 21420 4060 21700 4116
rect 20300 3378 20356 3388
rect 20860 3612 21252 3668
rect 20860 800 20916 3612
rect 21196 3556 21252 3612
rect 21532 3666 21588 3678
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3556 21588 3614
rect 21196 3500 21588 3556
rect 21084 3444 21140 3482
rect 21644 3388 21700 4060
rect 22316 3556 22372 3566
rect 22316 3462 22372 3500
rect 22652 3554 22708 4396
rect 24892 4452 24948 8372
rect 25228 8260 25284 8270
rect 25228 8258 25508 8260
rect 25228 8206 25230 8258
rect 25282 8206 25508 8258
rect 25228 8204 25508 8206
rect 25228 8194 25284 8204
rect 25340 7700 25396 7710
rect 25340 7606 25396 7644
rect 25026 7084 25290 7094
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25026 7018 25290 7028
rect 25452 5796 25508 8204
rect 26348 7700 26404 7710
rect 26236 7364 26292 7374
rect 26236 7270 26292 7308
rect 26348 6130 26404 7644
rect 26796 6466 26852 11116
rect 26908 8428 26964 12684
rect 27020 11508 27076 11518
rect 27020 11414 27076 11452
rect 27020 10388 27076 10398
rect 27132 10388 27188 14028
rect 27468 13858 27524 15260
rect 27580 15202 27636 15214
rect 27580 15150 27582 15202
rect 27634 15150 27636 15202
rect 27580 14532 27636 15150
rect 27692 14868 27748 16158
rect 28140 15876 28196 15886
rect 28140 15874 28308 15876
rect 28140 15822 28142 15874
rect 28194 15822 28308 15874
rect 28140 15820 28308 15822
rect 28140 15810 28196 15820
rect 27692 14802 27748 14812
rect 28028 15202 28084 15214
rect 28028 15150 28030 15202
rect 28082 15150 28084 15202
rect 27580 14466 27636 14476
rect 28028 14530 28084 15150
rect 28028 14478 28030 14530
rect 28082 14478 28084 14530
rect 27804 14418 27860 14430
rect 27804 14366 27806 14418
rect 27858 14366 27860 14418
rect 27804 14308 27860 14366
rect 27804 14242 27860 14252
rect 28028 14196 28084 14478
rect 28084 14140 28196 14196
rect 28028 14130 28084 14140
rect 27468 13806 27470 13858
rect 27522 13806 27524 13858
rect 27468 13794 27524 13806
rect 27356 13524 27412 13534
rect 27356 13074 27412 13468
rect 27356 13022 27358 13074
rect 27410 13022 27412 13074
rect 27356 13010 27412 13022
rect 28140 13074 28196 14140
rect 28140 13022 28142 13074
rect 28194 13022 28196 13074
rect 28140 13010 28196 13022
rect 27468 12738 27524 12750
rect 27468 12686 27470 12738
rect 27522 12686 27524 12738
rect 27244 12290 27300 12302
rect 27244 12238 27246 12290
rect 27298 12238 27300 12290
rect 27244 11508 27300 12238
rect 27244 11442 27300 11452
rect 27244 11284 27300 11294
rect 27244 10612 27300 11228
rect 27244 10546 27300 10556
rect 27468 10500 27524 12686
rect 28140 12180 28196 12190
rect 27580 11284 27636 11294
rect 27580 11190 27636 11228
rect 27692 11172 27748 11182
rect 27692 11078 27748 11116
rect 28140 10834 28196 12124
rect 28140 10782 28142 10834
rect 28194 10782 28196 10834
rect 28140 10770 28196 10782
rect 27580 10724 27636 10734
rect 27580 10722 28084 10724
rect 27580 10670 27582 10722
rect 27634 10670 28084 10722
rect 27580 10668 28084 10670
rect 27580 10658 27636 10668
rect 27468 10444 27748 10500
rect 27132 10332 27524 10388
rect 27020 9380 27076 10332
rect 27468 9714 27524 10332
rect 27468 9662 27470 9714
rect 27522 9662 27524 9714
rect 27468 9650 27524 9662
rect 27020 9324 27300 9380
rect 26908 8372 27076 8428
rect 26796 6414 26798 6466
rect 26850 6414 26852 6466
rect 26796 6402 26852 6414
rect 26348 6078 26350 6130
rect 26402 6078 26404 6130
rect 26348 6066 26404 6078
rect 27020 6020 27076 8372
rect 27244 7586 27300 9324
rect 27244 7534 27246 7586
rect 27298 7534 27300 7586
rect 27244 7522 27300 7534
rect 27468 9154 27524 9166
rect 27468 9102 27470 9154
rect 27522 9102 27524 9154
rect 27468 6690 27524 9102
rect 27692 8034 27748 10444
rect 28028 10164 28084 10668
rect 28252 10276 28308 15820
rect 28428 15708 28692 15718
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28428 15642 28692 15652
rect 28428 14140 28692 14150
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28428 14074 28692 14084
rect 28428 12572 28692 12582
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28428 12506 28692 12516
rect 28428 11004 28692 11014
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28428 10938 28692 10948
rect 28252 10220 28420 10276
rect 28028 10108 28308 10164
rect 28252 10050 28308 10108
rect 28252 9998 28254 10050
rect 28306 9998 28308 10050
rect 28252 9986 28308 9998
rect 28364 9828 28420 10220
rect 28252 9772 28420 9828
rect 28140 9268 28196 9278
rect 28140 9174 28196 9212
rect 28252 8370 28308 9772
rect 28428 9436 28692 9446
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28428 9370 28692 9380
rect 28252 8318 28254 8370
rect 28306 8318 28308 8370
rect 28252 8306 28308 8318
rect 27692 7982 27694 8034
rect 27746 7982 27748 8034
rect 27692 7970 27748 7982
rect 28428 7868 28692 7878
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28428 7802 28692 7812
rect 28140 7586 28196 7598
rect 28140 7534 28142 7586
rect 28194 7534 28196 7586
rect 27468 6638 27470 6690
rect 27522 6638 27524 6690
rect 27468 6626 27524 6638
rect 27692 6692 27748 6702
rect 27692 6598 27748 6636
rect 27804 6466 27860 6478
rect 27804 6414 27806 6466
rect 27858 6414 27860 6466
rect 27692 6020 27748 6030
rect 27020 6018 27748 6020
rect 27020 5966 27694 6018
rect 27746 5966 27748 6018
rect 27020 5964 27748 5966
rect 27692 5954 27748 5964
rect 26684 5796 26740 5806
rect 25452 5794 26740 5796
rect 25452 5742 26686 5794
rect 26738 5742 26740 5794
rect 25452 5740 26740 5742
rect 26684 5730 26740 5740
rect 25026 5516 25290 5526
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25026 5450 25290 5460
rect 25228 5236 25284 5246
rect 25228 5122 25284 5180
rect 25228 5070 25230 5122
rect 25282 5070 25284 5122
rect 25228 5058 25284 5070
rect 25340 5124 25396 5134
rect 25340 4564 25396 5068
rect 26236 4900 26292 4910
rect 25900 4564 25956 4574
rect 25340 4562 25956 4564
rect 25340 4510 25342 4562
rect 25394 4510 25902 4562
rect 25954 4510 25956 4562
rect 25340 4508 25956 4510
rect 25340 4498 25396 4508
rect 25900 4498 25956 4508
rect 26124 4564 26180 4574
rect 24892 4386 24948 4396
rect 25026 3948 25290 3958
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25026 3882 25290 3892
rect 23100 3668 23156 3678
rect 23100 3574 23156 3612
rect 26124 3666 26180 4508
rect 26236 4226 26292 4844
rect 27692 4900 27748 4910
rect 27804 4900 27860 6414
rect 28140 6132 28196 7534
rect 28428 6300 28692 6310
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28428 6234 28692 6244
rect 28140 6076 28532 6132
rect 28252 4900 28308 4910
rect 27692 4898 27860 4900
rect 27692 4846 27694 4898
rect 27746 4846 27860 4898
rect 27692 4844 27860 4846
rect 27916 4898 28308 4900
rect 27916 4846 28254 4898
rect 28306 4846 28308 4898
rect 27916 4844 28308 4846
rect 27692 4834 27748 4844
rect 27244 4452 27300 4462
rect 27244 4358 27300 4396
rect 26236 4174 26238 4226
rect 26290 4174 26292 4226
rect 26236 4162 26292 4174
rect 27916 4116 27972 4844
rect 28252 4834 28308 4844
rect 28476 4900 28532 6076
rect 28476 4834 28532 4844
rect 28428 4732 28692 4742
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28428 4666 28692 4676
rect 26124 3614 26126 3666
rect 26178 3614 26180 3666
rect 26124 3602 26180 3614
rect 27468 4060 27972 4116
rect 28140 4450 28196 4462
rect 28140 4398 28142 4450
rect 28194 4398 28196 4450
rect 22652 3502 22654 3554
rect 22706 3502 22708 3554
rect 22652 3490 22708 3502
rect 21084 3378 21140 3388
rect 21420 3332 21700 3388
rect 27468 3442 27524 4060
rect 27468 3390 27470 3442
rect 27522 3390 27524 3442
rect 27468 3378 27524 3390
rect 28140 3444 28196 4398
rect 28140 3378 28196 3388
rect 24780 3332 24836 3342
rect 21420 2436 21476 3332
rect 24780 3330 24948 3332
rect 24780 3278 24782 3330
rect 24834 3278 24948 3330
rect 24780 3276 24948 3278
rect 24780 3266 24836 3276
rect 21624 3164 21888 3174
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21624 3098 21888 3108
rect 21420 2380 21588 2436
rect 21532 800 21588 2380
rect 24892 800 24948 3276
rect 28428 3164 28692 3174
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28428 3098 28692 3108
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
<< via2 >>
rect 8016 26682 8072 26684
rect 8016 26630 8018 26682
rect 8018 26630 8070 26682
rect 8070 26630 8072 26682
rect 8016 26628 8072 26630
rect 8120 26682 8176 26684
rect 8120 26630 8122 26682
rect 8122 26630 8174 26682
rect 8174 26630 8176 26682
rect 8120 26628 8176 26630
rect 8224 26682 8280 26684
rect 8224 26630 8226 26682
rect 8226 26630 8278 26682
rect 8278 26630 8280 26682
rect 8224 26628 8280 26630
rect 4614 25898 4670 25900
rect 4614 25846 4616 25898
rect 4616 25846 4668 25898
rect 4668 25846 4670 25898
rect 4614 25844 4670 25846
rect 4718 25898 4774 25900
rect 4718 25846 4720 25898
rect 4720 25846 4772 25898
rect 4772 25846 4774 25898
rect 4718 25844 4774 25846
rect 4822 25898 4878 25900
rect 4822 25846 4824 25898
rect 4824 25846 4876 25898
rect 4876 25846 4878 25898
rect 4822 25844 4878 25846
rect 1708 25282 1764 25284
rect 1708 25230 1710 25282
rect 1710 25230 1762 25282
rect 1762 25230 1764 25282
rect 1708 25228 1764 25230
rect 8016 25114 8072 25116
rect 8016 25062 8018 25114
rect 8018 25062 8070 25114
rect 8070 25062 8072 25114
rect 8016 25060 8072 25062
rect 8120 25114 8176 25116
rect 8120 25062 8122 25114
rect 8122 25062 8174 25114
rect 8174 25062 8176 25114
rect 8120 25060 8176 25062
rect 8224 25114 8280 25116
rect 8224 25062 8226 25114
rect 8226 25062 8278 25114
rect 8278 25062 8280 25114
rect 8224 25060 8280 25062
rect 4614 24330 4670 24332
rect 4614 24278 4616 24330
rect 4616 24278 4668 24330
rect 4668 24278 4670 24330
rect 4614 24276 4670 24278
rect 4718 24330 4774 24332
rect 4718 24278 4720 24330
rect 4720 24278 4772 24330
rect 4772 24278 4774 24330
rect 4718 24276 4774 24278
rect 4822 24330 4878 24332
rect 4822 24278 4824 24330
rect 4824 24278 4876 24330
rect 4876 24278 4878 24330
rect 4822 24276 4878 24278
rect 9548 25228 9604 25284
rect 11418 25898 11474 25900
rect 11418 25846 11420 25898
rect 11420 25846 11472 25898
rect 11472 25846 11474 25898
rect 11418 25844 11474 25846
rect 11522 25898 11578 25900
rect 11522 25846 11524 25898
rect 11524 25846 11576 25898
rect 11576 25846 11578 25898
rect 11522 25844 11578 25846
rect 11626 25898 11682 25900
rect 11626 25846 11628 25898
rect 11628 25846 11680 25898
rect 11680 25846 11682 25898
rect 11626 25844 11682 25846
rect 13356 26514 13412 26516
rect 13356 26462 13358 26514
rect 13358 26462 13410 26514
rect 13410 26462 13412 26514
rect 13356 26460 13412 26462
rect 14028 26460 14084 26516
rect 12796 25676 12852 25732
rect 12908 26236 12964 26292
rect 13692 26290 13748 26292
rect 13692 26238 13694 26290
rect 13694 26238 13746 26290
rect 13746 26238 13748 26290
rect 13692 26236 13748 26238
rect 14820 26682 14876 26684
rect 14820 26630 14822 26682
rect 14822 26630 14874 26682
rect 14874 26630 14876 26682
rect 14820 26628 14876 26630
rect 14924 26682 14980 26684
rect 14924 26630 14926 26682
rect 14926 26630 14978 26682
rect 14978 26630 14980 26682
rect 14924 26628 14980 26630
rect 15028 26682 15084 26684
rect 15028 26630 15030 26682
rect 15030 26630 15082 26682
rect 15082 26630 15084 26682
rect 15028 26628 15084 26630
rect 13916 25676 13972 25732
rect 10332 25228 10388 25284
rect 11340 25282 11396 25284
rect 11340 25230 11342 25282
rect 11342 25230 11394 25282
rect 11394 25230 11396 25282
rect 11340 25228 11396 25230
rect 12796 25228 12852 25284
rect 14820 25114 14876 25116
rect 14820 25062 14822 25114
rect 14822 25062 14874 25114
rect 14874 25062 14876 25114
rect 14820 25060 14876 25062
rect 14924 25114 14980 25116
rect 14924 25062 14926 25114
rect 14926 25062 14978 25114
rect 14978 25062 14980 25114
rect 14924 25060 14980 25062
rect 15028 25114 15084 25116
rect 15028 25062 15030 25114
rect 15030 25062 15082 25114
rect 15082 25062 15084 25114
rect 15028 25060 15084 25062
rect 11418 24330 11474 24332
rect 11418 24278 11420 24330
rect 11420 24278 11472 24330
rect 11472 24278 11474 24330
rect 11418 24276 11474 24278
rect 11522 24330 11578 24332
rect 11522 24278 11524 24330
rect 11524 24278 11576 24330
rect 11576 24278 11578 24330
rect 11522 24276 11578 24278
rect 11626 24330 11682 24332
rect 11626 24278 11628 24330
rect 11628 24278 11680 24330
rect 11680 24278 11682 24330
rect 11626 24276 11682 24278
rect 8016 23546 8072 23548
rect 8016 23494 8018 23546
rect 8018 23494 8070 23546
rect 8070 23494 8072 23546
rect 8016 23492 8072 23494
rect 8120 23546 8176 23548
rect 8120 23494 8122 23546
rect 8122 23494 8174 23546
rect 8174 23494 8176 23546
rect 8120 23492 8176 23494
rect 8224 23546 8280 23548
rect 8224 23494 8226 23546
rect 8226 23494 8278 23546
rect 8278 23494 8280 23546
rect 8224 23492 8280 23494
rect 14820 23546 14876 23548
rect 14820 23494 14822 23546
rect 14822 23494 14874 23546
rect 14874 23494 14876 23546
rect 14820 23492 14876 23494
rect 14924 23546 14980 23548
rect 14924 23494 14926 23546
rect 14926 23494 14978 23546
rect 14978 23494 14980 23546
rect 14924 23492 14980 23494
rect 15028 23546 15084 23548
rect 15028 23494 15030 23546
rect 15030 23494 15082 23546
rect 15082 23494 15084 23546
rect 15028 23492 15084 23494
rect 4614 22762 4670 22764
rect 4614 22710 4616 22762
rect 4616 22710 4668 22762
rect 4668 22710 4670 22762
rect 4614 22708 4670 22710
rect 4718 22762 4774 22764
rect 4718 22710 4720 22762
rect 4720 22710 4772 22762
rect 4772 22710 4774 22762
rect 4718 22708 4774 22710
rect 4822 22762 4878 22764
rect 4822 22710 4824 22762
rect 4824 22710 4876 22762
rect 4876 22710 4878 22762
rect 4822 22708 4878 22710
rect 11418 22762 11474 22764
rect 11418 22710 11420 22762
rect 11420 22710 11472 22762
rect 11472 22710 11474 22762
rect 11418 22708 11474 22710
rect 11522 22762 11578 22764
rect 11522 22710 11524 22762
rect 11524 22710 11576 22762
rect 11576 22710 11578 22762
rect 11522 22708 11578 22710
rect 11626 22762 11682 22764
rect 11626 22710 11628 22762
rect 11628 22710 11680 22762
rect 11680 22710 11682 22762
rect 11626 22708 11682 22710
rect 8016 21978 8072 21980
rect 8016 21926 8018 21978
rect 8018 21926 8070 21978
rect 8070 21926 8072 21978
rect 8016 21924 8072 21926
rect 8120 21978 8176 21980
rect 8120 21926 8122 21978
rect 8122 21926 8174 21978
rect 8174 21926 8176 21978
rect 8120 21924 8176 21926
rect 8224 21978 8280 21980
rect 8224 21926 8226 21978
rect 8226 21926 8278 21978
rect 8278 21926 8280 21978
rect 8224 21924 8280 21926
rect 14820 21978 14876 21980
rect 14820 21926 14822 21978
rect 14822 21926 14874 21978
rect 14874 21926 14876 21978
rect 14820 21924 14876 21926
rect 14924 21978 14980 21980
rect 14924 21926 14926 21978
rect 14926 21926 14978 21978
rect 14978 21926 14980 21978
rect 14924 21924 14980 21926
rect 15028 21978 15084 21980
rect 15028 21926 15030 21978
rect 15030 21926 15082 21978
rect 15082 21926 15084 21978
rect 15028 21924 15084 21926
rect 15708 21810 15764 21812
rect 15708 21758 15710 21810
rect 15710 21758 15762 21810
rect 15762 21758 15764 21810
rect 15708 21756 15764 21758
rect 16268 26290 16324 26292
rect 16268 26238 16270 26290
rect 16270 26238 16322 26290
rect 16322 26238 16324 26290
rect 16268 26236 16324 26238
rect 16492 25564 16548 25620
rect 17164 26236 17220 26292
rect 18172 26796 18228 26852
rect 18956 26796 19012 26852
rect 17612 26460 17668 26516
rect 18222 25898 18278 25900
rect 18222 25846 18224 25898
rect 18224 25846 18276 25898
rect 18276 25846 18278 25898
rect 18222 25844 18278 25846
rect 18326 25898 18382 25900
rect 18326 25846 18328 25898
rect 18328 25846 18380 25898
rect 18380 25846 18382 25898
rect 18326 25844 18382 25846
rect 18430 25898 18486 25900
rect 18430 25846 18432 25898
rect 18432 25846 18484 25898
rect 18484 25846 18486 25898
rect 18430 25844 18486 25846
rect 18222 24330 18278 24332
rect 18222 24278 18224 24330
rect 18224 24278 18276 24330
rect 18276 24278 18278 24330
rect 18222 24276 18278 24278
rect 18326 24330 18382 24332
rect 18326 24278 18328 24330
rect 18328 24278 18380 24330
rect 18380 24278 18382 24330
rect 18326 24276 18382 24278
rect 18430 24330 18486 24332
rect 18430 24278 18432 24330
rect 18432 24278 18484 24330
rect 18484 24278 18486 24330
rect 18430 24276 18486 24278
rect 18222 22762 18278 22764
rect 18222 22710 18224 22762
rect 18224 22710 18276 22762
rect 18276 22710 18278 22762
rect 18222 22708 18278 22710
rect 18326 22762 18382 22764
rect 18326 22710 18328 22762
rect 18328 22710 18380 22762
rect 18380 22710 18382 22762
rect 18326 22708 18382 22710
rect 18430 22762 18486 22764
rect 18430 22710 18432 22762
rect 18432 22710 18484 22762
rect 18484 22710 18486 22762
rect 18430 22708 18486 22710
rect 18620 21756 18676 21812
rect 16380 21698 16436 21700
rect 16380 21646 16382 21698
rect 16382 21646 16434 21698
rect 16434 21646 16436 21698
rect 16380 21644 16436 21646
rect 19068 26460 19124 26516
rect 19516 26460 19572 26516
rect 19628 25452 19684 25508
rect 20188 25506 20244 25508
rect 20188 25454 20190 25506
rect 20190 25454 20242 25506
rect 20242 25454 20244 25506
rect 20188 25452 20244 25454
rect 19068 25340 19124 25396
rect 18956 25228 19012 25284
rect 21532 26796 21588 26852
rect 22764 26796 22820 26852
rect 21624 26682 21680 26684
rect 21624 26630 21626 26682
rect 21626 26630 21678 26682
rect 21678 26630 21680 26682
rect 21624 26628 21680 26630
rect 21728 26682 21784 26684
rect 21728 26630 21730 26682
rect 21730 26630 21782 26682
rect 21782 26630 21784 26682
rect 21728 26628 21784 26630
rect 21832 26682 21888 26684
rect 21832 26630 21834 26682
rect 21834 26630 21886 26682
rect 21886 26630 21888 26682
rect 21832 26628 21888 26630
rect 21196 26460 21252 26516
rect 20860 25452 20916 25508
rect 21308 25452 21364 25508
rect 20748 25340 20804 25396
rect 19964 25282 20020 25284
rect 19964 25230 19966 25282
rect 19966 25230 20018 25282
rect 20018 25230 20020 25282
rect 19964 25228 20020 25230
rect 22876 26460 22932 26516
rect 22652 25564 22708 25620
rect 22204 25506 22260 25508
rect 22204 25454 22206 25506
rect 22206 25454 22258 25506
rect 22258 25454 22260 25506
rect 22204 25452 22260 25454
rect 23884 26514 23940 26516
rect 23884 26462 23886 26514
rect 23886 26462 23938 26514
rect 23938 26462 23940 26514
rect 23884 26460 23940 26462
rect 28140 26796 28196 26852
rect 26236 26236 26292 26292
rect 25026 25898 25082 25900
rect 25026 25846 25028 25898
rect 25028 25846 25080 25898
rect 25080 25846 25082 25898
rect 25026 25844 25082 25846
rect 25130 25898 25186 25900
rect 25130 25846 25132 25898
rect 25132 25846 25184 25898
rect 25184 25846 25186 25898
rect 25130 25844 25186 25846
rect 25234 25898 25290 25900
rect 25234 25846 25236 25898
rect 25236 25846 25288 25898
rect 25288 25846 25290 25898
rect 25234 25844 25290 25846
rect 21420 25228 21476 25284
rect 21980 25282 22036 25284
rect 21980 25230 21982 25282
rect 21982 25230 22034 25282
rect 22034 25230 22036 25282
rect 21980 25228 22036 25230
rect 21624 25114 21680 25116
rect 21624 25062 21626 25114
rect 21626 25062 21678 25114
rect 21678 25062 21680 25114
rect 21624 25060 21680 25062
rect 21728 25114 21784 25116
rect 21728 25062 21730 25114
rect 21730 25062 21782 25114
rect 21782 25062 21784 25114
rect 21728 25060 21784 25062
rect 21832 25114 21888 25116
rect 21832 25062 21834 25114
rect 21834 25062 21886 25114
rect 21886 25062 21888 25114
rect 21832 25060 21888 25062
rect 27692 25564 27748 25620
rect 27132 25506 27188 25508
rect 27132 25454 27134 25506
rect 27134 25454 27186 25506
rect 27186 25454 27188 25506
rect 27132 25452 27188 25454
rect 28428 26682 28484 26684
rect 28428 26630 28430 26682
rect 28430 26630 28482 26682
rect 28482 26630 28484 26682
rect 28428 26628 28484 26630
rect 28532 26682 28588 26684
rect 28532 26630 28534 26682
rect 28534 26630 28586 26682
rect 28586 26630 28588 26682
rect 28532 26628 28588 26630
rect 28636 26682 28692 26684
rect 28636 26630 28638 26682
rect 28638 26630 28690 26682
rect 28690 26630 28692 26682
rect 28636 26628 28692 26630
rect 28140 25506 28196 25508
rect 28140 25454 28142 25506
rect 28142 25454 28194 25506
rect 28194 25454 28196 25506
rect 28140 25452 28196 25454
rect 27468 25282 27524 25284
rect 27468 25230 27470 25282
rect 27470 25230 27522 25282
rect 27522 25230 27524 25282
rect 27468 25228 27524 25230
rect 28428 25114 28484 25116
rect 28428 25062 28430 25114
rect 28430 25062 28482 25114
rect 28482 25062 28484 25114
rect 28428 25060 28484 25062
rect 28532 25114 28588 25116
rect 28532 25062 28534 25114
rect 28534 25062 28586 25114
rect 28586 25062 28588 25114
rect 28532 25060 28588 25062
rect 28636 25114 28692 25116
rect 28636 25062 28638 25114
rect 28638 25062 28690 25114
rect 28690 25062 28692 25114
rect 28636 25060 28692 25062
rect 25026 24330 25082 24332
rect 25026 24278 25028 24330
rect 25028 24278 25080 24330
rect 25080 24278 25082 24330
rect 25026 24276 25082 24278
rect 25130 24330 25186 24332
rect 25130 24278 25132 24330
rect 25132 24278 25184 24330
rect 25184 24278 25186 24330
rect 25130 24276 25186 24278
rect 25234 24330 25290 24332
rect 25234 24278 25236 24330
rect 25236 24278 25288 24330
rect 25288 24278 25290 24330
rect 25234 24276 25290 24278
rect 28140 24220 28196 24276
rect 27692 23714 27748 23716
rect 27692 23662 27694 23714
rect 27694 23662 27746 23714
rect 27746 23662 27748 23714
rect 27692 23660 27748 23662
rect 21624 23546 21680 23548
rect 21624 23494 21626 23546
rect 21626 23494 21678 23546
rect 21678 23494 21680 23546
rect 21624 23492 21680 23494
rect 21728 23546 21784 23548
rect 21728 23494 21730 23546
rect 21730 23494 21782 23546
rect 21782 23494 21784 23546
rect 21728 23492 21784 23494
rect 21832 23546 21888 23548
rect 21832 23494 21834 23546
rect 21834 23494 21886 23546
rect 21886 23494 21888 23546
rect 21832 23492 21888 23494
rect 26908 23042 26964 23044
rect 26908 22990 26910 23042
rect 26910 22990 26962 23042
rect 26962 22990 26964 23042
rect 26908 22988 26964 22990
rect 25026 22762 25082 22764
rect 25026 22710 25028 22762
rect 25028 22710 25080 22762
rect 25080 22710 25082 22762
rect 25026 22708 25082 22710
rect 25130 22762 25186 22764
rect 25130 22710 25132 22762
rect 25132 22710 25184 22762
rect 25184 22710 25186 22762
rect 25130 22708 25186 22710
rect 25234 22762 25290 22764
rect 25234 22710 25236 22762
rect 25236 22710 25288 22762
rect 25288 22710 25290 22762
rect 25234 22708 25290 22710
rect 28140 22988 28196 23044
rect 28028 22258 28084 22260
rect 28028 22206 28030 22258
rect 28030 22206 28082 22258
rect 28082 22206 28084 22258
rect 28028 22204 28084 22206
rect 21624 21978 21680 21980
rect 21624 21926 21626 21978
rect 21626 21926 21678 21978
rect 21678 21926 21680 21978
rect 21624 21924 21680 21926
rect 21728 21978 21784 21980
rect 21728 21926 21730 21978
rect 21730 21926 21782 21978
rect 21782 21926 21784 21978
rect 21728 21924 21784 21926
rect 21832 21978 21888 21980
rect 21832 21926 21834 21978
rect 21834 21926 21886 21978
rect 21886 21926 21888 21978
rect 21832 21924 21888 21926
rect 18732 21644 18788 21700
rect 24892 21644 24948 21700
rect 23660 21420 23716 21476
rect 4614 21194 4670 21196
rect 4614 21142 4616 21194
rect 4616 21142 4668 21194
rect 4668 21142 4670 21194
rect 4614 21140 4670 21142
rect 4718 21194 4774 21196
rect 4718 21142 4720 21194
rect 4720 21142 4772 21194
rect 4772 21142 4774 21194
rect 4718 21140 4774 21142
rect 4822 21194 4878 21196
rect 4822 21142 4824 21194
rect 4824 21142 4876 21194
rect 4876 21142 4878 21194
rect 4822 21140 4878 21142
rect 11418 21194 11474 21196
rect 11418 21142 11420 21194
rect 11420 21142 11472 21194
rect 11472 21142 11474 21194
rect 11418 21140 11474 21142
rect 11522 21194 11578 21196
rect 11522 21142 11524 21194
rect 11524 21142 11576 21194
rect 11576 21142 11578 21194
rect 11522 21140 11578 21142
rect 11626 21194 11682 21196
rect 11626 21142 11628 21194
rect 11628 21142 11680 21194
rect 11680 21142 11682 21194
rect 11626 21140 11682 21142
rect 18222 21194 18278 21196
rect 18222 21142 18224 21194
rect 18224 21142 18276 21194
rect 18276 21142 18278 21194
rect 18222 21140 18278 21142
rect 18326 21194 18382 21196
rect 18326 21142 18328 21194
rect 18328 21142 18380 21194
rect 18380 21142 18382 21194
rect 18326 21140 18382 21142
rect 18430 21194 18486 21196
rect 18430 21142 18432 21194
rect 18432 21142 18484 21194
rect 18484 21142 18486 21194
rect 18430 21140 18486 21142
rect 8016 20410 8072 20412
rect 8016 20358 8018 20410
rect 8018 20358 8070 20410
rect 8070 20358 8072 20410
rect 8016 20356 8072 20358
rect 8120 20410 8176 20412
rect 8120 20358 8122 20410
rect 8122 20358 8174 20410
rect 8174 20358 8176 20410
rect 8120 20356 8176 20358
rect 8224 20410 8280 20412
rect 8224 20358 8226 20410
rect 8226 20358 8278 20410
rect 8278 20358 8280 20410
rect 8224 20356 8280 20358
rect 14820 20410 14876 20412
rect 14820 20358 14822 20410
rect 14822 20358 14874 20410
rect 14874 20358 14876 20410
rect 14820 20356 14876 20358
rect 14924 20410 14980 20412
rect 14924 20358 14926 20410
rect 14926 20358 14978 20410
rect 14978 20358 14980 20410
rect 14924 20356 14980 20358
rect 15028 20410 15084 20412
rect 15028 20358 15030 20410
rect 15030 20358 15082 20410
rect 15082 20358 15084 20410
rect 15028 20356 15084 20358
rect 8764 19852 8820 19908
rect 4614 19626 4670 19628
rect 4614 19574 4616 19626
rect 4616 19574 4668 19626
rect 4668 19574 4670 19626
rect 4614 19572 4670 19574
rect 4718 19626 4774 19628
rect 4718 19574 4720 19626
rect 4720 19574 4772 19626
rect 4772 19574 4774 19626
rect 4718 19572 4774 19574
rect 4822 19626 4878 19628
rect 4822 19574 4824 19626
rect 4824 19574 4876 19626
rect 4876 19574 4878 19626
rect 4822 19572 4878 19574
rect 8016 18842 8072 18844
rect 8016 18790 8018 18842
rect 8018 18790 8070 18842
rect 8070 18790 8072 18842
rect 8016 18788 8072 18790
rect 8120 18842 8176 18844
rect 8120 18790 8122 18842
rect 8122 18790 8174 18842
rect 8174 18790 8176 18842
rect 8120 18788 8176 18790
rect 8224 18842 8280 18844
rect 8224 18790 8226 18842
rect 8226 18790 8278 18842
rect 8278 18790 8280 18842
rect 8224 18788 8280 18790
rect 2268 17666 2324 17668
rect 2268 17614 2270 17666
rect 2270 17614 2322 17666
rect 2322 17614 2324 17666
rect 2268 17612 2324 17614
rect 1708 16828 1764 16884
rect 2492 16828 2548 16884
rect 5292 18284 5348 18340
rect 4614 18058 4670 18060
rect 4614 18006 4616 18058
rect 4616 18006 4668 18058
rect 4668 18006 4670 18058
rect 4614 18004 4670 18006
rect 4718 18058 4774 18060
rect 4718 18006 4720 18058
rect 4720 18006 4772 18058
rect 4772 18006 4774 18058
rect 4718 18004 4774 18006
rect 4822 18058 4878 18060
rect 4822 18006 4824 18058
rect 4824 18006 4876 18058
rect 4876 18006 4878 18058
rect 4822 18004 4878 18006
rect 4620 16882 4676 16884
rect 4620 16830 4622 16882
rect 4622 16830 4674 16882
rect 4674 16830 4676 16882
rect 4620 16828 4676 16830
rect 5516 16716 5572 16772
rect 4614 16490 4670 16492
rect 4614 16438 4616 16490
rect 4616 16438 4668 16490
rect 4668 16438 4670 16490
rect 4614 16436 4670 16438
rect 4718 16490 4774 16492
rect 4718 16438 4720 16490
rect 4720 16438 4772 16490
rect 4772 16438 4774 16490
rect 4718 16436 4774 16438
rect 4822 16490 4878 16492
rect 4822 16438 4824 16490
rect 4824 16438 4876 16490
rect 4876 16438 4878 16490
rect 4822 16436 4878 16438
rect 8316 18620 8372 18676
rect 5964 18562 6020 18564
rect 5964 18510 5966 18562
rect 5966 18510 6018 18562
rect 6018 18510 6020 18562
rect 5964 18508 6020 18510
rect 7196 18338 7252 18340
rect 7196 18286 7198 18338
rect 7198 18286 7250 18338
rect 7250 18286 7252 18338
rect 7196 18284 7252 18286
rect 7308 17724 7364 17780
rect 5516 16044 5572 16100
rect 2828 15932 2884 15988
rect 4732 15986 4788 15988
rect 4732 15934 4734 15986
rect 4734 15934 4786 15986
rect 4786 15934 4788 15986
rect 4732 15932 4788 15934
rect 4172 15372 4228 15428
rect 4060 15260 4116 15316
rect 3052 14252 3108 14308
rect 5068 15314 5124 15316
rect 5068 15262 5070 15314
rect 5070 15262 5122 15314
rect 5122 15262 5124 15314
rect 5068 15260 5124 15262
rect 6636 16098 6692 16100
rect 6636 16046 6638 16098
rect 6638 16046 6690 16098
rect 6690 16046 6692 16098
rect 6636 16044 6692 16046
rect 7420 16828 7476 16884
rect 8428 18562 8484 18564
rect 8428 18510 8430 18562
rect 8430 18510 8482 18562
rect 8482 18510 8484 18562
rect 8428 18508 8484 18510
rect 8652 17948 8708 18004
rect 10668 19906 10724 19908
rect 10668 19854 10670 19906
rect 10670 19854 10722 19906
rect 10722 19854 10724 19906
rect 10668 19852 10724 19854
rect 11418 19626 11474 19628
rect 11418 19574 11420 19626
rect 11420 19574 11472 19626
rect 11472 19574 11474 19626
rect 11418 19572 11474 19574
rect 11522 19626 11578 19628
rect 11522 19574 11524 19626
rect 11524 19574 11576 19626
rect 11576 19574 11578 19626
rect 11522 19572 11578 19574
rect 11626 19626 11682 19628
rect 11626 19574 11628 19626
rect 11628 19574 11680 19626
rect 11680 19574 11682 19626
rect 11626 19572 11682 19574
rect 9660 18620 9716 18676
rect 10332 18172 10388 18228
rect 8016 17274 8072 17276
rect 8016 17222 8018 17274
rect 8018 17222 8070 17274
rect 8070 17222 8072 17274
rect 8016 17220 8072 17222
rect 8120 17274 8176 17276
rect 8120 17222 8122 17274
rect 8122 17222 8174 17274
rect 8174 17222 8176 17274
rect 8120 17220 8176 17222
rect 8224 17274 8280 17276
rect 8224 17222 8226 17274
rect 8226 17222 8278 17274
rect 8278 17222 8280 17274
rect 8224 17220 8280 17222
rect 7756 16044 7812 16100
rect 5292 15036 5348 15092
rect 6748 15426 6804 15428
rect 6748 15374 6750 15426
rect 6750 15374 6802 15426
rect 6802 15374 6804 15426
rect 6748 15372 6804 15374
rect 8988 16828 9044 16884
rect 8016 15706 8072 15708
rect 8016 15654 8018 15706
rect 8018 15654 8070 15706
rect 8070 15654 8072 15706
rect 8016 15652 8072 15654
rect 8120 15706 8176 15708
rect 8120 15654 8122 15706
rect 8122 15654 8174 15706
rect 8174 15654 8176 15706
rect 8120 15652 8176 15654
rect 8224 15706 8280 15708
rect 8224 15654 8226 15706
rect 8226 15654 8278 15706
rect 8278 15654 8280 15706
rect 8224 15652 8280 15654
rect 7868 15372 7924 15428
rect 6188 15036 6244 15092
rect 4614 14922 4670 14924
rect 4614 14870 4616 14922
rect 4616 14870 4668 14922
rect 4668 14870 4670 14922
rect 4614 14868 4670 14870
rect 4718 14922 4774 14924
rect 4718 14870 4720 14922
rect 4720 14870 4772 14922
rect 4772 14870 4774 14922
rect 4718 14868 4774 14870
rect 4822 14922 4878 14924
rect 4822 14870 4824 14922
rect 4824 14870 4876 14922
rect 4876 14870 4878 14922
rect 4822 14868 4878 14870
rect 4956 14364 5012 14420
rect 6076 14418 6132 14420
rect 6076 14366 6078 14418
rect 6078 14366 6130 14418
rect 6130 14366 6132 14418
rect 6076 14364 6132 14366
rect 6636 14306 6692 14308
rect 6636 14254 6638 14306
rect 6638 14254 6690 14306
rect 6690 14254 6692 14306
rect 6636 14252 6692 14254
rect 7420 14306 7476 14308
rect 7420 14254 7422 14306
rect 7422 14254 7474 14306
rect 7474 14254 7476 14306
rect 7420 14252 7476 14254
rect 6412 13580 6468 13636
rect 4614 13354 4670 13356
rect 4614 13302 4616 13354
rect 4616 13302 4668 13354
rect 4668 13302 4670 13354
rect 4614 13300 4670 13302
rect 4718 13354 4774 13356
rect 4718 13302 4720 13354
rect 4720 13302 4772 13354
rect 4772 13302 4774 13354
rect 4718 13300 4774 13302
rect 4822 13354 4878 13356
rect 4822 13302 4824 13354
rect 4824 13302 4876 13354
rect 4876 13302 4878 13354
rect 4822 13300 4878 13302
rect 7980 14812 8036 14868
rect 9772 16882 9828 16884
rect 9772 16830 9774 16882
rect 9774 16830 9826 16882
rect 9826 16830 9828 16882
rect 9772 16828 9828 16830
rect 14140 20076 14196 20132
rect 11676 18172 11732 18228
rect 11418 18058 11474 18060
rect 11418 18006 11420 18058
rect 11420 18006 11472 18058
rect 11472 18006 11474 18058
rect 11418 18004 11474 18006
rect 11522 18058 11578 18060
rect 11522 18006 11524 18058
rect 11524 18006 11576 18058
rect 11576 18006 11578 18058
rect 11522 18004 11578 18006
rect 11626 18058 11682 18060
rect 11626 18006 11628 18058
rect 11628 18006 11680 18058
rect 11680 18006 11682 18058
rect 11626 18004 11682 18006
rect 11228 17500 11284 17556
rect 12012 17554 12068 17556
rect 12012 17502 12014 17554
rect 12014 17502 12066 17554
rect 12066 17502 12068 17554
rect 12012 17500 12068 17502
rect 10668 16716 10724 16772
rect 8988 14364 9044 14420
rect 8652 14252 8708 14308
rect 8016 14138 8072 14140
rect 8016 14086 8018 14138
rect 8018 14086 8070 14138
rect 8070 14086 8072 14138
rect 8016 14084 8072 14086
rect 8120 14138 8176 14140
rect 8120 14086 8122 14138
rect 8122 14086 8174 14138
rect 8174 14086 8176 14138
rect 8120 14084 8176 14086
rect 8224 14138 8280 14140
rect 8224 14086 8226 14138
rect 8226 14086 8278 14138
rect 8278 14086 8280 14138
rect 8224 14084 8280 14086
rect 8652 13580 8708 13636
rect 4060 12908 4116 12964
rect 1820 12178 1876 12180
rect 1820 12126 1822 12178
rect 1822 12126 1874 12178
rect 1874 12126 1876 12178
rect 1820 12124 1876 12126
rect 3724 12684 3780 12740
rect 6076 12850 6132 12852
rect 6076 12798 6078 12850
rect 6078 12798 6130 12850
rect 6130 12798 6132 12850
rect 6076 12796 6132 12798
rect 7084 12796 7140 12852
rect 5852 12684 5908 12740
rect 6524 12738 6580 12740
rect 6524 12686 6526 12738
rect 6526 12686 6578 12738
rect 6578 12686 6580 12738
rect 6524 12684 6580 12686
rect 3052 11900 3108 11956
rect 4614 11786 4670 11788
rect 4614 11734 4616 11786
rect 4616 11734 4668 11786
rect 4668 11734 4670 11786
rect 4614 11732 4670 11734
rect 4718 11786 4774 11788
rect 4718 11734 4720 11786
rect 4720 11734 4772 11786
rect 4772 11734 4774 11786
rect 4718 11732 4774 11734
rect 4822 11786 4878 11788
rect 4822 11734 4824 11786
rect 4824 11734 4876 11786
rect 4876 11734 4878 11786
rect 4822 11732 4878 11734
rect 4396 11564 4452 11620
rect 5628 11340 5684 11396
rect 1820 10332 1876 10388
rect 2492 10332 2548 10388
rect 2380 9660 2436 9716
rect 1596 8092 1652 8148
rect 5628 10332 5684 10388
rect 4614 10218 4670 10220
rect 4614 10166 4616 10218
rect 4616 10166 4668 10218
rect 4668 10166 4670 10218
rect 4614 10164 4670 10166
rect 4718 10218 4774 10220
rect 4718 10166 4720 10218
rect 4720 10166 4772 10218
rect 4772 10166 4774 10218
rect 4718 10164 4774 10166
rect 4822 10218 4878 10220
rect 4822 10166 4824 10218
rect 4824 10166 4876 10218
rect 4876 10166 4878 10218
rect 4822 10164 4878 10166
rect 4284 9714 4340 9716
rect 4284 9662 4286 9714
rect 4286 9662 4338 9714
rect 4338 9662 4340 9714
rect 4284 9660 4340 9662
rect 4614 8650 4670 8652
rect 4614 8598 4616 8650
rect 4616 8598 4668 8650
rect 4668 8598 4670 8650
rect 4614 8596 4670 8598
rect 4718 8650 4774 8652
rect 4718 8598 4720 8650
rect 4720 8598 4772 8650
rect 4772 8598 4774 8650
rect 4718 8596 4774 8598
rect 4822 8650 4878 8652
rect 4822 8598 4824 8650
rect 4824 8598 4876 8650
rect 4876 8598 4878 8650
rect 4822 8596 4878 8598
rect 5068 8428 5124 8484
rect 2828 8316 2884 8372
rect 3612 8370 3668 8372
rect 3612 8318 3614 8370
rect 3614 8318 3666 8370
rect 3666 8318 3668 8370
rect 3612 8316 3668 8318
rect 4732 8316 4788 8372
rect 2492 8146 2548 8148
rect 2492 8094 2494 8146
rect 2494 8094 2546 8146
rect 2546 8094 2548 8146
rect 2492 8092 2548 8094
rect 6076 8876 6132 8932
rect 6076 8428 6132 8484
rect 5964 7532 6020 7588
rect 8016 12570 8072 12572
rect 8016 12518 8018 12570
rect 8018 12518 8070 12570
rect 8070 12518 8072 12570
rect 8016 12516 8072 12518
rect 8120 12570 8176 12572
rect 8120 12518 8122 12570
rect 8122 12518 8174 12570
rect 8174 12518 8176 12570
rect 8120 12516 8176 12518
rect 8224 12570 8280 12572
rect 8224 12518 8226 12570
rect 8226 12518 8278 12570
rect 8278 12518 8280 12570
rect 8224 12516 8280 12518
rect 8988 13580 9044 13636
rect 9324 15372 9380 15428
rect 8764 13468 8820 13524
rect 11116 16604 11172 16660
rect 11418 16490 11474 16492
rect 11418 16438 11420 16490
rect 11420 16438 11472 16490
rect 11472 16438 11474 16490
rect 11418 16436 11474 16438
rect 11522 16490 11578 16492
rect 11522 16438 11524 16490
rect 11524 16438 11576 16490
rect 11576 16438 11578 16490
rect 11522 16436 11578 16438
rect 11626 16490 11682 16492
rect 11626 16438 11628 16490
rect 11628 16438 11680 16490
rect 11680 16438 11682 16490
rect 11626 16436 11682 16438
rect 12572 15986 12628 15988
rect 12572 15934 12574 15986
rect 12574 15934 12626 15986
rect 12626 15934 12628 15986
rect 12572 15932 12628 15934
rect 10444 15372 10500 15428
rect 9660 14812 9716 14868
rect 11418 14922 11474 14924
rect 11418 14870 11420 14922
rect 11420 14870 11472 14922
rect 11472 14870 11474 14922
rect 11418 14868 11474 14870
rect 11522 14922 11578 14924
rect 11522 14870 11524 14922
rect 11524 14870 11576 14922
rect 11576 14870 11578 14922
rect 11522 14868 11578 14870
rect 11626 14922 11682 14924
rect 11626 14870 11628 14922
rect 11628 14870 11680 14922
rect 11680 14870 11682 14922
rect 11626 14868 11682 14870
rect 14028 19852 14084 19908
rect 16268 20130 16324 20132
rect 16268 20078 16270 20130
rect 16270 20078 16322 20130
rect 16322 20078 16324 20130
rect 16268 20076 16324 20078
rect 15260 19906 15316 19908
rect 15260 19854 15262 19906
rect 15262 19854 15314 19906
rect 15314 19854 15316 19906
rect 15260 19852 15316 19854
rect 21624 20410 21680 20412
rect 21624 20358 21626 20410
rect 21626 20358 21678 20410
rect 21678 20358 21680 20410
rect 21624 20356 21680 20358
rect 21728 20410 21784 20412
rect 21728 20358 21730 20410
rect 21730 20358 21782 20410
rect 21782 20358 21784 20410
rect 21728 20356 21784 20358
rect 21832 20410 21888 20412
rect 21832 20358 21834 20410
rect 21834 20358 21886 20410
rect 21886 20358 21888 20410
rect 21832 20356 21888 20358
rect 14476 18284 14532 18340
rect 14588 19404 14644 19460
rect 14364 17612 14420 17668
rect 14140 16994 14196 16996
rect 14140 16942 14142 16994
rect 14142 16942 14194 16994
rect 14194 16942 14196 16994
rect 14140 16940 14196 16942
rect 13468 16716 13524 16772
rect 12796 15426 12852 15428
rect 12796 15374 12798 15426
rect 12798 15374 12850 15426
rect 12850 15374 12852 15426
rect 12796 15372 12852 15374
rect 14028 16716 14084 16772
rect 13468 15372 13524 15428
rect 14364 15372 14420 15428
rect 11900 14418 11956 14420
rect 11900 14366 11902 14418
rect 11902 14366 11954 14418
rect 11954 14366 11956 14418
rect 11900 14364 11956 14366
rect 12796 14364 12852 14420
rect 13916 14418 13972 14420
rect 13916 14366 13918 14418
rect 13918 14366 13970 14418
rect 13970 14366 13972 14418
rect 13916 14364 13972 14366
rect 11116 13522 11172 13524
rect 11116 13470 11118 13522
rect 11118 13470 11170 13522
rect 11170 13470 11172 13522
rect 11116 13468 11172 13470
rect 11418 13354 11474 13356
rect 11418 13302 11420 13354
rect 11420 13302 11472 13354
rect 11472 13302 11474 13354
rect 11418 13300 11474 13302
rect 11522 13354 11578 13356
rect 11522 13302 11524 13354
rect 11524 13302 11576 13354
rect 11576 13302 11578 13354
rect 11522 13300 11578 13302
rect 11626 13354 11682 13356
rect 11626 13302 11628 13354
rect 11628 13302 11680 13354
rect 11680 13302 11682 13354
rect 11626 13300 11682 13302
rect 9660 12962 9716 12964
rect 9660 12910 9662 12962
rect 9662 12910 9714 12962
rect 9714 12910 9716 12962
rect 9660 12908 9716 12910
rect 14252 13580 14308 13636
rect 12796 13186 12852 13188
rect 12796 13134 12798 13186
rect 12798 13134 12850 13186
rect 12850 13134 12852 13186
rect 12796 13132 12852 13134
rect 15484 19292 15540 19348
rect 14820 18842 14876 18844
rect 14820 18790 14822 18842
rect 14822 18790 14874 18842
rect 14874 18790 14876 18842
rect 14820 18788 14876 18790
rect 14924 18842 14980 18844
rect 14924 18790 14926 18842
rect 14926 18790 14978 18842
rect 14978 18790 14980 18842
rect 14924 18788 14980 18790
rect 15028 18842 15084 18844
rect 15028 18790 15030 18842
rect 15030 18790 15082 18842
rect 15082 18790 15084 18842
rect 15028 18788 15084 18790
rect 15036 18396 15092 18452
rect 15372 18338 15428 18340
rect 15372 18286 15374 18338
rect 15374 18286 15426 18338
rect 15426 18286 15428 18338
rect 15372 18284 15428 18286
rect 17052 19122 17108 19124
rect 17052 19070 17054 19122
rect 17054 19070 17106 19122
rect 17106 19070 17108 19122
rect 17052 19068 17108 19070
rect 17500 18450 17556 18452
rect 17500 18398 17502 18450
rect 17502 18398 17554 18450
rect 17554 18398 17556 18450
rect 17500 18396 17556 18398
rect 16044 18284 16100 18340
rect 16716 18338 16772 18340
rect 16716 18286 16718 18338
rect 16718 18286 16770 18338
rect 16770 18286 16772 18338
rect 16716 18284 16772 18286
rect 16716 17612 16772 17668
rect 17612 17612 17668 17668
rect 18222 19626 18278 19628
rect 18222 19574 18224 19626
rect 18224 19574 18276 19626
rect 18276 19574 18278 19626
rect 18222 19572 18278 19574
rect 18326 19626 18382 19628
rect 18326 19574 18328 19626
rect 18328 19574 18380 19626
rect 18380 19574 18382 19626
rect 18326 19572 18382 19574
rect 18430 19626 18486 19628
rect 18430 19574 18432 19626
rect 18432 19574 18484 19626
rect 18484 19574 18486 19626
rect 18430 19572 18486 19574
rect 18284 19346 18340 19348
rect 18284 19294 18286 19346
rect 18286 19294 18338 19346
rect 18338 19294 18340 19346
rect 18284 19292 18340 19294
rect 18956 19180 19012 19236
rect 18620 18620 18676 18676
rect 17836 18284 17892 18340
rect 17948 18396 18004 18452
rect 14820 17274 14876 17276
rect 14820 17222 14822 17274
rect 14822 17222 14874 17274
rect 14874 17222 14876 17274
rect 14820 17220 14876 17222
rect 14924 17274 14980 17276
rect 14924 17222 14926 17274
rect 14926 17222 14978 17274
rect 14978 17222 14980 17274
rect 14924 17220 14980 17222
rect 15028 17274 15084 17276
rect 15028 17222 15030 17274
rect 15030 17222 15082 17274
rect 15082 17222 15084 17274
rect 15028 17220 15084 17222
rect 18222 18058 18278 18060
rect 18222 18006 18224 18058
rect 18224 18006 18276 18058
rect 18276 18006 18278 18058
rect 18222 18004 18278 18006
rect 18326 18058 18382 18060
rect 18326 18006 18328 18058
rect 18328 18006 18380 18058
rect 18380 18006 18382 18058
rect 18326 18004 18382 18006
rect 18430 18058 18486 18060
rect 18430 18006 18432 18058
rect 18432 18006 18484 18058
rect 18484 18006 18486 18058
rect 18430 18004 18486 18006
rect 19292 19122 19348 19124
rect 19292 19070 19294 19122
rect 19294 19070 19346 19122
rect 19346 19070 19348 19122
rect 19292 19068 19348 19070
rect 18956 18508 19012 18564
rect 19404 17724 19460 17780
rect 22428 20130 22484 20132
rect 22428 20078 22430 20130
rect 22430 20078 22482 20130
rect 22482 20078 22484 20130
rect 22428 20076 22484 20078
rect 21868 19852 21924 19908
rect 21420 19234 21476 19236
rect 21420 19182 21422 19234
rect 21422 19182 21474 19234
rect 21474 19182 21476 19234
rect 21420 19180 21476 19182
rect 27244 21698 27300 21700
rect 27244 21646 27246 21698
rect 27246 21646 27298 21698
rect 27298 21646 27300 21698
rect 27244 21644 27300 21646
rect 28428 23546 28484 23548
rect 28428 23494 28430 23546
rect 28430 23494 28482 23546
rect 28482 23494 28484 23546
rect 28428 23492 28484 23494
rect 28532 23546 28588 23548
rect 28532 23494 28534 23546
rect 28534 23494 28586 23546
rect 28586 23494 28588 23546
rect 28532 23492 28588 23494
rect 28636 23546 28692 23548
rect 28636 23494 28638 23546
rect 28638 23494 28690 23546
rect 28690 23494 28692 23546
rect 28636 23492 28692 23494
rect 28252 22876 28308 22932
rect 28428 21978 28484 21980
rect 28428 21926 28430 21978
rect 28430 21926 28482 21978
rect 28482 21926 28484 21978
rect 28428 21924 28484 21926
rect 28532 21978 28588 21980
rect 28532 21926 28534 21978
rect 28534 21926 28586 21978
rect 28586 21926 28588 21978
rect 28532 21924 28588 21926
rect 28636 21978 28692 21980
rect 28636 21926 28638 21978
rect 28638 21926 28690 21978
rect 28690 21926 28692 21978
rect 28636 21924 28692 21926
rect 28140 21532 28196 21588
rect 25026 21194 25082 21196
rect 25026 21142 25028 21194
rect 25028 21142 25080 21194
rect 25080 21142 25082 21194
rect 25026 21140 25082 21142
rect 25130 21194 25186 21196
rect 25130 21142 25132 21194
rect 25132 21142 25184 21194
rect 25184 21142 25186 21194
rect 25130 21140 25186 21142
rect 25234 21194 25290 21196
rect 25234 21142 25236 21194
rect 25236 21142 25288 21194
rect 25288 21142 25290 21194
rect 25234 21140 25290 21142
rect 26236 21474 26292 21476
rect 26236 21422 26238 21474
rect 26238 21422 26290 21474
rect 26290 21422 26292 21474
rect 26236 21420 26292 21422
rect 26124 20636 26180 20692
rect 26908 20690 26964 20692
rect 26908 20638 26910 20690
rect 26910 20638 26962 20690
rect 26962 20638 26964 20690
rect 26908 20636 26964 20638
rect 25026 19626 25082 19628
rect 25026 19574 25028 19626
rect 25028 19574 25080 19626
rect 25080 19574 25082 19626
rect 25026 19572 25082 19574
rect 25130 19626 25186 19628
rect 25130 19574 25132 19626
rect 25132 19574 25184 19626
rect 25184 19574 25186 19626
rect 25130 19572 25186 19574
rect 25234 19626 25290 19628
rect 25234 19574 25236 19626
rect 25236 19574 25288 19626
rect 25288 19574 25290 19626
rect 25234 19572 25290 19574
rect 22764 19180 22820 19236
rect 21624 18842 21680 18844
rect 21624 18790 21626 18842
rect 21626 18790 21678 18842
rect 21678 18790 21680 18842
rect 21624 18788 21680 18790
rect 21728 18842 21784 18844
rect 21728 18790 21730 18842
rect 21730 18790 21782 18842
rect 21782 18790 21784 18842
rect 21728 18788 21784 18790
rect 21832 18842 21888 18844
rect 21832 18790 21834 18842
rect 21834 18790 21886 18842
rect 21886 18790 21888 18842
rect 21832 18788 21888 18790
rect 22764 18508 22820 18564
rect 23212 18620 23268 18676
rect 25900 20018 25956 20020
rect 25900 19966 25902 20018
rect 25902 19966 25954 20018
rect 25954 19966 25956 20018
rect 25900 19964 25956 19966
rect 22204 18338 22260 18340
rect 22204 18286 22206 18338
rect 22206 18286 22258 18338
rect 22258 18286 22260 18338
rect 22204 18284 22260 18286
rect 24892 18396 24948 18452
rect 24108 18284 24164 18340
rect 20972 18226 21028 18228
rect 20972 18174 20974 18226
rect 20974 18174 21026 18226
rect 21026 18174 21028 18226
rect 20972 18172 21028 18174
rect 23548 18172 23604 18228
rect 22316 17778 22372 17780
rect 22316 17726 22318 17778
rect 22318 17726 22370 17778
rect 22370 17726 22372 17778
rect 22316 17724 22372 17726
rect 16380 16994 16436 16996
rect 16380 16942 16382 16994
rect 16382 16942 16434 16994
rect 16434 16942 16436 16994
rect 16380 16940 16436 16942
rect 15372 16770 15428 16772
rect 15372 16718 15374 16770
rect 15374 16718 15426 16770
rect 15426 16718 15428 16770
rect 15372 16716 15428 16718
rect 15708 16716 15764 16772
rect 15708 15932 15764 15988
rect 14820 15706 14876 15708
rect 14820 15654 14822 15706
rect 14822 15654 14874 15706
rect 14874 15654 14876 15706
rect 14820 15652 14876 15654
rect 14924 15706 14980 15708
rect 14924 15654 14926 15706
rect 14926 15654 14978 15706
rect 14978 15654 14980 15706
rect 14924 15652 14980 15654
rect 15028 15706 15084 15708
rect 15028 15654 15030 15706
rect 15030 15654 15082 15706
rect 15082 15654 15084 15706
rect 15028 15652 15084 15654
rect 16268 16156 16324 16212
rect 14700 15372 14756 15428
rect 15148 15426 15204 15428
rect 15148 15374 15150 15426
rect 15150 15374 15202 15426
rect 15202 15374 15204 15426
rect 15148 15372 15204 15374
rect 15148 14476 15204 14532
rect 14820 14138 14876 14140
rect 14820 14086 14822 14138
rect 14822 14086 14874 14138
rect 14874 14086 14876 14138
rect 14820 14084 14876 14086
rect 14924 14138 14980 14140
rect 14924 14086 14926 14138
rect 14926 14086 14978 14138
rect 14978 14086 14980 14138
rect 14924 14084 14980 14086
rect 15028 14138 15084 14140
rect 15028 14086 15030 14138
rect 15030 14086 15082 14138
rect 15082 14086 15084 14138
rect 15028 14084 15084 14086
rect 15820 14530 15876 14532
rect 15820 14478 15822 14530
rect 15822 14478 15874 14530
rect 15874 14478 15876 14530
rect 15820 14476 15876 14478
rect 17052 15986 17108 15988
rect 17052 15934 17054 15986
rect 17054 15934 17106 15986
rect 17106 15934 17108 15986
rect 17052 15932 17108 15934
rect 16492 15874 16548 15876
rect 16492 15822 16494 15874
rect 16494 15822 16546 15874
rect 16546 15822 16548 15874
rect 16492 15820 16548 15822
rect 18284 16716 18340 16772
rect 18620 16604 18676 16660
rect 18222 16490 18278 16492
rect 18222 16438 18224 16490
rect 18224 16438 18276 16490
rect 18276 16438 18278 16490
rect 18222 16436 18278 16438
rect 18326 16490 18382 16492
rect 18326 16438 18328 16490
rect 18328 16438 18380 16490
rect 18380 16438 18382 16490
rect 18326 16436 18382 16438
rect 18430 16490 18486 16492
rect 18430 16438 18432 16490
rect 18432 16438 18484 16490
rect 18484 16438 18486 16490
rect 18430 16436 18486 16438
rect 18284 16210 18340 16212
rect 18284 16158 18286 16210
rect 18286 16158 18338 16210
rect 18338 16158 18340 16210
rect 18284 16156 18340 16158
rect 18396 15314 18452 15316
rect 18396 15262 18398 15314
rect 18398 15262 18450 15314
rect 18450 15262 18452 15314
rect 18396 15260 18452 15262
rect 18222 14922 18278 14924
rect 18222 14870 18224 14922
rect 18224 14870 18276 14922
rect 18276 14870 18278 14922
rect 18222 14868 18278 14870
rect 18326 14922 18382 14924
rect 18326 14870 18328 14922
rect 18328 14870 18380 14922
rect 18380 14870 18382 14922
rect 18326 14868 18382 14870
rect 18430 14922 18486 14924
rect 18430 14870 18432 14922
rect 18432 14870 18484 14922
rect 18484 14870 18486 14922
rect 18430 14868 18486 14870
rect 17836 14476 17892 14532
rect 19628 17666 19684 17668
rect 19628 17614 19630 17666
rect 19630 17614 19682 17666
rect 19682 17614 19684 17666
rect 19628 17612 19684 17614
rect 20524 17666 20580 17668
rect 20524 17614 20526 17666
rect 20526 17614 20578 17666
rect 20578 17614 20580 17666
rect 20524 17612 20580 17614
rect 21420 17666 21476 17668
rect 21420 17614 21422 17666
rect 21422 17614 21474 17666
rect 21474 17614 21476 17666
rect 21420 17612 21476 17614
rect 21868 17666 21924 17668
rect 21868 17614 21870 17666
rect 21870 17614 21922 17666
rect 21922 17614 21924 17666
rect 21868 17612 21924 17614
rect 26236 19906 26292 19908
rect 26236 19854 26238 19906
rect 26238 19854 26290 19906
rect 26290 19854 26292 19906
rect 26236 19852 26292 19854
rect 25900 18284 25956 18340
rect 24220 17612 24276 17668
rect 21624 17274 21680 17276
rect 21624 17222 21626 17274
rect 21626 17222 21678 17274
rect 21678 17222 21680 17274
rect 21624 17220 21680 17222
rect 21728 17274 21784 17276
rect 21728 17222 21730 17274
rect 21730 17222 21782 17274
rect 21782 17222 21784 17274
rect 21728 17220 21784 17222
rect 21832 17274 21888 17276
rect 21832 17222 21834 17274
rect 21834 17222 21886 17274
rect 21886 17222 21888 17274
rect 21832 17220 21888 17222
rect 18956 16828 19012 16884
rect 19740 16828 19796 16884
rect 19292 15986 19348 15988
rect 19292 15934 19294 15986
rect 19294 15934 19346 15986
rect 19346 15934 19348 15986
rect 19292 15932 19348 15934
rect 19292 15372 19348 15428
rect 24444 17052 24500 17108
rect 23436 16940 23492 16996
rect 24220 16994 24276 16996
rect 24220 16942 24222 16994
rect 24222 16942 24274 16994
rect 24274 16942 24276 16994
rect 24220 16940 24276 16942
rect 20300 16716 20356 16772
rect 19964 15932 20020 15988
rect 20300 15874 20356 15876
rect 20300 15822 20302 15874
rect 20302 15822 20354 15874
rect 20354 15822 20356 15874
rect 20300 15820 20356 15822
rect 20524 15484 20580 15540
rect 25026 18058 25082 18060
rect 25026 18006 25028 18058
rect 25028 18006 25080 18058
rect 25080 18006 25082 18058
rect 25026 18004 25082 18006
rect 25130 18058 25186 18060
rect 25130 18006 25132 18058
rect 25132 18006 25184 18058
rect 25184 18006 25186 18058
rect 25130 18004 25186 18006
rect 25234 18058 25290 18060
rect 25234 18006 25236 18058
rect 25236 18006 25288 18058
rect 25288 18006 25290 18058
rect 25234 18004 25290 18006
rect 27244 20130 27300 20132
rect 27244 20078 27246 20130
rect 27246 20078 27298 20130
rect 27298 20078 27300 20130
rect 27244 20076 27300 20078
rect 27356 19964 27412 20020
rect 26908 19068 26964 19124
rect 28428 20410 28484 20412
rect 28428 20358 28430 20410
rect 28430 20358 28482 20410
rect 28482 20358 28484 20410
rect 28428 20356 28484 20358
rect 28532 20410 28588 20412
rect 28532 20358 28534 20410
rect 28534 20358 28586 20410
rect 28586 20358 28588 20410
rect 28532 20356 28588 20358
rect 28636 20410 28692 20412
rect 28636 20358 28638 20410
rect 28638 20358 28690 20410
rect 28690 20358 28692 20410
rect 28636 20356 28692 20358
rect 27692 19122 27748 19124
rect 27692 19070 27694 19122
rect 27694 19070 27746 19122
rect 27746 19070 27748 19122
rect 27692 19068 27748 19070
rect 28428 18842 28484 18844
rect 28428 18790 28430 18842
rect 28430 18790 28482 18842
rect 28482 18790 28484 18842
rect 28428 18788 28484 18790
rect 28532 18842 28588 18844
rect 28532 18790 28534 18842
rect 28534 18790 28586 18842
rect 28586 18790 28588 18842
rect 28532 18788 28588 18790
rect 28636 18842 28692 18844
rect 28636 18790 28638 18842
rect 28638 18790 28690 18842
rect 28690 18790 28692 18842
rect 28636 18788 28692 18790
rect 28428 17274 28484 17276
rect 28428 17222 28430 17274
rect 28430 17222 28482 17274
rect 28482 17222 28484 17274
rect 28428 17220 28484 17222
rect 28532 17274 28588 17276
rect 28532 17222 28534 17274
rect 28534 17222 28586 17274
rect 28586 17222 28588 17274
rect 28532 17220 28588 17222
rect 28636 17274 28692 17276
rect 28636 17222 28638 17274
rect 28638 17222 28690 17274
rect 28690 17222 28692 17274
rect 28636 17220 28692 17222
rect 25340 17106 25396 17108
rect 25340 17054 25342 17106
rect 25342 17054 25394 17106
rect 25394 17054 25396 17106
rect 25340 17052 25396 17054
rect 27132 17052 27188 17108
rect 24892 16828 24948 16884
rect 21624 15706 21680 15708
rect 21624 15654 21626 15706
rect 21626 15654 21678 15706
rect 21678 15654 21680 15706
rect 21624 15652 21680 15654
rect 21728 15706 21784 15708
rect 21728 15654 21730 15706
rect 21730 15654 21782 15706
rect 21782 15654 21784 15706
rect 21728 15652 21784 15654
rect 21832 15706 21888 15708
rect 21832 15654 21834 15706
rect 21834 15654 21886 15706
rect 21886 15654 21888 15706
rect 21832 15652 21888 15654
rect 19740 14306 19796 14308
rect 19740 14254 19742 14306
rect 19742 14254 19794 14306
rect 19794 14254 19796 14306
rect 19740 14252 19796 14254
rect 20636 14252 20692 14308
rect 18396 13634 18452 13636
rect 18396 13582 18398 13634
rect 18398 13582 18450 13634
rect 18450 13582 18452 13634
rect 18396 13580 18452 13582
rect 14476 13020 14532 13076
rect 18222 13354 18278 13356
rect 18222 13302 18224 13354
rect 18224 13302 18276 13354
rect 18276 13302 18278 13354
rect 18222 13300 18278 13302
rect 18326 13354 18382 13356
rect 18326 13302 18328 13354
rect 18328 13302 18380 13354
rect 18380 13302 18382 13354
rect 18326 13300 18382 13302
rect 18430 13354 18486 13356
rect 18430 13302 18432 13354
rect 18432 13302 18484 13354
rect 18484 13302 18486 13354
rect 18430 13300 18486 13302
rect 19404 13132 19460 13188
rect 20076 13020 20132 13076
rect 14820 12570 14876 12572
rect 14820 12518 14822 12570
rect 14822 12518 14874 12570
rect 14874 12518 14876 12570
rect 14820 12516 14876 12518
rect 14924 12570 14980 12572
rect 14924 12518 14926 12570
rect 14926 12518 14978 12570
rect 14978 12518 14980 12570
rect 14924 12516 14980 12518
rect 15028 12570 15084 12572
rect 15028 12518 15030 12570
rect 15030 12518 15082 12570
rect 15082 12518 15084 12570
rect 15028 12516 15084 12518
rect 20076 12348 20132 12404
rect 8876 12066 8932 12068
rect 8876 12014 8878 12066
rect 8878 12014 8930 12066
rect 8930 12014 8932 12066
rect 8876 12012 8932 12014
rect 7196 11900 7252 11956
rect 7980 11676 8036 11732
rect 8016 11002 8072 11004
rect 8016 10950 8018 11002
rect 8018 10950 8070 11002
rect 8070 10950 8072 11002
rect 8016 10948 8072 10950
rect 8120 11002 8176 11004
rect 8120 10950 8122 11002
rect 8122 10950 8174 11002
rect 8174 10950 8176 11002
rect 8120 10948 8176 10950
rect 8224 11002 8280 11004
rect 8224 10950 8226 11002
rect 8226 10950 8278 11002
rect 8278 10950 8280 11002
rect 8224 10948 8280 10950
rect 8316 10834 8372 10836
rect 8316 10782 8318 10834
rect 8318 10782 8370 10834
rect 8370 10782 8372 10834
rect 8316 10780 8372 10782
rect 8016 9434 8072 9436
rect 8016 9382 8018 9434
rect 8018 9382 8070 9434
rect 8070 9382 8072 9434
rect 8016 9380 8072 9382
rect 8120 9434 8176 9436
rect 8120 9382 8122 9434
rect 8122 9382 8174 9434
rect 8174 9382 8176 9434
rect 8120 9380 8176 9382
rect 8224 9434 8280 9436
rect 8224 9382 8226 9434
rect 8226 9382 8278 9434
rect 8278 9382 8280 9434
rect 8224 9380 8280 9382
rect 7532 8930 7588 8932
rect 7532 8878 7534 8930
rect 7534 8878 7586 8930
rect 7586 8878 7588 8930
rect 7532 8876 7588 8878
rect 6524 8428 6580 8484
rect 7420 8370 7476 8372
rect 7420 8318 7422 8370
rect 7422 8318 7474 8370
rect 7474 8318 7476 8370
rect 7420 8316 7476 8318
rect 4614 7082 4670 7084
rect 4614 7030 4616 7082
rect 4616 7030 4668 7082
rect 4668 7030 4670 7082
rect 4614 7028 4670 7030
rect 4718 7082 4774 7084
rect 4718 7030 4720 7082
rect 4720 7030 4772 7082
rect 4772 7030 4774 7082
rect 4718 7028 4774 7030
rect 4822 7082 4878 7084
rect 4822 7030 4824 7082
rect 4824 7030 4876 7082
rect 4876 7030 4878 7082
rect 4822 7028 4878 7030
rect 8016 7866 8072 7868
rect 8016 7814 8018 7866
rect 8018 7814 8070 7866
rect 8070 7814 8072 7866
rect 8016 7812 8072 7814
rect 8120 7866 8176 7868
rect 8120 7814 8122 7866
rect 8122 7814 8174 7866
rect 8174 7814 8176 7866
rect 8120 7812 8176 7814
rect 8224 7866 8280 7868
rect 8224 7814 8226 7866
rect 8226 7814 8278 7866
rect 8278 7814 8280 7866
rect 8224 7812 8280 7814
rect 11418 11786 11474 11788
rect 10108 11676 10164 11732
rect 10668 11676 10724 11732
rect 11418 11734 11420 11786
rect 11420 11734 11472 11786
rect 11472 11734 11474 11786
rect 11418 11732 11474 11734
rect 11522 11786 11578 11788
rect 11522 11734 11524 11786
rect 11524 11734 11576 11786
rect 11576 11734 11578 11786
rect 11522 11732 11578 11734
rect 11626 11786 11682 11788
rect 11626 11734 11628 11786
rect 11628 11734 11680 11786
rect 11680 11734 11682 11786
rect 11626 11732 11682 11734
rect 10332 11394 10388 11396
rect 10332 11342 10334 11394
rect 10334 11342 10386 11394
rect 10386 11342 10388 11394
rect 10332 11340 10388 11342
rect 10108 11116 10164 11172
rect 9324 9100 9380 9156
rect 7196 7586 7252 7588
rect 7196 7534 7198 7586
rect 7198 7534 7250 7586
rect 7250 7534 7252 7586
rect 7196 7532 7252 7534
rect 6524 6636 6580 6692
rect 7980 6690 8036 6692
rect 7980 6638 7982 6690
rect 7982 6638 8034 6690
rect 8034 6638 8036 6690
rect 7980 6636 8036 6638
rect 14588 11340 14644 11396
rect 11900 11116 11956 11172
rect 11116 10780 11172 10836
rect 10668 10556 10724 10612
rect 12460 10610 12516 10612
rect 12460 10558 12462 10610
rect 12462 10558 12514 10610
rect 12514 10558 12516 10610
rect 12460 10556 12516 10558
rect 11228 10498 11284 10500
rect 11228 10446 11230 10498
rect 11230 10446 11282 10498
rect 11282 10446 11284 10498
rect 11228 10444 11284 10446
rect 11418 10218 11474 10220
rect 11418 10166 11420 10218
rect 11420 10166 11472 10218
rect 11472 10166 11474 10218
rect 11418 10164 11474 10166
rect 11522 10218 11578 10220
rect 11522 10166 11524 10218
rect 11524 10166 11576 10218
rect 11576 10166 11578 10218
rect 11522 10164 11578 10166
rect 11626 10218 11682 10220
rect 11626 10166 11628 10218
rect 11628 10166 11680 10218
rect 11680 10166 11682 10218
rect 11626 10164 11682 10166
rect 11116 9772 11172 9828
rect 10108 9154 10164 9156
rect 10108 9102 10110 9154
rect 10110 9102 10162 9154
rect 10162 9102 10164 9154
rect 10108 9100 10164 9102
rect 10108 8034 10164 8036
rect 10108 7982 10110 8034
rect 10110 7982 10162 8034
rect 10162 7982 10164 8034
rect 10108 7980 10164 7982
rect 12348 9826 12404 9828
rect 12348 9774 12350 9826
rect 12350 9774 12402 9826
rect 12402 9774 12404 9826
rect 12348 9772 12404 9774
rect 13020 10444 13076 10500
rect 12908 10108 12964 10164
rect 11452 8988 11508 9044
rect 11418 8650 11474 8652
rect 11418 8598 11420 8650
rect 11420 8598 11472 8650
rect 11472 8598 11474 8650
rect 11418 8596 11474 8598
rect 11522 8650 11578 8652
rect 11522 8598 11524 8650
rect 11524 8598 11576 8650
rect 11576 8598 11578 8650
rect 11522 8596 11578 8598
rect 11626 8650 11682 8652
rect 11626 8598 11628 8650
rect 11628 8598 11680 8650
rect 11680 8598 11682 8650
rect 11626 8596 11682 8598
rect 12460 8258 12516 8260
rect 12460 8206 12462 8258
rect 12462 8206 12514 8258
rect 12514 8206 12516 8258
rect 12460 8204 12516 8206
rect 13244 9042 13300 9044
rect 13244 8990 13246 9042
rect 13246 8990 13298 9042
rect 13298 8990 13300 9042
rect 13244 8988 13300 8990
rect 12460 7980 12516 8036
rect 14140 7980 14196 8036
rect 14476 8204 14532 8260
rect 13244 7362 13300 7364
rect 13244 7310 13246 7362
rect 13246 7310 13298 7362
rect 13298 7310 13300 7362
rect 13244 7308 13300 7310
rect 11418 7082 11474 7084
rect 11418 7030 11420 7082
rect 11420 7030 11472 7082
rect 11472 7030 11474 7082
rect 11418 7028 11474 7030
rect 11522 7082 11578 7084
rect 11522 7030 11524 7082
rect 11524 7030 11576 7082
rect 11576 7030 11578 7082
rect 11522 7028 11578 7030
rect 11626 7082 11682 7084
rect 11626 7030 11628 7082
rect 11628 7030 11680 7082
rect 11680 7030 11682 7082
rect 11626 7028 11682 7030
rect 12684 6748 12740 6804
rect 14820 11002 14876 11004
rect 14820 10950 14822 11002
rect 14822 10950 14874 11002
rect 14874 10950 14876 11002
rect 14820 10948 14876 10950
rect 14924 11002 14980 11004
rect 14924 10950 14926 11002
rect 14926 10950 14978 11002
rect 14978 10950 14980 11002
rect 14924 10948 14980 10950
rect 15028 11002 15084 11004
rect 15028 10950 15030 11002
rect 15030 10950 15082 11002
rect 15082 10950 15084 11002
rect 15028 10948 15084 10950
rect 15596 10834 15652 10836
rect 15596 10782 15598 10834
rect 15598 10782 15650 10834
rect 15650 10782 15652 10834
rect 15596 10780 15652 10782
rect 15148 10108 15204 10164
rect 14820 9434 14876 9436
rect 14820 9382 14822 9434
rect 14822 9382 14874 9434
rect 14874 9382 14876 9434
rect 14820 9380 14876 9382
rect 14924 9434 14980 9436
rect 14924 9382 14926 9434
rect 14926 9382 14978 9434
rect 14978 9382 14980 9434
rect 14924 9380 14980 9382
rect 15028 9434 15084 9436
rect 15028 9382 15030 9434
rect 15030 9382 15082 9434
rect 15082 9382 15084 9434
rect 15028 9380 15084 9382
rect 14820 7866 14876 7868
rect 14820 7814 14822 7866
rect 14822 7814 14874 7866
rect 14874 7814 14876 7866
rect 14820 7812 14876 7814
rect 14924 7866 14980 7868
rect 14924 7814 14926 7866
rect 14926 7814 14978 7866
rect 14978 7814 14980 7866
rect 14924 7812 14980 7814
rect 15028 7866 15084 7868
rect 15028 7814 15030 7866
rect 15030 7814 15082 7866
rect 15082 7814 15084 7866
rect 15028 7812 15084 7814
rect 15148 7308 15204 7364
rect 8652 6690 8708 6692
rect 8652 6638 8654 6690
rect 8654 6638 8706 6690
rect 8706 6638 8708 6690
rect 8652 6636 8708 6638
rect 8016 6298 8072 6300
rect 8016 6246 8018 6298
rect 8018 6246 8070 6298
rect 8070 6246 8072 6298
rect 8016 6244 8072 6246
rect 8120 6298 8176 6300
rect 8120 6246 8122 6298
rect 8122 6246 8174 6298
rect 8174 6246 8176 6298
rect 8120 6244 8176 6246
rect 8224 6298 8280 6300
rect 8224 6246 8226 6298
rect 8226 6246 8278 6298
rect 8278 6246 8280 6298
rect 8224 6244 8280 6246
rect 14820 6298 14876 6300
rect 14820 6246 14822 6298
rect 14822 6246 14874 6298
rect 14874 6246 14876 6298
rect 14820 6244 14876 6246
rect 14924 6298 14980 6300
rect 14924 6246 14926 6298
rect 14926 6246 14978 6298
rect 14978 6246 14980 6298
rect 14924 6244 14980 6246
rect 15028 6298 15084 6300
rect 15028 6246 15030 6298
rect 15030 6246 15082 6298
rect 15082 6246 15084 6298
rect 15028 6244 15084 6246
rect 12572 5852 12628 5908
rect 4614 5514 4670 5516
rect 4614 5462 4616 5514
rect 4616 5462 4668 5514
rect 4668 5462 4670 5514
rect 4614 5460 4670 5462
rect 4718 5514 4774 5516
rect 4718 5462 4720 5514
rect 4720 5462 4772 5514
rect 4772 5462 4774 5514
rect 4718 5460 4774 5462
rect 4822 5514 4878 5516
rect 4822 5462 4824 5514
rect 4824 5462 4876 5514
rect 4876 5462 4878 5514
rect 4822 5460 4878 5462
rect 11418 5514 11474 5516
rect 11418 5462 11420 5514
rect 11420 5462 11472 5514
rect 11472 5462 11474 5514
rect 11418 5460 11474 5462
rect 11522 5514 11578 5516
rect 11522 5462 11524 5514
rect 11524 5462 11576 5514
rect 11576 5462 11578 5514
rect 11522 5460 11578 5462
rect 11626 5514 11682 5516
rect 11626 5462 11628 5514
rect 11628 5462 11680 5514
rect 11680 5462 11682 5514
rect 11626 5460 11682 5462
rect 8016 4730 8072 4732
rect 8016 4678 8018 4730
rect 8018 4678 8070 4730
rect 8070 4678 8072 4730
rect 8016 4676 8072 4678
rect 8120 4730 8176 4732
rect 8120 4678 8122 4730
rect 8122 4678 8174 4730
rect 8174 4678 8176 4730
rect 8120 4676 8176 4678
rect 8224 4730 8280 4732
rect 8224 4678 8226 4730
rect 8226 4678 8278 4730
rect 8278 4678 8280 4730
rect 8224 4676 8280 4678
rect 4614 3946 4670 3948
rect 4614 3894 4616 3946
rect 4616 3894 4668 3946
rect 4668 3894 4670 3946
rect 4614 3892 4670 3894
rect 4718 3946 4774 3948
rect 4718 3894 4720 3946
rect 4720 3894 4772 3946
rect 4772 3894 4774 3946
rect 4718 3892 4774 3894
rect 4822 3946 4878 3948
rect 4822 3894 4824 3946
rect 4824 3894 4876 3946
rect 4876 3894 4878 3946
rect 4822 3892 4878 3894
rect 11418 3946 11474 3948
rect 11418 3894 11420 3946
rect 11420 3894 11472 3946
rect 11472 3894 11474 3946
rect 11418 3892 11474 3894
rect 11522 3946 11578 3948
rect 11522 3894 11524 3946
rect 11524 3894 11576 3946
rect 11576 3894 11578 3946
rect 11522 3892 11578 3894
rect 11626 3946 11682 3948
rect 11626 3894 11628 3946
rect 11628 3894 11680 3946
rect 11680 3894 11682 3946
rect 11626 3892 11682 3894
rect 8016 3162 8072 3164
rect 8016 3110 8018 3162
rect 8018 3110 8070 3162
rect 8070 3110 8072 3162
rect 8016 3108 8072 3110
rect 8120 3162 8176 3164
rect 8120 3110 8122 3162
rect 8122 3110 8174 3162
rect 8174 3110 8176 3162
rect 8120 3108 8176 3110
rect 8224 3162 8280 3164
rect 8224 3110 8226 3162
rect 8226 3110 8278 3162
rect 8278 3110 8280 3162
rect 8224 3108 8280 3110
rect 13468 5906 13524 5908
rect 13468 5854 13470 5906
rect 13470 5854 13522 5906
rect 13522 5854 13524 5906
rect 13468 5852 13524 5854
rect 15708 8988 15764 9044
rect 16380 10780 16436 10836
rect 16716 10498 16772 10500
rect 16716 10446 16718 10498
rect 16718 10446 16770 10498
rect 16770 10446 16772 10498
rect 16716 10444 16772 10446
rect 16268 9996 16324 10052
rect 16156 8316 16212 8372
rect 16380 8092 16436 8148
rect 16828 8034 16884 8036
rect 16828 7982 16830 8034
rect 16830 7982 16882 8034
rect 16882 7982 16884 8034
rect 16828 7980 16884 7982
rect 16268 7586 16324 7588
rect 16268 7534 16270 7586
rect 16270 7534 16322 7586
rect 16322 7534 16324 7586
rect 16268 7532 16324 7534
rect 19628 12124 19684 12180
rect 18222 11786 18278 11788
rect 18222 11734 18224 11786
rect 18224 11734 18276 11786
rect 18276 11734 18278 11786
rect 18222 11732 18278 11734
rect 18326 11786 18382 11788
rect 18326 11734 18328 11786
rect 18328 11734 18380 11786
rect 18380 11734 18382 11786
rect 18326 11732 18382 11734
rect 18430 11786 18486 11788
rect 18430 11734 18432 11786
rect 18432 11734 18484 11786
rect 18484 11734 18486 11786
rect 18430 11732 18486 11734
rect 18060 11452 18116 11508
rect 19180 11394 19236 11396
rect 19180 11342 19182 11394
rect 19182 11342 19234 11394
rect 19234 11342 19236 11394
rect 19180 11340 19236 11342
rect 18620 11228 18676 11284
rect 19404 11282 19460 11284
rect 19404 11230 19406 11282
rect 19406 11230 19458 11282
rect 19458 11230 19460 11282
rect 19404 11228 19460 11230
rect 17500 10498 17556 10500
rect 17500 10446 17502 10498
rect 17502 10446 17554 10498
rect 17554 10446 17556 10498
rect 17500 10444 17556 10446
rect 20300 12124 20356 12180
rect 20412 12236 20468 12292
rect 20748 13580 20804 13636
rect 20188 11452 20244 11508
rect 18222 10218 18278 10220
rect 18222 10166 18224 10218
rect 18224 10166 18276 10218
rect 18276 10166 18278 10218
rect 18222 10164 18278 10166
rect 18326 10218 18382 10220
rect 18326 10166 18328 10218
rect 18328 10166 18380 10218
rect 18380 10166 18382 10218
rect 18326 10164 18382 10166
rect 18430 10218 18486 10220
rect 18430 10166 18432 10218
rect 18432 10166 18484 10218
rect 18484 10166 18486 10218
rect 18430 10164 18486 10166
rect 18620 9660 18676 9716
rect 19180 9602 19236 9604
rect 19180 9550 19182 9602
rect 19182 9550 19234 9602
rect 19234 9550 19236 9602
rect 19180 9548 19236 9550
rect 17500 9042 17556 9044
rect 17500 8990 17502 9042
rect 17502 8990 17554 9042
rect 17554 8990 17556 9042
rect 17500 8988 17556 8990
rect 19740 9938 19796 9940
rect 19740 9886 19742 9938
rect 19742 9886 19794 9938
rect 19794 9886 19796 9938
rect 19740 9884 19796 9886
rect 20300 9884 20356 9940
rect 19404 9714 19460 9716
rect 19404 9662 19406 9714
rect 19406 9662 19458 9714
rect 19458 9662 19460 9714
rect 19404 9660 19460 9662
rect 19292 8988 19348 9044
rect 18172 8876 18228 8932
rect 18222 8650 18278 8652
rect 18222 8598 18224 8650
rect 18224 8598 18276 8650
rect 18276 8598 18278 8650
rect 18222 8596 18278 8598
rect 18326 8650 18382 8652
rect 18326 8598 18328 8650
rect 18328 8598 18380 8650
rect 18380 8598 18382 8650
rect 18326 8596 18382 8598
rect 18430 8650 18486 8652
rect 18430 8598 18432 8650
rect 18432 8598 18484 8650
rect 18484 8598 18486 8650
rect 18430 8596 18486 8598
rect 17612 8370 17668 8372
rect 17612 8318 17614 8370
rect 17614 8318 17666 8370
rect 17666 8318 17668 8370
rect 17612 8316 17668 8318
rect 18620 8146 18676 8148
rect 18620 8094 18622 8146
rect 18622 8094 18674 8146
rect 18674 8094 18676 8146
rect 18620 8092 18676 8094
rect 21420 15314 21476 15316
rect 21420 15262 21422 15314
rect 21422 15262 21474 15314
rect 21474 15262 21476 15314
rect 21420 15260 21476 15262
rect 21756 15538 21812 15540
rect 21756 15486 21758 15538
rect 21758 15486 21810 15538
rect 21810 15486 21812 15538
rect 21756 15484 21812 15486
rect 21868 14252 21924 14308
rect 21624 14138 21680 14140
rect 21624 14086 21626 14138
rect 21626 14086 21678 14138
rect 21678 14086 21680 14138
rect 21624 14084 21680 14086
rect 21728 14138 21784 14140
rect 21728 14086 21730 14138
rect 21730 14086 21782 14138
rect 21782 14086 21784 14138
rect 21728 14084 21784 14086
rect 21832 14138 21888 14140
rect 21832 14086 21834 14138
rect 21834 14086 21886 14138
rect 21886 14086 21888 14138
rect 21832 14084 21888 14086
rect 21624 12570 21680 12572
rect 21624 12518 21626 12570
rect 21626 12518 21678 12570
rect 21678 12518 21680 12570
rect 21624 12516 21680 12518
rect 21728 12570 21784 12572
rect 21728 12518 21730 12570
rect 21730 12518 21782 12570
rect 21782 12518 21784 12570
rect 21728 12516 21784 12518
rect 21832 12570 21888 12572
rect 21832 12518 21834 12570
rect 21834 12518 21886 12570
rect 21886 12518 21888 12570
rect 21832 12516 21888 12518
rect 23212 15932 23268 15988
rect 22652 15202 22708 15204
rect 22652 15150 22654 15202
rect 22654 15150 22706 15202
rect 22706 15150 22708 15202
rect 22652 15148 22708 15150
rect 23660 15426 23716 15428
rect 23660 15374 23662 15426
rect 23662 15374 23714 15426
rect 23714 15374 23716 15426
rect 23660 15372 23716 15374
rect 23996 15372 24052 15428
rect 25026 16490 25082 16492
rect 25026 16438 25028 16490
rect 25028 16438 25080 16490
rect 25080 16438 25082 16490
rect 25026 16436 25082 16438
rect 25130 16490 25186 16492
rect 25130 16438 25132 16490
rect 25132 16438 25184 16490
rect 25184 16438 25186 16490
rect 25130 16436 25186 16438
rect 25234 16490 25290 16492
rect 25234 16438 25236 16490
rect 25236 16438 25288 16490
rect 25288 16438 25290 16490
rect 25234 16436 25290 16438
rect 24892 15484 24948 15540
rect 23772 14700 23828 14756
rect 22316 14252 22372 14308
rect 22652 13916 22708 13972
rect 25340 15426 25396 15428
rect 25340 15374 25342 15426
rect 25342 15374 25394 15426
rect 25394 15374 25396 15426
rect 25340 15372 25396 15374
rect 25026 14922 25082 14924
rect 25026 14870 25028 14922
rect 25028 14870 25080 14922
rect 25080 14870 25082 14922
rect 25026 14868 25082 14870
rect 25130 14922 25186 14924
rect 25130 14870 25132 14922
rect 25132 14870 25184 14922
rect 25184 14870 25186 14922
rect 25130 14868 25186 14870
rect 25234 14922 25290 14924
rect 25234 14870 25236 14922
rect 25236 14870 25288 14922
rect 25288 14870 25290 14922
rect 25234 14868 25290 14870
rect 24892 14476 24948 14532
rect 23996 14306 24052 14308
rect 23996 14254 23998 14306
rect 23998 14254 24050 14306
rect 24050 14254 24052 14306
rect 23996 14252 24052 14254
rect 23436 13132 23492 13188
rect 21868 12348 21924 12404
rect 21084 12178 21140 12180
rect 21084 12126 21086 12178
rect 21086 12126 21138 12178
rect 21138 12126 21140 12178
rect 21084 12124 21140 12126
rect 20860 10444 20916 10500
rect 21980 12124 22036 12180
rect 21624 11002 21680 11004
rect 21624 10950 21626 11002
rect 21626 10950 21678 11002
rect 21678 10950 21680 11002
rect 21624 10948 21680 10950
rect 21728 11002 21784 11004
rect 21728 10950 21730 11002
rect 21730 10950 21782 11002
rect 21782 10950 21784 11002
rect 21728 10948 21784 10950
rect 21832 11002 21888 11004
rect 21832 10950 21834 11002
rect 21834 10950 21886 11002
rect 21886 10950 21888 11002
rect 21832 10948 21888 10950
rect 20636 9212 20692 9268
rect 21196 8092 21252 8148
rect 20412 7980 20468 8036
rect 17276 7532 17332 7588
rect 18222 7082 18278 7084
rect 18222 7030 18224 7082
rect 18224 7030 18276 7082
rect 18276 7030 18278 7082
rect 18222 7028 18278 7030
rect 18326 7082 18382 7084
rect 18326 7030 18328 7082
rect 18328 7030 18380 7082
rect 18380 7030 18382 7082
rect 18326 7028 18382 7030
rect 18430 7082 18486 7084
rect 18430 7030 18432 7082
rect 18432 7030 18484 7082
rect 18484 7030 18486 7082
rect 18430 7028 18486 7030
rect 20524 6636 20580 6692
rect 18844 6524 18900 6580
rect 18222 5514 18278 5516
rect 18222 5462 18224 5514
rect 18224 5462 18276 5514
rect 18276 5462 18278 5514
rect 18222 5460 18278 5462
rect 18326 5514 18382 5516
rect 18326 5462 18328 5514
rect 18328 5462 18380 5514
rect 18380 5462 18382 5514
rect 18326 5460 18382 5462
rect 18430 5514 18486 5516
rect 18430 5462 18432 5514
rect 18432 5462 18484 5514
rect 18484 5462 18486 5514
rect 18430 5460 18486 5462
rect 14820 4730 14876 4732
rect 14820 4678 14822 4730
rect 14822 4678 14874 4730
rect 14874 4678 14876 4730
rect 14820 4676 14876 4678
rect 14924 4730 14980 4732
rect 14924 4678 14926 4730
rect 14926 4678 14978 4730
rect 14978 4678 14980 4730
rect 14924 4676 14980 4678
rect 15028 4730 15084 4732
rect 15028 4678 15030 4730
rect 15030 4678 15082 4730
rect 15082 4678 15084 4730
rect 15028 4676 15084 4678
rect 14700 4338 14756 4340
rect 14700 4286 14702 4338
rect 14702 4286 14754 4338
rect 14754 4286 14756 4338
rect 14700 4284 14756 4286
rect 16940 4284 16996 4340
rect 16492 3500 16548 3556
rect 14820 3162 14876 3164
rect 14820 3110 14822 3162
rect 14822 3110 14874 3162
rect 14874 3110 14876 3162
rect 14820 3108 14876 3110
rect 14924 3162 14980 3164
rect 14924 3110 14926 3162
rect 14926 3110 14978 3162
rect 14978 3110 14980 3162
rect 14924 3108 14980 3110
rect 15028 3162 15084 3164
rect 15028 3110 15030 3162
rect 15030 3110 15082 3162
rect 15082 3110 15084 3162
rect 15028 3108 15084 3110
rect 17164 3554 17220 3556
rect 17164 3502 17166 3554
rect 17166 3502 17218 3554
rect 17218 3502 17220 3554
rect 17164 3500 17220 3502
rect 18222 3946 18278 3948
rect 18222 3894 18224 3946
rect 18224 3894 18276 3946
rect 18276 3894 18278 3946
rect 18222 3892 18278 3894
rect 18326 3946 18382 3948
rect 18326 3894 18328 3946
rect 18328 3894 18380 3946
rect 18380 3894 18382 3946
rect 18326 3892 18382 3894
rect 18430 3946 18486 3948
rect 18430 3894 18432 3946
rect 18432 3894 18484 3946
rect 18484 3894 18486 3946
rect 18430 3892 18486 3894
rect 19628 6412 19684 6468
rect 19404 5964 19460 6020
rect 19292 4450 19348 4452
rect 19292 4398 19294 4450
rect 19294 4398 19346 4450
rect 19346 4398 19348 4450
rect 19292 4396 19348 4398
rect 19516 3612 19572 3668
rect 18508 2716 18564 2772
rect 20188 3500 20244 3556
rect 20860 6018 20916 6020
rect 20860 5966 20862 6018
rect 20862 5966 20914 6018
rect 20914 5966 20916 6018
rect 20860 5964 20916 5966
rect 21084 5964 21140 6020
rect 21084 5628 21140 5684
rect 21624 9434 21680 9436
rect 21624 9382 21626 9434
rect 21626 9382 21678 9434
rect 21678 9382 21680 9434
rect 21624 9380 21680 9382
rect 21728 9434 21784 9436
rect 21728 9382 21730 9434
rect 21730 9382 21782 9434
rect 21782 9382 21784 9434
rect 21728 9380 21784 9382
rect 21832 9434 21888 9436
rect 21832 9382 21834 9434
rect 21834 9382 21886 9434
rect 21886 9382 21888 9434
rect 21832 9380 21888 9382
rect 22764 12124 22820 12180
rect 23548 12124 23604 12180
rect 23996 11676 24052 11732
rect 24220 12012 24276 12068
rect 22316 9212 22372 9268
rect 21980 8988 22036 9044
rect 21532 7980 21588 8036
rect 21624 7866 21680 7868
rect 21624 7814 21626 7866
rect 21626 7814 21678 7866
rect 21678 7814 21680 7866
rect 21624 7812 21680 7814
rect 21728 7866 21784 7868
rect 21728 7814 21730 7866
rect 21730 7814 21782 7866
rect 21782 7814 21784 7866
rect 21728 7812 21784 7814
rect 21832 7866 21888 7868
rect 21832 7814 21834 7866
rect 21834 7814 21886 7866
rect 21886 7814 21888 7866
rect 21832 7812 21888 7814
rect 23660 10386 23716 10388
rect 23660 10334 23662 10386
rect 23662 10334 23714 10386
rect 23714 10334 23716 10386
rect 23660 10332 23716 10334
rect 23548 9938 23604 9940
rect 23548 9886 23550 9938
rect 23550 9886 23602 9938
rect 23602 9886 23604 9938
rect 23548 9884 23604 9886
rect 23100 9212 23156 9268
rect 23548 9548 23604 9604
rect 22428 8930 22484 8932
rect 22428 8878 22430 8930
rect 22430 8878 22482 8930
rect 22482 8878 22484 8930
rect 22428 8876 22484 8878
rect 24556 10610 24612 10612
rect 24556 10558 24558 10610
rect 24558 10558 24610 10610
rect 24610 10558 24612 10610
rect 24556 10556 24612 10558
rect 24220 9212 24276 9268
rect 24332 8988 24388 9044
rect 24444 9884 24500 9940
rect 23996 8204 24052 8260
rect 23548 8146 23604 8148
rect 23548 8094 23550 8146
rect 23550 8094 23602 8146
rect 23602 8094 23604 8146
rect 23548 8092 23604 8094
rect 21532 6636 21588 6692
rect 24220 7308 24276 7364
rect 25026 13354 25082 13356
rect 25026 13302 25028 13354
rect 25028 13302 25080 13354
rect 25080 13302 25082 13354
rect 25026 13300 25082 13302
rect 25130 13354 25186 13356
rect 25130 13302 25132 13354
rect 25132 13302 25184 13354
rect 25184 13302 25186 13354
rect 25130 13300 25186 13302
rect 25234 13354 25290 13356
rect 25234 13302 25236 13354
rect 25236 13302 25288 13354
rect 25288 13302 25290 13354
rect 25234 13300 25290 13302
rect 25340 12066 25396 12068
rect 25340 12014 25342 12066
rect 25342 12014 25394 12066
rect 25394 12014 25396 12066
rect 25340 12012 25396 12014
rect 25026 11786 25082 11788
rect 25026 11734 25028 11786
rect 25028 11734 25080 11786
rect 25080 11734 25082 11786
rect 25026 11732 25082 11734
rect 25130 11786 25186 11788
rect 25130 11734 25132 11786
rect 25132 11734 25184 11786
rect 25184 11734 25186 11786
rect 25130 11732 25186 11734
rect 25234 11786 25290 11788
rect 25234 11734 25236 11786
rect 25236 11734 25288 11786
rect 25288 11734 25290 11786
rect 25234 11732 25290 11734
rect 25026 10218 25082 10220
rect 25026 10166 25028 10218
rect 25028 10166 25080 10218
rect 25080 10166 25082 10218
rect 25026 10164 25082 10166
rect 25130 10218 25186 10220
rect 25130 10166 25132 10218
rect 25132 10166 25184 10218
rect 25184 10166 25186 10218
rect 25130 10164 25186 10166
rect 25234 10218 25290 10220
rect 25234 10166 25236 10218
rect 25236 10166 25288 10218
rect 25288 10166 25290 10218
rect 25234 10164 25290 10166
rect 25788 16882 25844 16884
rect 25788 16830 25790 16882
rect 25790 16830 25842 16882
rect 25842 16830 25844 16882
rect 25788 16828 25844 16830
rect 25900 13970 25956 13972
rect 25900 13918 25902 13970
rect 25902 13918 25954 13970
rect 25954 13918 25956 13970
rect 25900 13916 25956 13918
rect 28140 16882 28196 16884
rect 28140 16830 28142 16882
rect 28142 16830 28194 16882
rect 28194 16830 28196 16882
rect 28140 16828 28196 16830
rect 27244 14700 27300 14756
rect 27468 15260 27524 15316
rect 26684 14530 26740 14532
rect 26684 14478 26686 14530
rect 26686 14478 26738 14530
rect 26738 14478 26740 14530
rect 26684 14476 26740 14478
rect 26908 14140 26964 14196
rect 26236 13634 26292 13636
rect 26236 13582 26238 13634
rect 26238 13582 26290 13634
rect 26290 13582 26292 13634
rect 26236 13580 26292 13582
rect 26124 13132 26180 13188
rect 26908 13468 26964 13524
rect 26236 12236 26292 12292
rect 25900 12066 25956 12068
rect 25900 12014 25902 12066
rect 25902 12014 25954 12066
rect 25954 12014 25956 12066
rect 25900 12012 25956 12014
rect 26796 11116 26852 11172
rect 26236 10498 26292 10500
rect 26236 10446 26238 10498
rect 26238 10446 26290 10498
rect 26290 10446 26292 10498
rect 26236 10444 26292 10446
rect 26236 9996 26292 10052
rect 24780 9212 24836 9268
rect 25026 8650 25082 8652
rect 25026 8598 25028 8650
rect 25028 8598 25080 8650
rect 25080 8598 25082 8650
rect 25026 8596 25082 8598
rect 25130 8650 25186 8652
rect 25130 8598 25132 8650
rect 25132 8598 25184 8650
rect 25184 8598 25186 8650
rect 25130 8596 25186 8598
rect 25234 8650 25290 8652
rect 25234 8598 25236 8650
rect 25236 8598 25288 8650
rect 25288 8598 25290 8650
rect 25234 8596 25290 8598
rect 24556 8258 24612 8260
rect 24556 8206 24558 8258
rect 24558 8206 24610 8258
rect 24610 8206 24612 8258
rect 24556 8204 24612 8206
rect 24556 7644 24612 7700
rect 24332 6636 24388 6692
rect 21980 6578 22036 6580
rect 21980 6526 21982 6578
rect 21982 6526 22034 6578
rect 22034 6526 22036 6578
rect 21980 6524 22036 6526
rect 22316 6466 22372 6468
rect 22316 6414 22318 6466
rect 22318 6414 22370 6466
rect 22370 6414 22372 6466
rect 22316 6412 22372 6414
rect 21624 6298 21680 6300
rect 21624 6246 21626 6298
rect 21626 6246 21678 6298
rect 21678 6246 21680 6298
rect 21624 6244 21680 6246
rect 21728 6298 21784 6300
rect 21728 6246 21730 6298
rect 21730 6246 21782 6298
rect 21782 6246 21784 6298
rect 21728 6244 21784 6246
rect 21832 6298 21888 6300
rect 21832 6246 21834 6298
rect 21834 6246 21886 6298
rect 21886 6246 21888 6298
rect 21832 6244 21888 6246
rect 23100 6076 23156 6132
rect 22540 6018 22596 6020
rect 22540 5966 22542 6018
rect 22542 5966 22594 6018
rect 22594 5966 22596 6018
rect 22540 5964 22596 5966
rect 21084 4508 21140 4564
rect 23324 5234 23380 5236
rect 23324 5182 23326 5234
rect 23326 5182 23378 5234
rect 23378 5182 23380 5234
rect 23324 5180 23380 5182
rect 21196 4284 21252 4340
rect 21308 5068 21364 5124
rect 22316 5010 22372 5012
rect 22316 4958 22318 5010
rect 22318 4958 22370 5010
rect 22370 4958 22372 5010
rect 22316 4956 22372 4958
rect 20412 4226 20468 4228
rect 20412 4174 20414 4226
rect 20414 4174 20466 4226
rect 20466 4174 20468 4226
rect 20412 4172 20468 4174
rect 21624 4730 21680 4732
rect 21624 4678 21626 4730
rect 21626 4678 21678 4730
rect 21678 4678 21680 4730
rect 21624 4676 21680 4678
rect 21728 4730 21784 4732
rect 21728 4678 21730 4730
rect 21730 4678 21782 4730
rect 21782 4678 21784 4730
rect 21728 4676 21784 4678
rect 21832 4730 21888 4732
rect 21832 4678 21834 4730
rect 21834 4678 21886 4730
rect 21886 4678 21888 4730
rect 21832 4676 21888 4678
rect 24668 6636 24724 6692
rect 24556 5122 24612 5124
rect 24556 5070 24558 5122
rect 24558 5070 24610 5122
rect 24610 5070 24612 5122
rect 24556 5068 24612 5070
rect 24444 4844 24500 4900
rect 24780 4956 24836 5012
rect 22652 4396 22708 4452
rect 21644 4338 21700 4340
rect 21644 4286 21646 4338
rect 21646 4286 21698 4338
rect 21698 4286 21700 4338
rect 21644 4284 21700 4286
rect 20300 3388 20356 3444
rect 21084 3442 21140 3444
rect 21084 3390 21086 3442
rect 21086 3390 21138 3442
rect 21138 3390 21140 3442
rect 21084 3388 21140 3390
rect 22316 3554 22372 3556
rect 22316 3502 22318 3554
rect 22318 3502 22370 3554
rect 22370 3502 22372 3554
rect 22316 3500 22372 3502
rect 25340 7698 25396 7700
rect 25340 7646 25342 7698
rect 25342 7646 25394 7698
rect 25394 7646 25396 7698
rect 25340 7644 25396 7646
rect 25026 7082 25082 7084
rect 25026 7030 25028 7082
rect 25028 7030 25080 7082
rect 25080 7030 25082 7082
rect 25026 7028 25082 7030
rect 25130 7082 25186 7084
rect 25130 7030 25132 7082
rect 25132 7030 25184 7082
rect 25184 7030 25186 7082
rect 25130 7028 25186 7030
rect 25234 7082 25290 7084
rect 25234 7030 25236 7082
rect 25236 7030 25288 7082
rect 25288 7030 25290 7082
rect 25234 7028 25290 7030
rect 26348 7644 26404 7700
rect 26236 7362 26292 7364
rect 26236 7310 26238 7362
rect 26238 7310 26290 7362
rect 26290 7310 26292 7362
rect 26236 7308 26292 7310
rect 27020 11506 27076 11508
rect 27020 11454 27022 11506
rect 27022 11454 27074 11506
rect 27074 11454 27076 11506
rect 27020 11452 27076 11454
rect 27020 10332 27076 10388
rect 27692 14812 27748 14868
rect 27580 14476 27636 14532
rect 27804 14252 27860 14308
rect 28028 14140 28084 14196
rect 27356 13468 27412 13524
rect 27244 11452 27300 11508
rect 27244 11282 27300 11284
rect 27244 11230 27246 11282
rect 27246 11230 27298 11282
rect 27298 11230 27300 11282
rect 27244 11228 27300 11230
rect 27244 10556 27300 10612
rect 28140 12124 28196 12180
rect 27580 11282 27636 11284
rect 27580 11230 27582 11282
rect 27582 11230 27634 11282
rect 27634 11230 27636 11282
rect 27580 11228 27636 11230
rect 27692 11170 27748 11172
rect 27692 11118 27694 11170
rect 27694 11118 27746 11170
rect 27746 11118 27748 11170
rect 27692 11116 27748 11118
rect 28428 15706 28484 15708
rect 28428 15654 28430 15706
rect 28430 15654 28482 15706
rect 28482 15654 28484 15706
rect 28428 15652 28484 15654
rect 28532 15706 28588 15708
rect 28532 15654 28534 15706
rect 28534 15654 28586 15706
rect 28586 15654 28588 15706
rect 28532 15652 28588 15654
rect 28636 15706 28692 15708
rect 28636 15654 28638 15706
rect 28638 15654 28690 15706
rect 28690 15654 28692 15706
rect 28636 15652 28692 15654
rect 28428 14138 28484 14140
rect 28428 14086 28430 14138
rect 28430 14086 28482 14138
rect 28482 14086 28484 14138
rect 28428 14084 28484 14086
rect 28532 14138 28588 14140
rect 28532 14086 28534 14138
rect 28534 14086 28586 14138
rect 28586 14086 28588 14138
rect 28532 14084 28588 14086
rect 28636 14138 28692 14140
rect 28636 14086 28638 14138
rect 28638 14086 28690 14138
rect 28690 14086 28692 14138
rect 28636 14084 28692 14086
rect 28428 12570 28484 12572
rect 28428 12518 28430 12570
rect 28430 12518 28482 12570
rect 28482 12518 28484 12570
rect 28428 12516 28484 12518
rect 28532 12570 28588 12572
rect 28532 12518 28534 12570
rect 28534 12518 28586 12570
rect 28586 12518 28588 12570
rect 28532 12516 28588 12518
rect 28636 12570 28692 12572
rect 28636 12518 28638 12570
rect 28638 12518 28690 12570
rect 28690 12518 28692 12570
rect 28636 12516 28692 12518
rect 28428 11002 28484 11004
rect 28428 10950 28430 11002
rect 28430 10950 28482 11002
rect 28482 10950 28484 11002
rect 28428 10948 28484 10950
rect 28532 11002 28588 11004
rect 28532 10950 28534 11002
rect 28534 10950 28586 11002
rect 28586 10950 28588 11002
rect 28532 10948 28588 10950
rect 28636 11002 28692 11004
rect 28636 10950 28638 11002
rect 28638 10950 28690 11002
rect 28690 10950 28692 11002
rect 28636 10948 28692 10950
rect 28140 9266 28196 9268
rect 28140 9214 28142 9266
rect 28142 9214 28194 9266
rect 28194 9214 28196 9266
rect 28140 9212 28196 9214
rect 28428 9434 28484 9436
rect 28428 9382 28430 9434
rect 28430 9382 28482 9434
rect 28482 9382 28484 9434
rect 28428 9380 28484 9382
rect 28532 9434 28588 9436
rect 28532 9382 28534 9434
rect 28534 9382 28586 9434
rect 28586 9382 28588 9434
rect 28532 9380 28588 9382
rect 28636 9434 28692 9436
rect 28636 9382 28638 9434
rect 28638 9382 28690 9434
rect 28690 9382 28692 9434
rect 28636 9380 28692 9382
rect 28428 7866 28484 7868
rect 28428 7814 28430 7866
rect 28430 7814 28482 7866
rect 28482 7814 28484 7866
rect 28428 7812 28484 7814
rect 28532 7866 28588 7868
rect 28532 7814 28534 7866
rect 28534 7814 28586 7866
rect 28586 7814 28588 7866
rect 28532 7812 28588 7814
rect 28636 7866 28692 7868
rect 28636 7814 28638 7866
rect 28638 7814 28690 7866
rect 28690 7814 28692 7866
rect 28636 7812 28692 7814
rect 27692 6690 27748 6692
rect 27692 6638 27694 6690
rect 27694 6638 27746 6690
rect 27746 6638 27748 6690
rect 27692 6636 27748 6638
rect 25026 5514 25082 5516
rect 25026 5462 25028 5514
rect 25028 5462 25080 5514
rect 25080 5462 25082 5514
rect 25026 5460 25082 5462
rect 25130 5514 25186 5516
rect 25130 5462 25132 5514
rect 25132 5462 25184 5514
rect 25184 5462 25186 5514
rect 25130 5460 25186 5462
rect 25234 5514 25290 5516
rect 25234 5462 25236 5514
rect 25236 5462 25288 5514
rect 25288 5462 25290 5514
rect 25234 5460 25290 5462
rect 25228 5180 25284 5236
rect 25340 5068 25396 5124
rect 26236 4844 26292 4900
rect 26124 4508 26180 4564
rect 24892 4396 24948 4452
rect 25026 3946 25082 3948
rect 25026 3894 25028 3946
rect 25028 3894 25080 3946
rect 25080 3894 25082 3946
rect 25026 3892 25082 3894
rect 25130 3946 25186 3948
rect 25130 3894 25132 3946
rect 25132 3894 25184 3946
rect 25184 3894 25186 3946
rect 25130 3892 25186 3894
rect 25234 3946 25290 3948
rect 25234 3894 25236 3946
rect 25236 3894 25288 3946
rect 25288 3894 25290 3946
rect 25234 3892 25290 3894
rect 23100 3666 23156 3668
rect 23100 3614 23102 3666
rect 23102 3614 23154 3666
rect 23154 3614 23156 3666
rect 23100 3612 23156 3614
rect 28428 6298 28484 6300
rect 28428 6246 28430 6298
rect 28430 6246 28482 6298
rect 28482 6246 28484 6298
rect 28428 6244 28484 6246
rect 28532 6298 28588 6300
rect 28532 6246 28534 6298
rect 28534 6246 28586 6298
rect 28586 6246 28588 6298
rect 28532 6244 28588 6246
rect 28636 6298 28692 6300
rect 28636 6246 28638 6298
rect 28638 6246 28690 6298
rect 28690 6246 28692 6298
rect 28636 6244 28692 6246
rect 27244 4450 27300 4452
rect 27244 4398 27246 4450
rect 27246 4398 27298 4450
rect 27298 4398 27300 4450
rect 27244 4396 27300 4398
rect 28476 4844 28532 4900
rect 28428 4730 28484 4732
rect 28428 4678 28430 4730
rect 28430 4678 28482 4730
rect 28482 4678 28484 4730
rect 28428 4676 28484 4678
rect 28532 4730 28588 4732
rect 28532 4678 28534 4730
rect 28534 4678 28586 4730
rect 28586 4678 28588 4730
rect 28532 4676 28588 4678
rect 28636 4730 28692 4732
rect 28636 4678 28638 4730
rect 28638 4678 28690 4730
rect 28690 4678 28692 4730
rect 28636 4676 28692 4678
rect 28140 3388 28196 3444
rect 21624 3162 21680 3164
rect 21624 3110 21626 3162
rect 21626 3110 21678 3162
rect 21678 3110 21680 3162
rect 21624 3108 21680 3110
rect 21728 3162 21784 3164
rect 21728 3110 21730 3162
rect 21730 3110 21782 3162
rect 21782 3110 21784 3162
rect 21728 3108 21784 3110
rect 21832 3162 21888 3164
rect 21832 3110 21834 3162
rect 21834 3110 21886 3162
rect 21886 3110 21888 3162
rect 21832 3108 21888 3110
rect 28428 3162 28484 3164
rect 28428 3110 28430 3162
rect 28430 3110 28482 3162
rect 28482 3110 28484 3162
rect 28428 3108 28484 3110
rect 28532 3162 28588 3164
rect 28532 3110 28534 3162
rect 28534 3110 28586 3162
rect 28586 3110 28588 3162
rect 28532 3108 28588 3110
rect 28636 3162 28692 3164
rect 28636 3110 28638 3162
rect 28638 3110 28690 3162
rect 28690 3110 28692 3162
rect 28636 3108 28692 3110
<< metal3 >>
rect 29200 26964 30000 26992
rect 28140 26908 30000 26964
rect 28140 26852 28196 26908
rect 29200 26880 30000 26908
rect 18162 26796 18172 26852
rect 18228 26796 18956 26852
rect 19012 26796 19022 26852
rect 21522 26796 21532 26852
rect 21588 26796 22764 26852
rect 22820 26796 22830 26852
rect 28130 26796 28140 26852
rect 28196 26796 28206 26852
rect 8006 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8290 26684
rect 14810 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15094 26684
rect 21614 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21898 26684
rect 28418 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28702 26684
rect 13346 26460 13356 26516
rect 13412 26460 14028 26516
rect 14084 26460 14094 26516
rect 17602 26460 17612 26516
rect 17668 26460 19068 26516
rect 19124 26460 19134 26516
rect 19506 26460 19516 26516
rect 19572 26460 21196 26516
rect 21252 26460 21262 26516
rect 22866 26460 22876 26516
rect 22932 26460 23884 26516
rect 23940 26460 23950 26516
rect 29200 26292 30000 26320
rect 12898 26236 12908 26292
rect 12964 26236 13692 26292
rect 13748 26236 13758 26292
rect 16258 26236 16268 26292
rect 16324 26236 17164 26292
rect 17220 26236 17230 26292
rect 26226 26236 26236 26292
rect 26292 26236 30000 26292
rect 29200 26208 30000 26236
rect 4604 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4888 25900
rect 11408 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11692 25900
rect 18212 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18496 25900
rect 25016 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25300 25900
rect 12786 25676 12796 25732
rect 12852 25676 13916 25732
rect 13972 25676 13982 25732
rect 29200 25620 30000 25648
rect 16482 25564 16492 25620
rect 16548 25564 22652 25620
rect 22708 25564 22718 25620
rect 27682 25564 27692 25620
rect 27748 25564 30000 25620
rect 29200 25536 30000 25564
rect 19618 25452 19628 25508
rect 19684 25452 20188 25508
rect 20244 25452 20254 25508
rect 20850 25452 20860 25508
rect 20916 25452 21308 25508
rect 21364 25452 22204 25508
rect 22260 25452 22270 25508
rect 27122 25452 27132 25508
rect 27188 25452 28140 25508
rect 28196 25452 28206 25508
rect 19058 25340 19068 25396
rect 19124 25340 20748 25396
rect 20804 25340 20814 25396
rect 1698 25228 1708 25284
rect 1764 25228 1774 25284
rect 9538 25228 9548 25284
rect 9604 25228 10332 25284
rect 10388 25228 10398 25284
rect 11330 25228 11340 25284
rect 11396 25228 12796 25284
rect 12852 25228 12862 25284
rect 18946 25228 18956 25284
rect 19012 25228 19964 25284
rect 20020 25228 20030 25284
rect 21410 25228 21420 25284
rect 21476 25228 21980 25284
rect 22036 25228 22046 25284
rect 27458 25228 27468 25284
rect 27524 25228 27534 25284
rect 0 24948 800 24976
rect 1708 24948 1764 25228
rect 8006 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8290 25116
rect 14810 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15094 25116
rect 21614 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21898 25116
rect 0 24892 1764 24948
rect 27468 24948 27524 25228
rect 28418 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28702 25116
rect 29200 24948 30000 24976
rect 27468 24892 30000 24948
rect 0 24864 800 24892
rect 29200 24864 30000 24892
rect 4604 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4888 24332
rect 11408 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11692 24332
rect 18212 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18496 24332
rect 25016 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25300 24332
rect 29200 24276 30000 24304
rect 28130 24220 28140 24276
rect 28196 24220 30000 24276
rect 29200 24192 30000 24220
rect 27682 23660 27692 23716
rect 27748 23660 28868 23716
rect 28812 23604 28868 23660
rect 29200 23604 30000 23632
rect 28812 23548 30000 23604
rect 8006 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8290 23548
rect 14810 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15094 23548
rect 21614 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21898 23548
rect 28418 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28702 23548
rect 29200 23520 30000 23548
rect 26898 22988 26908 23044
rect 26964 22988 28140 23044
rect 28196 22988 28206 23044
rect 29200 22932 30000 22960
rect 28242 22876 28252 22932
rect 28308 22876 30000 22932
rect 29200 22848 30000 22876
rect 4604 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4888 22764
rect 11408 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11692 22764
rect 18212 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18496 22764
rect 25016 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25300 22764
rect 29200 22260 30000 22288
rect 28018 22204 28028 22260
rect 28084 22204 30000 22260
rect 29200 22176 30000 22204
rect 8006 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8290 21980
rect 14810 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15094 21980
rect 21614 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21898 21980
rect 28418 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28702 21980
rect 15698 21756 15708 21812
rect 15764 21756 18620 21812
rect 18676 21756 18686 21812
rect 16370 21644 16380 21700
rect 16436 21644 18732 21700
rect 18788 21644 18798 21700
rect 24882 21644 24892 21700
rect 24948 21644 27244 21700
rect 27300 21644 27310 21700
rect 29200 21588 30000 21616
rect 28130 21532 28140 21588
rect 28196 21532 30000 21588
rect 29200 21504 30000 21532
rect 23650 21420 23660 21476
rect 23716 21420 26236 21476
rect 26292 21420 26302 21476
rect 4604 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4888 21196
rect 11408 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11692 21196
rect 18212 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18496 21196
rect 25016 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25300 21196
rect 26114 20636 26124 20692
rect 26180 20636 26908 20692
rect 26964 20636 26974 20692
rect 8006 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8290 20412
rect 14810 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15094 20412
rect 21614 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21898 20412
rect 28418 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28702 20412
rect 14130 20076 14140 20132
rect 14196 20076 16268 20132
rect 16324 20076 16334 20132
rect 22418 20076 22428 20132
rect 22484 20076 27244 20132
rect 27300 20076 27310 20132
rect 25890 19964 25900 20020
rect 25956 19964 27356 20020
rect 27412 19964 27422 20020
rect 8754 19852 8764 19908
rect 8820 19852 10668 19908
rect 10724 19852 10734 19908
rect 14018 19852 14028 19908
rect 14084 19852 15260 19908
rect 15316 19852 15326 19908
rect 21858 19852 21868 19908
rect 21924 19852 26236 19908
rect 26292 19852 26302 19908
rect 0 19572 800 19600
rect 4604 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4888 19628
rect 11408 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11692 19628
rect 18212 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18496 19628
rect 25016 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25300 19628
rect 0 19516 4228 19572
rect 0 19488 800 19516
rect 4172 19460 4228 19516
rect 4172 19404 14588 19460
rect 14644 19404 14654 19460
rect 15474 19292 15484 19348
rect 15540 19292 18284 19348
rect 18340 19292 18350 19348
rect 18946 19180 18956 19236
rect 19012 19180 21420 19236
rect 21476 19180 22764 19236
rect 22820 19180 22830 19236
rect 17042 19068 17052 19124
rect 17108 19068 19292 19124
rect 19348 19068 19358 19124
rect 26898 19068 26908 19124
rect 26964 19068 27692 19124
rect 27748 19068 27758 19124
rect 8006 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8290 18844
rect 14810 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15094 18844
rect 21614 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21898 18844
rect 28418 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28702 18844
rect 8306 18620 8316 18676
rect 8372 18620 9660 18676
rect 9716 18620 9726 18676
rect 18610 18620 18620 18676
rect 18676 18620 23212 18676
rect 23268 18620 23278 18676
rect 5954 18508 5964 18564
rect 6020 18508 8428 18564
rect 8484 18508 8494 18564
rect 18396 18508 18956 18564
rect 19012 18508 19022 18564
rect 22754 18508 22764 18564
rect 22820 18508 23604 18564
rect 18396 18452 18452 18508
rect 15026 18396 15036 18452
rect 15092 18396 17500 18452
rect 17556 18396 17948 18452
rect 18004 18396 18452 18452
rect 23548 18452 23604 18508
rect 23548 18396 24892 18452
rect 24948 18396 24958 18452
rect 5282 18284 5292 18340
rect 5348 18284 7196 18340
rect 7252 18284 7262 18340
rect 14466 18284 14476 18340
rect 14532 18284 15372 18340
rect 15428 18284 16044 18340
rect 16100 18284 16716 18340
rect 16772 18284 16782 18340
rect 17826 18284 17836 18340
rect 17892 18284 22204 18340
rect 22260 18284 22270 18340
rect 24098 18284 24108 18340
rect 24164 18284 25900 18340
rect 25956 18284 25966 18340
rect 10322 18172 10332 18228
rect 10388 18172 11676 18228
rect 11732 18172 11742 18228
rect 20962 18172 20972 18228
rect 21028 18172 23548 18228
rect 23604 18172 23614 18228
rect 4604 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4888 18060
rect 11408 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11692 18060
rect 18212 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18496 18060
rect 25016 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25300 18060
rect 8372 17948 8652 18004
rect 8708 17948 8718 18004
rect 8372 17780 8428 17948
rect 7298 17724 7308 17780
rect 7364 17724 8428 17780
rect 19394 17724 19404 17780
rect 19460 17724 22316 17780
rect 22372 17724 22382 17780
rect 2258 17612 2268 17668
rect 2324 17612 14364 17668
rect 14420 17612 14430 17668
rect 16706 17612 16716 17668
rect 16772 17612 17612 17668
rect 17668 17612 19628 17668
rect 19684 17612 20524 17668
rect 20580 17612 21420 17668
rect 21476 17612 21868 17668
rect 21924 17612 24220 17668
rect 24276 17612 24286 17668
rect 11218 17500 11228 17556
rect 11284 17500 12012 17556
rect 12068 17500 12078 17556
rect 8006 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8290 17276
rect 14810 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15094 17276
rect 21614 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21898 17276
rect 28418 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28702 17276
rect 24434 17052 24444 17108
rect 24500 17052 25340 17108
rect 25396 17052 27132 17108
rect 27188 17052 27198 17108
rect 14130 16940 14140 16996
rect 14196 16940 16380 16996
rect 16436 16940 16446 16996
rect 23426 16940 23436 16996
rect 23492 16940 24220 16996
rect 24276 16940 24286 16996
rect 0 16884 800 16912
rect 0 16828 1708 16884
rect 1764 16828 1774 16884
rect 2482 16828 2492 16884
rect 2548 16828 4620 16884
rect 4676 16828 5460 16884
rect 7410 16828 7420 16884
rect 7476 16828 8988 16884
rect 9044 16828 9772 16884
rect 9828 16828 9838 16884
rect 18284 16828 18956 16884
rect 19012 16828 19740 16884
rect 19796 16828 20188 16884
rect 24882 16828 24892 16884
rect 24948 16828 25788 16884
rect 25844 16828 28140 16884
rect 28196 16828 28206 16884
rect 0 16800 800 16828
rect 5404 16772 5460 16828
rect 18284 16772 18340 16828
rect 20132 16772 20188 16828
rect 5404 16716 5516 16772
rect 5572 16716 5582 16772
rect 10658 16716 10668 16772
rect 10724 16716 13468 16772
rect 13524 16716 13534 16772
rect 14018 16716 14028 16772
rect 14084 16716 15372 16772
rect 15428 16716 15438 16772
rect 15698 16716 15708 16772
rect 15764 16716 18284 16772
rect 18340 16716 18350 16772
rect 20132 16716 20300 16772
rect 20356 16716 20366 16772
rect 11106 16604 11116 16660
rect 11172 16604 18620 16660
rect 18676 16604 18686 16660
rect 4604 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4888 16492
rect 11408 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11692 16492
rect 18212 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18496 16492
rect 25016 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25300 16492
rect 16258 16156 16268 16212
rect 16324 16156 18284 16212
rect 18340 16156 18350 16212
rect 5506 16044 5516 16100
rect 5572 16044 6636 16100
rect 6692 16044 7756 16100
rect 7812 16044 7822 16100
rect 2818 15932 2828 15988
rect 2884 15932 4732 15988
rect 4788 15932 4798 15988
rect 12562 15932 12572 15988
rect 12628 15932 15708 15988
rect 15764 15932 15774 15988
rect 17042 15932 17052 15988
rect 17108 15932 19292 15988
rect 19348 15932 19358 15988
rect 19954 15932 19964 15988
rect 20020 15932 23212 15988
rect 23268 15932 23278 15988
rect 16482 15820 16492 15876
rect 16548 15820 20300 15876
rect 20356 15820 20366 15876
rect 8006 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8290 15708
rect 14810 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15094 15708
rect 21614 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21898 15708
rect 28418 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28702 15708
rect 20514 15484 20524 15540
rect 20580 15484 21756 15540
rect 21812 15484 24892 15540
rect 24948 15484 24958 15540
rect 4162 15372 4172 15428
rect 4228 15372 6748 15428
rect 6804 15372 6814 15428
rect 7858 15372 7868 15428
rect 7924 15372 9324 15428
rect 9380 15372 10444 15428
rect 10500 15372 10510 15428
rect 12786 15372 12796 15428
rect 12852 15372 13468 15428
rect 13524 15372 13534 15428
rect 14354 15372 14364 15428
rect 14420 15372 14700 15428
rect 14756 15372 15148 15428
rect 15204 15372 15214 15428
rect 19282 15372 19292 15428
rect 19348 15372 23660 15428
rect 23716 15372 23726 15428
rect 23986 15372 23996 15428
rect 24052 15372 25340 15428
rect 25396 15372 25406 15428
rect 4050 15260 4060 15316
rect 4116 15260 5068 15316
rect 5124 15260 5134 15316
rect 18386 15260 18396 15316
rect 18452 15260 20188 15316
rect 21410 15260 21420 15316
rect 21476 15260 27468 15316
rect 27524 15260 27534 15316
rect 20132 15204 20188 15260
rect 20132 15148 22652 15204
rect 22708 15148 22718 15204
rect 5282 15036 5292 15092
rect 5348 15036 6188 15092
rect 6244 15036 6254 15092
rect 4604 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4888 14924
rect 11408 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11692 14924
rect 18212 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18496 14924
rect 25016 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25300 14924
rect 29200 14868 30000 14896
rect 7970 14812 7980 14868
rect 8036 14812 9660 14868
rect 9716 14812 9726 14868
rect 27682 14812 27692 14868
rect 27748 14812 30000 14868
rect 29200 14784 30000 14812
rect 23762 14700 23772 14756
rect 23828 14700 27244 14756
rect 27300 14700 27310 14756
rect 15138 14476 15148 14532
rect 15204 14476 15820 14532
rect 15876 14476 17836 14532
rect 17892 14476 17902 14532
rect 24882 14476 24892 14532
rect 24948 14476 26684 14532
rect 26740 14476 27580 14532
rect 27636 14476 27646 14532
rect 4946 14364 4956 14420
rect 5012 14364 6076 14420
rect 6132 14364 6142 14420
rect 8978 14364 8988 14420
rect 9044 14364 11900 14420
rect 11956 14364 12796 14420
rect 12852 14364 13916 14420
rect 13972 14364 13982 14420
rect 3042 14252 3052 14308
rect 3108 14252 6636 14308
rect 6692 14252 6702 14308
rect 7410 14252 7420 14308
rect 7476 14252 8652 14308
rect 8708 14252 8718 14308
rect 19730 14252 19740 14308
rect 19796 14252 20636 14308
rect 20692 14252 21868 14308
rect 21924 14252 22316 14308
rect 22372 14252 22382 14308
rect 23986 14252 23996 14308
rect 24052 14252 27804 14308
rect 27860 14252 27870 14308
rect 25900 14140 26908 14196
rect 26964 14140 28028 14196
rect 28084 14140 28094 14196
rect 8006 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8290 14140
rect 14810 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15094 14140
rect 21614 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21898 14140
rect 25900 13972 25956 14140
rect 28418 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28702 14140
rect 22642 13916 22652 13972
rect 22708 13916 25900 13972
rect 25956 13916 25966 13972
rect 6402 13580 6412 13636
rect 6468 13580 8652 13636
rect 8708 13580 8988 13636
rect 9044 13580 9054 13636
rect 14242 13580 14252 13636
rect 14308 13580 18396 13636
rect 18452 13580 18462 13636
rect 20738 13580 20748 13636
rect 20804 13580 26236 13636
rect 26292 13580 26302 13636
rect 8754 13468 8764 13524
rect 8820 13468 11116 13524
rect 11172 13468 11182 13524
rect 26898 13468 26908 13524
rect 26964 13468 27356 13524
rect 27412 13468 27422 13524
rect 4604 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4888 13356
rect 11408 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11692 13356
rect 18212 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18496 13356
rect 25016 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25300 13356
rect 12786 13132 12796 13188
rect 12852 13132 19404 13188
rect 19460 13132 19470 13188
rect 23426 13132 23436 13188
rect 23492 13132 26124 13188
rect 26180 13132 26190 13188
rect 14466 13020 14476 13076
rect 14532 13020 20076 13076
rect 20132 13020 20142 13076
rect 4050 12908 4060 12964
rect 4116 12908 9660 12964
rect 9716 12908 9726 12964
rect 6066 12796 6076 12852
rect 6132 12796 7084 12852
rect 7140 12796 7150 12852
rect 3714 12684 3724 12740
rect 3780 12684 5852 12740
rect 5908 12684 6524 12740
rect 6580 12684 6590 12740
rect 8006 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8290 12572
rect 14810 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15094 12572
rect 21614 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21898 12572
rect 28418 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28702 12572
rect 20066 12348 20076 12404
rect 20132 12348 21868 12404
rect 21924 12348 21934 12404
rect 20402 12236 20412 12292
rect 20468 12236 26236 12292
rect 26292 12236 26302 12292
rect 0 12180 800 12208
rect 0 12124 1820 12180
rect 1876 12124 1886 12180
rect 19618 12124 19628 12180
rect 19684 12124 20300 12180
rect 20356 12124 21084 12180
rect 21140 12124 21980 12180
rect 22036 12124 22764 12180
rect 22820 12124 23548 12180
rect 23604 12124 23614 12180
rect 26852 12124 28140 12180
rect 28196 12124 28206 12180
rect 0 12096 800 12124
rect 26852 12068 26908 12124
rect 7868 12012 8428 12068
rect 8484 12012 8494 12068
rect 8652 12012 8876 12068
rect 8932 12012 8942 12068
rect 24210 12012 24220 12068
rect 24276 12012 25340 12068
rect 25396 12012 25900 12068
rect 25956 12012 26908 12068
rect 3042 11900 3052 11956
rect 3108 11900 7196 11956
rect 7252 11900 7262 11956
rect 7868 11844 7924 12012
rect 8652 11844 8708 12012
rect 7756 11788 7924 11844
rect 7980 11788 8708 11844
rect 4604 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4888 11788
rect 7756 11620 7812 11788
rect 7980 11732 8036 11788
rect 11408 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11692 11788
rect 18212 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18496 11788
rect 25016 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25300 11788
rect 7970 11676 7980 11732
rect 8036 11676 8046 11732
rect 8418 11676 8428 11732
rect 8484 11676 10108 11732
rect 10164 11676 10668 11732
rect 10724 11676 10734 11732
rect 23986 11676 23996 11732
rect 24052 11676 24062 11732
rect 4386 11564 4396 11620
rect 4452 11564 7812 11620
rect 8428 11396 8484 11676
rect 23996 11508 24052 11676
rect 18050 11452 18060 11508
rect 18116 11452 20188 11508
rect 20244 11452 20254 11508
rect 23996 11452 27020 11508
rect 27076 11452 27086 11508
rect 27234 11452 27244 11508
rect 27300 11452 27310 11508
rect 27244 11396 27300 11452
rect 5618 11340 5628 11396
rect 5684 11340 8484 11396
rect 10322 11340 10332 11396
rect 10388 11340 14588 11396
rect 14644 11340 14654 11396
rect 19170 11340 19180 11396
rect 19236 11340 27300 11396
rect 18610 11228 18620 11284
rect 18676 11228 19404 11284
rect 19460 11228 19470 11284
rect 27234 11228 27244 11284
rect 27300 11228 27580 11284
rect 27636 11228 27646 11284
rect 10098 11116 10108 11172
rect 10164 11116 11900 11172
rect 11956 11116 11966 11172
rect 26786 11116 26796 11172
rect 26852 11116 27692 11172
rect 27748 11116 27758 11172
rect 8006 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8290 11004
rect 14810 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15094 11004
rect 21614 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21898 11004
rect 28418 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28702 11004
rect 8306 10780 8316 10836
rect 8372 10780 11116 10836
rect 11172 10780 11182 10836
rect 15586 10780 15596 10836
rect 15652 10780 16380 10836
rect 16436 10780 16446 10836
rect 10658 10556 10668 10612
rect 10724 10556 12460 10612
rect 12516 10556 12526 10612
rect 24546 10556 24556 10612
rect 24612 10556 27244 10612
rect 27300 10556 27310 10612
rect 11218 10444 11228 10500
rect 11284 10444 13020 10500
rect 13076 10444 13086 10500
rect 15092 10444 16716 10500
rect 16772 10444 17500 10500
rect 17556 10444 17566 10500
rect 20850 10444 20860 10500
rect 20916 10444 26236 10500
rect 26292 10444 26302 10500
rect 1810 10332 1820 10388
rect 1876 10332 2492 10388
rect 2548 10332 5628 10388
rect 5684 10332 5694 10388
rect 4604 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4888 10220
rect 11408 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11692 10220
rect 15092 10164 15148 10444
rect 23650 10332 23660 10388
rect 23716 10332 27020 10388
rect 27076 10332 27086 10388
rect 18212 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18496 10220
rect 25016 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25300 10220
rect 12898 10108 12908 10164
rect 12964 10108 15148 10164
rect 15204 10108 15214 10164
rect 16258 9996 16268 10052
rect 16324 9996 26236 10052
rect 26292 9996 26302 10052
rect 19730 9884 19740 9940
rect 19796 9884 20300 9940
rect 20356 9884 23548 9940
rect 23604 9884 24444 9940
rect 24500 9884 24510 9940
rect 11106 9772 11116 9828
rect 11172 9772 12348 9828
rect 12404 9772 12414 9828
rect 2370 9660 2380 9716
rect 2436 9660 4284 9716
rect 4340 9660 4350 9716
rect 18610 9660 18620 9716
rect 18676 9660 19404 9716
rect 19460 9660 19470 9716
rect 19170 9548 19180 9604
rect 19236 9548 23548 9604
rect 23604 9548 23614 9604
rect 8006 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8290 9436
rect 14810 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15094 9436
rect 21614 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21898 9436
rect 28418 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28702 9436
rect 20626 9212 20636 9268
rect 20692 9212 22316 9268
rect 22372 9212 22382 9268
rect 23090 9212 23100 9268
rect 23156 9212 24220 9268
rect 24276 9212 24286 9268
rect 24770 9212 24780 9268
rect 24836 9212 28140 9268
rect 28196 9212 28206 9268
rect 9314 9100 9324 9156
rect 9380 9100 10108 9156
rect 10164 9100 10174 9156
rect 11442 8988 11452 9044
rect 11508 8988 13244 9044
rect 13300 8988 13310 9044
rect 15698 8988 15708 9044
rect 15764 8988 17500 9044
rect 17556 8988 19292 9044
rect 19348 8988 19358 9044
rect 21970 8988 21980 9044
rect 22036 8988 24332 9044
rect 24388 8988 24398 9044
rect 6066 8876 6076 8932
rect 6132 8876 7532 8932
rect 7588 8876 7598 8932
rect 18162 8876 18172 8932
rect 18228 8876 22428 8932
rect 22484 8876 22494 8932
rect 4604 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4888 8652
rect 11408 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11692 8652
rect 18212 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18496 8652
rect 25016 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25300 8652
rect 5058 8428 5068 8484
rect 5124 8428 6076 8484
rect 6132 8428 6524 8484
rect 6580 8428 6590 8484
rect 2818 8316 2828 8372
rect 2884 8316 3612 8372
rect 3668 8316 3678 8372
rect 4722 8316 4732 8372
rect 4788 8316 7420 8372
rect 7476 8316 7486 8372
rect 16146 8316 16156 8372
rect 16212 8316 17612 8372
rect 17668 8316 17678 8372
rect 12450 8204 12460 8260
rect 12516 8204 14476 8260
rect 14532 8204 14542 8260
rect 23986 8204 23996 8260
rect 24052 8204 24556 8260
rect 24612 8204 24622 8260
rect 1586 8092 1596 8148
rect 1652 8092 2492 8148
rect 2548 8092 2558 8148
rect 16370 8092 16380 8148
rect 16436 8092 18620 8148
rect 18676 8092 18686 8148
rect 21186 8092 21196 8148
rect 21252 8092 23548 8148
rect 23604 8092 23614 8148
rect 10098 7980 10108 8036
rect 10164 7980 12460 8036
rect 12516 7980 12526 8036
rect 14130 7980 14140 8036
rect 14196 7980 16828 8036
rect 16884 7980 20412 8036
rect 20468 7980 21532 8036
rect 21588 7980 21598 8036
rect 8006 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8290 7868
rect 14810 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15094 7868
rect 21614 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21898 7868
rect 28418 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28702 7868
rect 24546 7644 24556 7700
rect 24612 7644 25340 7700
rect 25396 7644 26348 7700
rect 26404 7644 26414 7700
rect 5954 7532 5964 7588
rect 6020 7532 7196 7588
rect 7252 7532 7262 7588
rect 16258 7532 16268 7588
rect 16324 7532 17276 7588
rect 17332 7532 17342 7588
rect 29200 7392 30000 7504
rect 13234 7308 13244 7364
rect 13300 7308 15148 7364
rect 15204 7308 15214 7364
rect 24210 7308 24220 7364
rect 24276 7308 26236 7364
rect 26292 7308 26302 7364
rect 4604 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4888 7084
rect 11408 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11692 7084
rect 18212 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18496 7084
rect 25016 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25300 7084
rect 8652 6748 12684 6804
rect 12740 6748 12750 6804
rect 8652 6692 8708 6748
rect 29200 6720 30000 6832
rect 6514 6636 6524 6692
rect 6580 6636 7980 6692
rect 8036 6636 8652 6692
rect 8708 6636 8718 6692
rect 20514 6636 20524 6692
rect 20580 6636 21532 6692
rect 21588 6636 21598 6692
rect 24322 6636 24332 6692
rect 24388 6636 24668 6692
rect 24724 6636 27692 6692
rect 27748 6636 27758 6692
rect 18834 6524 18844 6580
rect 18900 6524 21980 6580
rect 22036 6524 22046 6580
rect 19618 6412 19628 6468
rect 19684 6412 22316 6468
rect 22372 6412 22382 6468
rect 8006 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8290 6300
rect 14810 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15094 6300
rect 21614 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21898 6300
rect 28418 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28702 6300
rect 29200 6132 30000 6160
rect 23090 6076 23100 6132
rect 23156 6076 30000 6132
rect 29200 6048 30000 6076
rect 19394 5964 19404 6020
rect 19460 5964 20860 6020
rect 20916 5964 20926 6020
rect 21074 5964 21084 6020
rect 21140 5964 22540 6020
rect 22596 5964 22606 6020
rect 12562 5852 12572 5908
rect 12628 5852 13468 5908
rect 13524 5852 13534 5908
rect 21074 5628 21084 5684
rect 21140 5628 26908 5684
rect 4604 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4888 5516
rect 11408 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11692 5516
rect 18212 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18496 5516
rect 25016 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25300 5516
rect 26852 5460 26908 5628
rect 29200 5460 30000 5488
rect 26852 5404 30000 5460
rect 29200 5376 30000 5404
rect 23314 5180 23324 5236
rect 23380 5180 25228 5236
rect 25284 5180 25294 5236
rect 21298 5068 21308 5124
rect 21364 5068 24556 5124
rect 24612 5068 25340 5124
rect 25396 5068 25406 5124
rect 22306 4956 22316 5012
rect 22372 4956 24780 5012
rect 24836 4956 24846 5012
rect 24434 4844 24444 4900
rect 24500 4844 26236 4900
rect 26292 4844 26302 4900
rect 28466 4844 28476 4900
rect 28532 4844 28868 4900
rect 28812 4788 28868 4844
rect 29200 4788 30000 4816
rect 28812 4732 30000 4788
rect 8006 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8290 4732
rect 14810 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15094 4732
rect 21614 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21898 4732
rect 28418 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28702 4732
rect 29200 4704 30000 4732
rect 21074 4508 21084 4564
rect 21140 4508 26124 4564
rect 26180 4508 26190 4564
rect 19282 4396 19292 4452
rect 19348 4396 22652 4452
rect 22708 4396 22718 4452
rect 24882 4396 24892 4452
rect 24948 4396 27244 4452
rect 27300 4396 27310 4452
rect 14690 4284 14700 4340
rect 14756 4284 16940 4340
rect 16996 4284 17006 4340
rect 21186 4284 21196 4340
rect 21252 4284 21644 4340
rect 21700 4284 21710 4340
rect 20402 4172 20412 4228
rect 20468 4172 26908 4228
rect 26852 4116 26908 4172
rect 29200 4116 30000 4144
rect 26852 4060 30000 4116
rect 29200 4032 30000 4060
rect 4604 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4888 3948
rect 11408 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11692 3948
rect 18212 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18496 3948
rect 25016 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25300 3948
rect 19506 3612 19516 3668
rect 19572 3612 23100 3668
rect 23156 3612 23166 3668
rect 16482 3500 16492 3556
rect 16548 3500 17164 3556
rect 17220 3500 17230 3556
rect 20178 3500 20188 3556
rect 20244 3500 22316 3556
rect 22372 3500 22382 3556
rect 29200 3444 30000 3472
rect 20290 3388 20300 3444
rect 20356 3388 21084 3444
rect 21140 3388 21150 3444
rect 28130 3388 28140 3444
rect 28196 3388 30000 3444
rect 29200 3360 30000 3388
rect 8006 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8290 3164
rect 14810 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15094 3164
rect 21614 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21898 3164
rect 28418 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28702 3164
rect 29200 2772 30000 2800
rect 18498 2716 18508 2772
rect 18564 2716 30000 2772
rect 29200 2688 30000 2716
rect 29200 2016 30000 2128
rect 29200 1344 30000 1456
rect 29200 672 30000 784
rect 29200 0 30000 112
<< via3 >>
rect 8016 26628 8072 26684
rect 8120 26628 8176 26684
rect 8224 26628 8280 26684
rect 14820 26628 14876 26684
rect 14924 26628 14980 26684
rect 15028 26628 15084 26684
rect 21624 26628 21680 26684
rect 21728 26628 21784 26684
rect 21832 26628 21888 26684
rect 28428 26628 28484 26684
rect 28532 26628 28588 26684
rect 28636 26628 28692 26684
rect 4614 25844 4670 25900
rect 4718 25844 4774 25900
rect 4822 25844 4878 25900
rect 11418 25844 11474 25900
rect 11522 25844 11578 25900
rect 11626 25844 11682 25900
rect 18222 25844 18278 25900
rect 18326 25844 18382 25900
rect 18430 25844 18486 25900
rect 25026 25844 25082 25900
rect 25130 25844 25186 25900
rect 25234 25844 25290 25900
rect 8016 25060 8072 25116
rect 8120 25060 8176 25116
rect 8224 25060 8280 25116
rect 14820 25060 14876 25116
rect 14924 25060 14980 25116
rect 15028 25060 15084 25116
rect 21624 25060 21680 25116
rect 21728 25060 21784 25116
rect 21832 25060 21888 25116
rect 28428 25060 28484 25116
rect 28532 25060 28588 25116
rect 28636 25060 28692 25116
rect 4614 24276 4670 24332
rect 4718 24276 4774 24332
rect 4822 24276 4878 24332
rect 11418 24276 11474 24332
rect 11522 24276 11578 24332
rect 11626 24276 11682 24332
rect 18222 24276 18278 24332
rect 18326 24276 18382 24332
rect 18430 24276 18486 24332
rect 25026 24276 25082 24332
rect 25130 24276 25186 24332
rect 25234 24276 25290 24332
rect 8016 23492 8072 23548
rect 8120 23492 8176 23548
rect 8224 23492 8280 23548
rect 14820 23492 14876 23548
rect 14924 23492 14980 23548
rect 15028 23492 15084 23548
rect 21624 23492 21680 23548
rect 21728 23492 21784 23548
rect 21832 23492 21888 23548
rect 28428 23492 28484 23548
rect 28532 23492 28588 23548
rect 28636 23492 28692 23548
rect 4614 22708 4670 22764
rect 4718 22708 4774 22764
rect 4822 22708 4878 22764
rect 11418 22708 11474 22764
rect 11522 22708 11578 22764
rect 11626 22708 11682 22764
rect 18222 22708 18278 22764
rect 18326 22708 18382 22764
rect 18430 22708 18486 22764
rect 25026 22708 25082 22764
rect 25130 22708 25186 22764
rect 25234 22708 25290 22764
rect 8016 21924 8072 21980
rect 8120 21924 8176 21980
rect 8224 21924 8280 21980
rect 14820 21924 14876 21980
rect 14924 21924 14980 21980
rect 15028 21924 15084 21980
rect 21624 21924 21680 21980
rect 21728 21924 21784 21980
rect 21832 21924 21888 21980
rect 28428 21924 28484 21980
rect 28532 21924 28588 21980
rect 28636 21924 28692 21980
rect 4614 21140 4670 21196
rect 4718 21140 4774 21196
rect 4822 21140 4878 21196
rect 11418 21140 11474 21196
rect 11522 21140 11578 21196
rect 11626 21140 11682 21196
rect 18222 21140 18278 21196
rect 18326 21140 18382 21196
rect 18430 21140 18486 21196
rect 25026 21140 25082 21196
rect 25130 21140 25186 21196
rect 25234 21140 25290 21196
rect 8016 20356 8072 20412
rect 8120 20356 8176 20412
rect 8224 20356 8280 20412
rect 14820 20356 14876 20412
rect 14924 20356 14980 20412
rect 15028 20356 15084 20412
rect 21624 20356 21680 20412
rect 21728 20356 21784 20412
rect 21832 20356 21888 20412
rect 28428 20356 28484 20412
rect 28532 20356 28588 20412
rect 28636 20356 28692 20412
rect 4614 19572 4670 19628
rect 4718 19572 4774 19628
rect 4822 19572 4878 19628
rect 11418 19572 11474 19628
rect 11522 19572 11578 19628
rect 11626 19572 11682 19628
rect 18222 19572 18278 19628
rect 18326 19572 18382 19628
rect 18430 19572 18486 19628
rect 25026 19572 25082 19628
rect 25130 19572 25186 19628
rect 25234 19572 25290 19628
rect 8016 18788 8072 18844
rect 8120 18788 8176 18844
rect 8224 18788 8280 18844
rect 14820 18788 14876 18844
rect 14924 18788 14980 18844
rect 15028 18788 15084 18844
rect 21624 18788 21680 18844
rect 21728 18788 21784 18844
rect 21832 18788 21888 18844
rect 28428 18788 28484 18844
rect 28532 18788 28588 18844
rect 28636 18788 28692 18844
rect 4614 18004 4670 18060
rect 4718 18004 4774 18060
rect 4822 18004 4878 18060
rect 11418 18004 11474 18060
rect 11522 18004 11578 18060
rect 11626 18004 11682 18060
rect 18222 18004 18278 18060
rect 18326 18004 18382 18060
rect 18430 18004 18486 18060
rect 25026 18004 25082 18060
rect 25130 18004 25186 18060
rect 25234 18004 25290 18060
rect 8016 17220 8072 17276
rect 8120 17220 8176 17276
rect 8224 17220 8280 17276
rect 14820 17220 14876 17276
rect 14924 17220 14980 17276
rect 15028 17220 15084 17276
rect 21624 17220 21680 17276
rect 21728 17220 21784 17276
rect 21832 17220 21888 17276
rect 28428 17220 28484 17276
rect 28532 17220 28588 17276
rect 28636 17220 28692 17276
rect 4614 16436 4670 16492
rect 4718 16436 4774 16492
rect 4822 16436 4878 16492
rect 11418 16436 11474 16492
rect 11522 16436 11578 16492
rect 11626 16436 11682 16492
rect 18222 16436 18278 16492
rect 18326 16436 18382 16492
rect 18430 16436 18486 16492
rect 25026 16436 25082 16492
rect 25130 16436 25186 16492
rect 25234 16436 25290 16492
rect 8016 15652 8072 15708
rect 8120 15652 8176 15708
rect 8224 15652 8280 15708
rect 14820 15652 14876 15708
rect 14924 15652 14980 15708
rect 15028 15652 15084 15708
rect 21624 15652 21680 15708
rect 21728 15652 21784 15708
rect 21832 15652 21888 15708
rect 28428 15652 28484 15708
rect 28532 15652 28588 15708
rect 28636 15652 28692 15708
rect 4614 14868 4670 14924
rect 4718 14868 4774 14924
rect 4822 14868 4878 14924
rect 11418 14868 11474 14924
rect 11522 14868 11578 14924
rect 11626 14868 11682 14924
rect 18222 14868 18278 14924
rect 18326 14868 18382 14924
rect 18430 14868 18486 14924
rect 25026 14868 25082 14924
rect 25130 14868 25186 14924
rect 25234 14868 25290 14924
rect 8016 14084 8072 14140
rect 8120 14084 8176 14140
rect 8224 14084 8280 14140
rect 14820 14084 14876 14140
rect 14924 14084 14980 14140
rect 15028 14084 15084 14140
rect 21624 14084 21680 14140
rect 21728 14084 21784 14140
rect 21832 14084 21888 14140
rect 28428 14084 28484 14140
rect 28532 14084 28588 14140
rect 28636 14084 28692 14140
rect 4614 13300 4670 13356
rect 4718 13300 4774 13356
rect 4822 13300 4878 13356
rect 11418 13300 11474 13356
rect 11522 13300 11578 13356
rect 11626 13300 11682 13356
rect 18222 13300 18278 13356
rect 18326 13300 18382 13356
rect 18430 13300 18486 13356
rect 25026 13300 25082 13356
rect 25130 13300 25186 13356
rect 25234 13300 25290 13356
rect 8016 12516 8072 12572
rect 8120 12516 8176 12572
rect 8224 12516 8280 12572
rect 14820 12516 14876 12572
rect 14924 12516 14980 12572
rect 15028 12516 15084 12572
rect 21624 12516 21680 12572
rect 21728 12516 21784 12572
rect 21832 12516 21888 12572
rect 28428 12516 28484 12572
rect 28532 12516 28588 12572
rect 28636 12516 28692 12572
rect 8428 12012 8484 12068
rect 4614 11732 4670 11788
rect 4718 11732 4774 11788
rect 4822 11732 4878 11788
rect 11418 11732 11474 11788
rect 11522 11732 11578 11788
rect 11626 11732 11682 11788
rect 18222 11732 18278 11788
rect 18326 11732 18382 11788
rect 18430 11732 18486 11788
rect 25026 11732 25082 11788
rect 25130 11732 25186 11788
rect 25234 11732 25290 11788
rect 8428 11676 8484 11732
rect 8016 10948 8072 11004
rect 8120 10948 8176 11004
rect 8224 10948 8280 11004
rect 14820 10948 14876 11004
rect 14924 10948 14980 11004
rect 15028 10948 15084 11004
rect 21624 10948 21680 11004
rect 21728 10948 21784 11004
rect 21832 10948 21888 11004
rect 28428 10948 28484 11004
rect 28532 10948 28588 11004
rect 28636 10948 28692 11004
rect 4614 10164 4670 10220
rect 4718 10164 4774 10220
rect 4822 10164 4878 10220
rect 11418 10164 11474 10220
rect 11522 10164 11578 10220
rect 11626 10164 11682 10220
rect 18222 10164 18278 10220
rect 18326 10164 18382 10220
rect 18430 10164 18486 10220
rect 25026 10164 25082 10220
rect 25130 10164 25186 10220
rect 25234 10164 25290 10220
rect 8016 9380 8072 9436
rect 8120 9380 8176 9436
rect 8224 9380 8280 9436
rect 14820 9380 14876 9436
rect 14924 9380 14980 9436
rect 15028 9380 15084 9436
rect 21624 9380 21680 9436
rect 21728 9380 21784 9436
rect 21832 9380 21888 9436
rect 28428 9380 28484 9436
rect 28532 9380 28588 9436
rect 28636 9380 28692 9436
rect 4614 8596 4670 8652
rect 4718 8596 4774 8652
rect 4822 8596 4878 8652
rect 11418 8596 11474 8652
rect 11522 8596 11578 8652
rect 11626 8596 11682 8652
rect 18222 8596 18278 8652
rect 18326 8596 18382 8652
rect 18430 8596 18486 8652
rect 25026 8596 25082 8652
rect 25130 8596 25186 8652
rect 25234 8596 25290 8652
rect 8016 7812 8072 7868
rect 8120 7812 8176 7868
rect 8224 7812 8280 7868
rect 14820 7812 14876 7868
rect 14924 7812 14980 7868
rect 15028 7812 15084 7868
rect 21624 7812 21680 7868
rect 21728 7812 21784 7868
rect 21832 7812 21888 7868
rect 28428 7812 28484 7868
rect 28532 7812 28588 7868
rect 28636 7812 28692 7868
rect 4614 7028 4670 7084
rect 4718 7028 4774 7084
rect 4822 7028 4878 7084
rect 11418 7028 11474 7084
rect 11522 7028 11578 7084
rect 11626 7028 11682 7084
rect 18222 7028 18278 7084
rect 18326 7028 18382 7084
rect 18430 7028 18486 7084
rect 25026 7028 25082 7084
rect 25130 7028 25186 7084
rect 25234 7028 25290 7084
rect 8016 6244 8072 6300
rect 8120 6244 8176 6300
rect 8224 6244 8280 6300
rect 14820 6244 14876 6300
rect 14924 6244 14980 6300
rect 15028 6244 15084 6300
rect 21624 6244 21680 6300
rect 21728 6244 21784 6300
rect 21832 6244 21888 6300
rect 28428 6244 28484 6300
rect 28532 6244 28588 6300
rect 28636 6244 28692 6300
rect 4614 5460 4670 5516
rect 4718 5460 4774 5516
rect 4822 5460 4878 5516
rect 11418 5460 11474 5516
rect 11522 5460 11578 5516
rect 11626 5460 11682 5516
rect 18222 5460 18278 5516
rect 18326 5460 18382 5516
rect 18430 5460 18486 5516
rect 25026 5460 25082 5516
rect 25130 5460 25186 5516
rect 25234 5460 25290 5516
rect 8016 4676 8072 4732
rect 8120 4676 8176 4732
rect 8224 4676 8280 4732
rect 14820 4676 14876 4732
rect 14924 4676 14980 4732
rect 15028 4676 15084 4732
rect 21624 4676 21680 4732
rect 21728 4676 21784 4732
rect 21832 4676 21888 4732
rect 28428 4676 28484 4732
rect 28532 4676 28588 4732
rect 28636 4676 28692 4732
rect 4614 3892 4670 3948
rect 4718 3892 4774 3948
rect 4822 3892 4878 3948
rect 11418 3892 11474 3948
rect 11522 3892 11578 3948
rect 11626 3892 11682 3948
rect 18222 3892 18278 3948
rect 18326 3892 18382 3948
rect 18430 3892 18486 3948
rect 25026 3892 25082 3948
rect 25130 3892 25186 3948
rect 25234 3892 25290 3948
rect 8016 3108 8072 3164
rect 8120 3108 8176 3164
rect 8224 3108 8280 3164
rect 14820 3108 14876 3164
rect 14924 3108 14980 3164
rect 15028 3108 15084 3164
rect 21624 3108 21680 3164
rect 21728 3108 21784 3164
rect 21832 3108 21888 3164
rect 28428 3108 28484 3164
rect 28532 3108 28588 3164
rect 28636 3108 28692 3164
<< metal4 >>
rect 4586 25900 4906 26716
rect 4586 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4906 25900
rect 4586 24332 4906 25844
rect 4586 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4906 24332
rect 4586 22764 4906 24276
rect 4586 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4906 22764
rect 4586 21196 4906 22708
rect 4586 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4906 21196
rect 4586 19628 4906 21140
rect 4586 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4906 19628
rect 4586 18060 4906 19572
rect 4586 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4906 18060
rect 4586 16492 4906 18004
rect 4586 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4906 16492
rect 4586 14924 4906 16436
rect 4586 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4906 14924
rect 4586 13356 4906 14868
rect 4586 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4906 13356
rect 4586 11788 4906 13300
rect 4586 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4906 11788
rect 4586 10220 4906 11732
rect 4586 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4906 10220
rect 4586 8652 4906 10164
rect 4586 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4906 8652
rect 4586 7084 4906 8596
rect 4586 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4906 7084
rect 4586 5516 4906 7028
rect 4586 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4906 5516
rect 4586 3948 4906 5460
rect 4586 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4906 3948
rect 4586 3076 4906 3892
rect 7988 26684 8308 26716
rect 7988 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8308 26684
rect 7988 25116 8308 26628
rect 7988 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8308 25116
rect 7988 23548 8308 25060
rect 7988 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8308 23548
rect 7988 21980 8308 23492
rect 7988 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8308 21980
rect 7988 20412 8308 21924
rect 7988 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8308 20412
rect 7988 18844 8308 20356
rect 7988 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8308 18844
rect 7988 17276 8308 18788
rect 7988 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8308 17276
rect 7988 15708 8308 17220
rect 7988 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8308 15708
rect 7988 14140 8308 15652
rect 7988 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8308 14140
rect 7988 12572 8308 14084
rect 7988 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8308 12572
rect 7988 11004 8308 12516
rect 11390 25900 11710 26716
rect 11390 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11710 25900
rect 11390 24332 11710 25844
rect 11390 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11710 24332
rect 11390 22764 11710 24276
rect 11390 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11710 22764
rect 11390 21196 11710 22708
rect 11390 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11710 21196
rect 11390 19628 11710 21140
rect 11390 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11710 19628
rect 11390 18060 11710 19572
rect 11390 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11710 18060
rect 11390 16492 11710 18004
rect 11390 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11710 16492
rect 11390 14924 11710 16436
rect 11390 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11710 14924
rect 11390 13356 11710 14868
rect 11390 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11710 13356
rect 8428 12068 8484 12078
rect 8428 11732 8484 12012
rect 8428 11666 8484 11676
rect 11390 11788 11710 13300
rect 11390 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11710 11788
rect 7988 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8308 11004
rect 7988 9436 8308 10948
rect 7988 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8308 9436
rect 7988 7868 8308 9380
rect 7988 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8308 7868
rect 7988 6300 8308 7812
rect 7988 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8308 6300
rect 7988 4732 8308 6244
rect 7988 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8308 4732
rect 7988 3164 8308 4676
rect 7988 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8308 3164
rect 7988 3076 8308 3108
rect 11390 10220 11710 11732
rect 11390 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11710 10220
rect 11390 8652 11710 10164
rect 11390 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11710 8652
rect 11390 7084 11710 8596
rect 11390 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11710 7084
rect 11390 5516 11710 7028
rect 11390 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11710 5516
rect 11390 3948 11710 5460
rect 11390 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11710 3948
rect 11390 3076 11710 3892
rect 14792 26684 15112 26716
rect 14792 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15112 26684
rect 14792 25116 15112 26628
rect 14792 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15112 25116
rect 14792 23548 15112 25060
rect 14792 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15112 23548
rect 14792 21980 15112 23492
rect 14792 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15112 21980
rect 14792 20412 15112 21924
rect 14792 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15112 20412
rect 14792 18844 15112 20356
rect 14792 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15112 18844
rect 14792 17276 15112 18788
rect 14792 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15112 17276
rect 14792 15708 15112 17220
rect 14792 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15112 15708
rect 14792 14140 15112 15652
rect 14792 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15112 14140
rect 14792 12572 15112 14084
rect 14792 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15112 12572
rect 14792 11004 15112 12516
rect 14792 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15112 11004
rect 14792 9436 15112 10948
rect 14792 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15112 9436
rect 14792 7868 15112 9380
rect 14792 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15112 7868
rect 14792 6300 15112 7812
rect 14792 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15112 6300
rect 14792 4732 15112 6244
rect 14792 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15112 4732
rect 14792 3164 15112 4676
rect 14792 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15112 3164
rect 14792 3076 15112 3108
rect 18194 25900 18514 26716
rect 18194 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18514 25900
rect 18194 24332 18514 25844
rect 18194 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18514 24332
rect 18194 22764 18514 24276
rect 18194 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18514 22764
rect 18194 21196 18514 22708
rect 18194 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18514 21196
rect 18194 19628 18514 21140
rect 18194 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18514 19628
rect 18194 18060 18514 19572
rect 18194 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18514 18060
rect 18194 16492 18514 18004
rect 18194 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18514 16492
rect 18194 14924 18514 16436
rect 18194 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18514 14924
rect 18194 13356 18514 14868
rect 18194 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18514 13356
rect 18194 11788 18514 13300
rect 18194 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18514 11788
rect 18194 10220 18514 11732
rect 18194 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18514 10220
rect 18194 8652 18514 10164
rect 18194 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18514 8652
rect 18194 7084 18514 8596
rect 18194 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18514 7084
rect 18194 5516 18514 7028
rect 18194 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18514 5516
rect 18194 3948 18514 5460
rect 18194 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18514 3948
rect 18194 3076 18514 3892
rect 21596 26684 21916 26716
rect 21596 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21916 26684
rect 21596 25116 21916 26628
rect 21596 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21916 25116
rect 21596 23548 21916 25060
rect 21596 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21916 23548
rect 21596 21980 21916 23492
rect 21596 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21916 21980
rect 21596 20412 21916 21924
rect 21596 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21916 20412
rect 21596 18844 21916 20356
rect 21596 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21916 18844
rect 21596 17276 21916 18788
rect 21596 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21916 17276
rect 21596 15708 21916 17220
rect 21596 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21916 15708
rect 21596 14140 21916 15652
rect 21596 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21916 14140
rect 21596 12572 21916 14084
rect 21596 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21916 12572
rect 21596 11004 21916 12516
rect 21596 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21916 11004
rect 21596 9436 21916 10948
rect 21596 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21916 9436
rect 21596 7868 21916 9380
rect 21596 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21916 7868
rect 21596 6300 21916 7812
rect 21596 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21916 6300
rect 21596 4732 21916 6244
rect 21596 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21916 4732
rect 21596 3164 21916 4676
rect 21596 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21916 3164
rect 21596 3076 21916 3108
rect 24998 25900 25318 26716
rect 24998 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25318 25900
rect 24998 24332 25318 25844
rect 24998 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25318 24332
rect 24998 22764 25318 24276
rect 24998 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25318 22764
rect 24998 21196 25318 22708
rect 24998 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25318 21196
rect 24998 19628 25318 21140
rect 24998 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25318 19628
rect 24998 18060 25318 19572
rect 24998 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25318 18060
rect 24998 16492 25318 18004
rect 24998 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25318 16492
rect 24998 14924 25318 16436
rect 24998 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25318 14924
rect 24998 13356 25318 14868
rect 24998 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25318 13356
rect 24998 11788 25318 13300
rect 24998 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25318 11788
rect 24998 10220 25318 11732
rect 24998 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25318 10220
rect 24998 8652 25318 10164
rect 24998 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25318 8652
rect 24998 7084 25318 8596
rect 24998 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25318 7084
rect 24998 5516 25318 7028
rect 24998 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25318 5516
rect 24998 3948 25318 5460
rect 24998 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25318 3948
rect 24998 3076 25318 3892
rect 28400 26684 28720 26716
rect 28400 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28720 26684
rect 28400 25116 28720 26628
rect 28400 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28720 25116
rect 28400 23548 28720 25060
rect 28400 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28720 23548
rect 28400 21980 28720 23492
rect 28400 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28720 21980
rect 28400 20412 28720 21924
rect 28400 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28720 20412
rect 28400 18844 28720 20356
rect 28400 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28720 18844
rect 28400 17276 28720 18788
rect 28400 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28720 17276
rect 28400 15708 28720 17220
rect 28400 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28720 15708
rect 28400 14140 28720 15652
rect 28400 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28720 14140
rect 28400 12572 28720 14084
rect 28400 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28720 12572
rect 28400 11004 28720 12516
rect 28400 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28720 11004
rect 28400 9436 28720 10948
rect 28400 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28720 9436
rect 28400 7868 28720 9380
rect 28400 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28720 7868
rect 28400 6300 28720 7812
rect 28400 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28720 6300
rect 28400 4732 28720 6244
rect 28400 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28720 4732
rect 28400 3164 28720 4676
rect 28400 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28720 3164
rect 28400 3076 28720 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _053_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _054_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _055_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _056_
timestamp 1698431365
transform 1 0 3472 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _057_
timestamp 1698431365
transform -1 0 6272 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _058_
timestamp 1698431365
transform -1 0 4816 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _059_
timestamp 1698431365
transform -1 0 11648 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _060_
timestamp 1698431365
transform 1 0 7728 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _061_
timestamp 1698431365
transform -1 0 16912 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _062_
timestamp 1698431365
transform -1 0 12432 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _063_
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _064_
timestamp 1698431365
transform -1 0 12992 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _065_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _066_
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _067_
timestamp 1698431365
transform -1 0 19936 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _068_
timestamp 1698431365
transform -1 0 24864 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _069_
timestamp 1698431365
transform -1 0 24752 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _070_
timestamp 1698431365
transform 1 0 27552 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _071_
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _072_
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _073_
timestamp 1698431365
transform -1 0 27440 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _074_
timestamp 1698431365
transform 1 0 19936 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _075_
timestamp 1698431365
transform -1 0 19936 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _076_
timestamp 1698431365
transform -1 0 14896 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _077_
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _078_
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _079_
timestamp 1698431365
transform -1 0 6608 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _080_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _081_
timestamp 1698431365
transform -1 0 5264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _082_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _083_
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _084_
timestamp 1698431365
transform -1 0 6160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _085_
timestamp 1698431365
transform -1 0 12544 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _086_
timestamp 1698431365
transform -1 0 10080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _087_
timestamp 1698431365
transform 1 0 14224 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _088_
timestamp 1698431365
transform 1 0 15792 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _089_
timestamp 1698431365
transform -1 0 14112 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _090_
timestamp 1698431365
transform 1 0 19376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _091_
timestamp 1698431365
transform 1 0 17472 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _092_
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _093_
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _094_
timestamp 1698431365
transform -1 0 28112 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _095_
timestamp 1698431365
transform -1 0 27440 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _096_
timestamp 1698431365
transform -1 0 24752 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _097_
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _098_
timestamp 1698431365
transform 1 0 12432 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _099_
timestamp 1698431365
transform -1 0 28336 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _100_
timestamp 1698431365
transform -1 0 19264 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _101_
timestamp 1698431365
transform -1 0 20608 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _102_
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _103_
timestamp 1698431365
transform -1 0 22176 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _104_
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _105_
timestamp 1698431365
transform -1 0 27216 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4144 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _107_
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _108_
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _109_
timestamp 1698431365
transform -1 0 5376 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _110_
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _111_
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _112_
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _113_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _114_
timestamp 1698431365
transform 1 0 12656 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _115_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _116_
timestamp 1698431365
transform 1 0 17472 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _117_
timestamp 1698431365
transform 1 0 15456 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _118_
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _119_
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _120_
timestamp 1698431365
transform 1 0 24528 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _121_
timestamp 1698431365
transform 1 0 21056 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _122_
timestamp 1698431365
transform 1 0 23744 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _123_
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _124_
timestamp 1698431365
transform -1 0 21056 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _125_
timestamp 1698431365
transform 1 0 15456 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _126_
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _127_
timestamp 1698431365
transform -1 0 10976 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _128_
timestamp 1698431365
transform -1 0 7952 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _129_
timestamp 1698431365
transform -1 0 14896 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _130_
timestamp 1698431365
transform -1 0 5824 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _131_
timestamp 1698431365
transform -1 0 10416 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _132_
timestamp 1698431365
transform 1 0 4592 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _133_
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _134_
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _135_
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _136_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _137_
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _138_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _139_
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _140_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _141_
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _142_
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _143_
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _144_
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _145_
timestamp 1698431365
transform 1 0 24528 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _146_
timestamp 1698431365
transform 1 0 10416 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _147_
timestamp 1698431365
transform -1 0 26992 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _148_
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _149_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _150_
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _151_
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _152_
timestamp 1698431365
transform 1 0 24528 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _153_
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1698431365
transform 1 0 18592 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _180_
timestamp 1698431365
transform 1 0 19152 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _183_
timestamp 1698431365
transform -1 0 27664 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1698431365
transform 1 0 19824 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _185_
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _187_
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _188_
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _189_
timestamp 1698431365
transform -1 0 27552 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _190_
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _191_
timestamp 1698431365
transform 1 0 14448 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _192_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _193_
timestamp 1698431365
transform -1 0 22176 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1698431365
transform -1 0 3472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1698431365
transform 1 0 11648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1698431365
transform 1 0 8624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I
timestamp 1698431365
transform 1 0 14784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1698431365
transform 1 0 13216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1698431365
transform 1 0 21504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1698431365
transform 1 0 14336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1698431365
transform 1 0 24192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I
timestamp 1698431365
transform 1 0 28112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I
timestamp 1698431365
transform 1 0 25872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1698431365
transform -1 0 12432 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1698431365
transform 1 0 28000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I
timestamp 1698431365
transform 1 0 25872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__I
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__CLK
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__CLK
timestamp 1698431365
transform 1 0 19712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__CLK
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__CLK
timestamp 1698431365
transform 1 0 25872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__CLK
timestamp 1698431365
transform 1 0 26320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__CLK
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__CLK
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__CLK
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__CLK
timestamp 1698431365
transform 1 0 21280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__CLK
timestamp 1698431365
transform 1 0 17808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__CLK
timestamp 1698431365
transform 1 0 25200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__CLK
timestamp 1698431365
transform 1 0 22736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__CLK
timestamp 1698431365
transform -1 0 26096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__CLK
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__CLK
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__CLK
timestamp 1698431365
transform -1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__CLK
timestamp 1698431365
transform 1 0 21728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__CLK
timestamp 1698431365
transform 1 0 25872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform -1 0 15008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 22512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 27216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 10864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 12096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 18816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 19600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 12768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 22288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 26992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 19712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1698431365
transform -1 0 15008 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_118 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_132
timestamp 1698431365
transform 1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_148
timestamp 1698431365
transform 1 0 17920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_150 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_163
timestamp 1698431365
transform 1 0 19600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_199
timestamp 1698431365
transform 1 0 23632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_211
timestamp 1698431365
transform 1 0 24976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_219
timestamp 1698431365
transform 1 0 25872 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_88
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_96
timestamp 1698431365
transform 1 0 12096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_100
timestamp 1698431365
transform 1 0 12544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_104
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_112
timestamp 1698431365
transform 1 0 13888 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_127
timestamp 1698431365
transform 1 0 15568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_135
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1698431365
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_152
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_162
timestamp 1698431365
transform 1 0 19488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_198
timestamp 1698431365
transform 1 0 23520 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_206
timestamp 1698431365
transform 1 0 24416 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_104
timestamp 1698431365
transform 1 0 12992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_106
timestamp 1698431365
transform 1 0 13216 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_113
timestamp 1698431365
transform 1 0 14000 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_117
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_119
timestamp 1698431365
transform 1 0 14672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_128
timestamp 1698431365
transform 1 0 15680 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_158
timestamp 1698431365
transform 1 0 19040 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_166
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_170
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_63
timestamp 1698431365
transform 1 0 8400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_67
timestamp 1698431365
transform 1 0 8848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_132
timestamp 1698431365
transform 1 0 16128 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_164
timestamp 1698431365
transform 1 0 19712 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_196
timestamp 1698431365
transform 1 0 23296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_36
timestamp 1698431365
transform 1 0 5376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_40
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_89
timestamp 1698431365
transform 1 0 11312 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_97
timestamp 1698431365
transform 1 0 12208 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_104
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_108
timestamp 1698431365
transform 1 0 13440 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_116
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_174
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_6
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_24
timestamp 1698431365
transform 1 0 4032 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_44
timestamp 1698431365
transform 1 0 6272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_48
timestamp 1698431365
transform 1 0 6720 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_52
timestamp 1698431365
transform 1 0 7168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_135
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_143
timestamp 1698431365
transform 1 0 17360 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_160
timestamp 1698431365
transform 1 0 19264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_202
timestamp 1698431365
transform 1 0 23968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_206
timestamp 1698431365
transform 1 0 24416 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_6
timestamp 1698431365
transform 1 0 2016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_42
timestamp 1698431365
transform 1 0 6048 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_50
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_92
timestamp 1698431365
transform 1 0 11648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_100
timestamp 1698431365
transform 1 0 12544 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_135
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_178
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_182
timestamp 1698431365
transform 1 0 21728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_186
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_237
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_22
timestamp 1698431365
transform 1 0 3808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_24
timestamp 1698431365
transform 1 0 4032 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_125
timestamp 1698431365
transform 1 0 15344 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_166
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_203
timestamp 1698431365
transform 1 0 24080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_90
timestamp 1698431365
transform 1 0 11424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_94
timestamp 1698431365
transform 1 0 11872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_98
timestamp 1698431365
transform 1 0 12320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_154
timestamp 1698431365
transform 1 0 18592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_162
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_200
timestamp 1698431365
transform 1 0 23744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_237
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_49
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_51
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_99
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_125
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_16
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_63
timestamp 1698431365
transform 1 0 8400 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_237
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_44
timestamp 1698431365
transform 1 0 6272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_48
timestamp 1698431365
transform 1 0 6720 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_52
timestamp 1698431365
transform 1 0 7168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_103
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_119
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_237
timestamp 1698431365
transform 1 0 27888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_22
timestamp 1698431365
transform 1 0 3808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_24
timestamp 1698431365
transform 1 0 4032 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_59
timestamp 1698431365
transform 1 0 7952 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_63
timestamp 1698431365
transform 1 0 8400 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_84
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_86
timestamp 1698431365
transform 1 0 10976 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_121
timestamp 1698431365
transform 1 0 14896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_125
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698431365
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_237
timestamp 1698431365
transform 1 0 27888 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_81
timestamp 1698431365
transform 1 0 10416 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_89
timestamp 1698431365
transform 1 0 11312 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_125
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_161
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_163
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_166
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_170
timestamp 1698431365
transform 1 0 20384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_179
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_186
timestamp 1698431365
transform 1 0 22176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_188
timestamp 1698431365
transform 1 0 22400 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_40
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_44
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_180
timestamp 1698431365
transform 1 0 21504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_184
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_186
timestamp 1698431365
transform 1 0 22176 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698431365
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_228
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_232
timestamp 1698431365
transform 1 0 27328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_236
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_240
timestamp 1698431365
transform 1 0 28224 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_18
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_43
timestamp 1698431365
transform 1 0 6160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_81
timestamp 1698431365
transform 1 0 10416 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_149
timestamp 1698431365
transform 1 0 18032 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_20
timestamp 1698431365
transform 1 0 3584 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_28
timestamp 1698431365
transform 1 0 4480 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_63
timestamp 1698431365
transform 1 0 8400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_67
timestamp 1698431365
transform 1 0 8848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_115
timestamp 1698431365
transform 1 0 14224 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_123
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_149
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_237
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_10
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_59
timestamp 1698431365
transform 1 0 7952 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_100
timestamp 1698431365
transform 1 0 12544 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_160
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_167
timestamp 1698431365
transform 1 0 20048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_202
timestamp 1698431365
transform 1 0 23968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_206
timestamp 1698431365
transform 1 0 24416 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_42
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_50
timestamp 1698431365
transform 1 0 6944 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_176
timestamp 1698431365
transform 1 0 21056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_180
timestamp 1698431365
transform 1 0 21504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_184
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_224
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_63
timestamp 1698431365
transform 1 0 8400 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_80
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_88
timestamp 1698431365
transform 1 0 11200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_141
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_149
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_166
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_211
timestamp 1698431365
transform 1 0 24976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_215
timestamp 1698431365
transform 1 0 25424 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_98
timestamp 1698431365
transform 1 0 12320 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_106
timestamp 1698431365
transform 1 0 13216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_114
timestamp 1698431365
transform 1 0 14112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_118
timestamp 1698431365
transform 1 0 14560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_122
timestamp 1698431365
transform 1 0 15008 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_189
timestamp 1698431365
transform 1 0 22512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_193
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_237
timestamp 1698431365
transform 1 0 27888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_141
timestamp 1698431365
transform 1 0 17136 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_144
timestamp 1698431365
transform 1 0 17472 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_160
timestamp 1698431365
transform 1 0 19264 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_120
timestamp 1698431365
transform 1 0 14784 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698431365
transform 1 0 25760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_237
timestamp 1698431365
transform 1 0 27888 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_209
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_225
timestamp 1698431365
transform 1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_224
timestamp 1698431365
transform 1 0 26432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_75
timestamp 1698431365
transform 1 0 9744 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_91
timestamp 1698431365
transform 1 0 11536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_99
timestamp 1698431365
transform 1 0 12432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_139
timestamp 1698431365
transform 1 0 16912 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_147
timestamp 1698431365
transform 1 0 17808 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_151
timestamp 1698431365
transform 1 0 18256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_153
timestamp 1698431365
transform 1 0 18480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_160
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_209
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_225
timestamp 1698431365
transform 1 0 26544 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698431365
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_96
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_100
timestamp 1698431365
transform 1 0 12544 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_107
timestamp 1698431365
transform 1 0 13328 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_178
timestamp 1698431365
transform 1 0 21280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_180
timestamp 1698431365
transform 1 0 21504 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_183
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_189
timestamp 1698431365
transform 1 0 22512 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_234
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_236
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_6
timestamp 1698431365
transform 1 0 2016 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_30
timestamp 1698431365
transform 1 0 4704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_81
timestamp 1698431365
transform 1 0 10416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_95
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_117
timestamp 1698431365
transform 1 0 14448 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_129
timestamp 1698431365
transform 1 0 15792 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_132
timestamp 1698431365
transform 1 0 16128 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_143
timestamp 1698431365
transform 1 0 17360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_195
timestamp 1698431365
transform 1 0 23184 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_227
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_54
timestamp 1698431365
transform 1 0 7392 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_70
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_89
timestamp 1698431365
transform 1 0 11312 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_93
timestamp 1698431365
transform 1 0 11760 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_104
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_119
timestamp 1698431365
transform 1 0 14672 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_123
timestamp 1698431365
transform 1 0 15120 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_149
timestamp 1698431365
transform 1 0 18032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_167
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_169
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_182
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_210
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_215
timestamp 1698431365
transform 1 0 25424 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_219
timestamp 1698431365
transform 1 0 25872 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_240
timestamp 1698431365
transform 1 0 28224 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27888 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 20048 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 19936 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 19264 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 19936 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform -1 0 27888 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 16912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 7840 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 27888 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform 1 0 21728 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 23856 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 27888 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 24304 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform 1 0 9520 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform -1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 24080 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 10304 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 5264 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 23968 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform -1 0 8848 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 6384 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 27888 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 23968 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 12320 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 23184 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 9184 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 28336 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 16576 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 27888 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 28336 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 9072 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform -1 0 28336 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform -1 0 16128 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform -1 0 27888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform -1 0 20272 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 27776 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 10192 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 23184 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 28336 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 10864 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 12096 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 18256 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 22512 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 17472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 15904 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 21392 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 20496 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 16576 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 28336 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 19600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output19 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28336 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output20
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output21
timestamp 1698431365
transform 1 0 22176 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output22
timestamp 1698431365
transform 1 0 20608 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output23
timestamp 1698431365
transform -1 0 14560 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output24
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output25
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output27
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output29
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output30
timestamp 1698431365
transform 1 0 13552 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output31
timestamp 1698431365
transform 1 0 10192 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output32
timestamp 1698431365
transform -1 0 21056 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output33
timestamp 1698431365
transform 1 0 22176 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output34
timestamp 1698431365
transform 1 0 15008 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output35
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_30 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 28560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_31
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_32
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_33
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_34
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_35
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_36
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_37
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_38
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_39
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_40
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_41
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 28560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_42
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_43
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_44
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_45
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_46
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_47
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_48
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_49
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_50
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 28560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 28560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27888 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__37
timestamp 1698431365
transform -1 0 18368 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__38
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__39
timestamp 1698431365
transform -1 0 14448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__40
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__41
timestamp 1698431365
transform -1 0 7952 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__42
timestamp 1698431365
transform -1 0 13440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__43
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__44
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__45
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__46
timestamp 1698431365
transform -1 0 25424 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__47
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__48
timestamp 1698431365
transform 1 0 21280 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__49
timestamp 1698431365
transform 1 0 24528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__50
timestamp 1698431365
transform -1 0 17920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__51
timestamp 1698431365
transform -1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__52
timestamp 1698431365
transform -1 0 24192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__53
timestamp 1698431365
transform -1 0 15568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__54
timestamp 1698431365
transform 1 0 27440 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__55
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__56
timestamp 1698431365
transform -1 0 15344 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__57
timestamp 1698431365
transform -1 0 2016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__58
timestamp 1698431365
transform -1 0 11984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__0__59
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_61
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_62
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_63
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_64
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_65
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_66
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_67
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_68
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_69
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_70
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_71
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_72
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_73
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_74
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_75
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_76
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_77
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_78
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_81
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_86
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_87
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_88
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_89
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_90
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_91
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_92
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_93
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_94
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_95
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_96
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_97
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_98
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_99
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_100
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_101
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_102
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_103
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_104
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_105
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_106
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_107
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_108
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_109
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_110
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_111
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_112
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_113
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_114
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_115
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_116
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_117
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_118
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_119
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_120
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_121
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_122
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_123
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_124
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_125
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_126
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_127
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_128
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_129
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_130
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_131
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_132
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_133
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_134
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_135
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_136
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_137
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_138
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_139
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_140
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_141
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_142
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_143
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_144
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_145
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_146
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_147
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_148
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_149
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_150
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_151
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_152
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_153
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_154
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_155
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_156
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_157
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 29200 14784 30000 14896 0 FreeSans 448 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 9408 29200 9520 30000 0 FreeSans 448 90 0 0 chanx_right_in[0]
port 2 nsew signal input
flabel metal2 s 22176 29200 22288 30000 0 FreeSans 448 90 0 0 chanx_right_in[10]
port 3 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 chanx_right_in[11]
port 4 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 chanx_right_in[12]
port 5 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 chanx_right_in[13]
port 6 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 chanx_right_in[14]
port 7 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 chanx_right_in[15]
port 8 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 chanx_right_in[16]
port 9 nsew signal input
flabel metal3 s 29200 26880 30000 26992 0 FreeSans 448 0 0 0 chanx_right_in[17]
port 10 nsew signal input
flabel metal2 s 10752 29200 10864 30000 0 FreeSans 448 90 0 0 chanx_right_in[18]
port 11 nsew signal input
flabel metal2 s 12096 29200 12208 30000 0 FreeSans 448 90 0 0 chanx_right_in[19]
port 12 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chanx_right_in[1]
port 13 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chanx_right_in[2]
port 14 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 chanx_right_in[3]
port 15 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 chanx_right_in[4]
port 16 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chanx_right_in[5]
port 17 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chanx_right_in[6]
port 18 nsew signal input
flabel metal3 s 29200 2688 30000 2800 0 FreeSans 448 0 0 0 chanx_right_in[7]
port 19 nsew signal input
flabel metal2 s 20832 29200 20944 30000 0 FreeSans 448 90 0 0 chanx_right_in[8]
port 20 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chanx_right_in[9]
port 21 nsew signal input
flabel metal3 s 29200 22848 30000 22960 0 FreeSans 448 0 0 0 chanx_right_out[0]
port 22 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chanx_right_out[10]
port 23 nsew signal tristate
flabel metal2 s 22848 29200 22960 30000 0 FreeSans 448 90 0 0 chanx_right_out[11]
port 24 nsew signal tristate
flabel metal2 s 8064 29200 8176 30000 0 FreeSans 448 90 0 0 chanx_right_out[12]
port 25 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chanx_right_out[13]
port 26 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 chanx_right_out[14]
port 27 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 chanx_right_out[15]
port 28 nsew signal tristate
flabel metal2 s 18144 29200 18256 30000 0 FreeSans 448 90 0 0 chanx_right_out[16]
port 29 nsew signal tristate
flabel metal3 s 29200 6048 30000 6160 0 FreeSans 448 0 0 0 chanx_right_out[17]
port 30 nsew signal tristate
flabel metal2 s 19488 29200 19600 30000 0 FreeSans 448 90 0 0 chanx_right_out[18]
port 31 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chanx_right_out[19]
port 32 nsew signal tristate
flabel metal2 s 11424 29200 11536 30000 0 FreeSans 448 90 0 0 chanx_right_out[1]
port 33 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 chanx_right_out[2]
port 34 nsew signal tristate
flabel metal2 s 14784 29200 14896 30000 0 FreeSans 448 90 0 0 chanx_right_out[3]
port 35 nsew signal tristate
flabel metal2 s 14112 29200 14224 30000 0 FreeSans 448 90 0 0 chanx_right_out[4]
port 36 nsew signal tristate
flabel metal3 s 29200 23520 30000 23632 0 FreeSans 448 0 0 0 chanx_right_out[5]
port 37 nsew signal tristate
flabel metal2 s 17472 29200 17584 30000 0 FreeSans 448 90 0 0 chanx_right_out[6]
port 38 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 chanx_right_out[7]
port 39 nsew signal tristate
flabel metal3 s 29200 22176 30000 22288 0 FreeSans 448 0 0 0 chanx_right_out[8]
port 40 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 chanx_right_out[9]
port 41 nsew signal tristate
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 chany_top_in[0]
port 42 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 chany_top_in[10]
port 43 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 chany_top_in[11]
port 44 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chany_top_in[12]
port 45 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chany_top_in[13]
port 46 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 chany_top_in[14]
port 47 nsew signal input
flabel metal2 s 15456 29200 15568 30000 0 FreeSans 448 90 0 0 chany_top_in[15]
port 48 nsew signal input
flabel metal3 s 29200 5376 30000 5488 0 FreeSans 448 0 0 0 chany_top_in[16]
port 49 nsew signal input
flabel metal2 s 18816 29200 18928 30000 0 FreeSans 448 90 0 0 chany_top_in[17]
port 50 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chany_top_in[18]
port 51 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 chany_top_in[19]
port 52 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 chany_top_in[1]
port 53 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 chany_top_in[2]
port 54 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 chany_top_in[3]
port 55 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 chany_top_in[4]
port 56 nsew signal input
flabel metal2 s 16128 29200 16240 30000 0 FreeSans 448 90 0 0 chany_top_in[5]
port 57 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chany_top_in[6]
port 58 nsew signal input
flabel metal3 s 29200 21504 30000 21616 0 FreeSans 448 0 0 0 chany_top_in[7]
port 59 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chany_top_in[8]
port 60 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 chany_top_in[9]
port 61 nsew signal input
flabel metal3 s 29200 26208 30000 26320 0 FreeSans 448 0 0 0 chany_top_out[0]
port 62 nsew signal tristate
flabel metal2 s 7392 29200 7504 30000 0 FreeSans 448 90 0 0 chany_top_out[10]
port 63 nsew signal tristate
flabel metal3 s 29200 24864 30000 24976 0 FreeSans 448 0 0 0 chany_top_out[11]
port 64 nsew signal tristate
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chany_top_out[12]
port 65 nsew signal tristate
flabel metal2 s 20160 29200 20272 30000 0 FreeSans 448 90 0 0 chany_top_out[13]
port 66 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chany_top_out[14]
port 67 nsew signal tristate
flabel metal3 s 29200 24192 30000 24304 0 FreeSans 448 0 0 0 chany_top_out[15]
port 68 nsew signal tristate
flabel metal3 s 29200 25536 30000 25648 0 FreeSans 448 0 0 0 chany_top_out[16]
port 69 nsew signal tristate
flabel metal2 s 12768 29200 12880 30000 0 FreeSans 448 90 0 0 chany_top_out[17]
port 70 nsew signal tristate
flabel metal2 s 13440 29200 13552 30000 0 FreeSans 448 90 0 0 chany_top_out[18]
port 71 nsew signal tristate
flabel metal2 s 10080 29200 10192 30000 0 FreeSans 448 90 0 0 chany_top_out[19]
port 72 nsew signal tristate
flabel metal2 s 24864 29200 24976 30000 0 FreeSans 448 90 0 0 chany_top_out[1]
port 73 nsew signal tristate
flabel metal2 s 8736 29200 8848 30000 0 FreeSans 448 90 0 0 chany_top_out[2]
port 74 nsew signal tristate
flabel metal3 s 29200 3360 30000 3472 0 FreeSans 448 0 0 0 chany_top_out[3]
port 75 nsew signal tristate
flabel metal3 s 29200 4704 30000 4816 0 FreeSans 448 0 0 0 chany_top_out[4]
port 76 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 chany_top_out[5]
port 77 nsew signal tristate
flabel metal3 s 29200 4032 30000 4144 0 FreeSans 448 0 0 0 chany_top_out[6]
port 78 nsew signal tristate
flabel metal2 s 21504 29200 21616 30000 0 FreeSans 448 90 0 0 chany_top_out[7]
port 79 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 chany_top_out[8]
port 80 nsew signal tristate
flabel metal2 s 16800 29200 16912 30000 0 FreeSans 448 90 0 0 chany_top_out[9]
port 81 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 pReset
port 82 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 prog_clk
port 83 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 84 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 85 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 86 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 87 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 88 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 89 nsew signal input
flabel metal3 s 29200 1344 30000 1456 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 90 nsew signal input
flabel metal3 s 29200 2016 30000 2128 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 91 nsew signal input
flabel metal3 s 29200 7392 30000 7504 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 92 nsew signal input
flabel metal3 s 29200 6720 30000 6832 0 FreeSans 448 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 93 nsew signal input
flabel metal3 s 29200 0 30000 112 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 94 nsew signal input
flabel metal3 s 29200 672 30000 784 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 95 nsew signal input
flabel metal4 s 4586 3076 4906 26716 0 FreeSans 1280 90 0 0 vdd
port 96 nsew power bidirectional
flabel metal4 s 11390 3076 11710 26716 0 FreeSans 1280 90 0 0 vdd
port 96 nsew power bidirectional
flabel metal4 s 18194 3076 18514 26716 0 FreeSans 1280 90 0 0 vdd
port 96 nsew power bidirectional
flabel metal4 s 24998 3076 25318 26716 0 FreeSans 1280 90 0 0 vdd
port 96 nsew power bidirectional
flabel metal4 s 7988 3076 8308 26716 0 FreeSans 1280 90 0 0 vss
port 97 nsew ground bidirectional
flabel metal4 s 14792 3076 15112 26716 0 FreeSans 1280 90 0 0 vss
port 97 nsew ground bidirectional
flabel metal4 s 21596 3076 21916 26716 0 FreeSans 1280 90 0 0 vss
port 97 nsew ground bidirectional
flabel metal4 s 28400 3076 28720 26716 0 FreeSans 1280 90 0 0 vss
port 97 nsew ground bidirectional
rlabel metal1 14952 25872 14952 25872 0 vdd
rlabel via1 15032 26656 15032 26656 0 vss
rlabel metal2 7112 12600 7112 12600 0 _000_
rlabel metal2 4536 11088 4536 11088 0 _001_
rlabel metal2 5600 9240 5600 9240 0 _002_
rlabel metal3 3360 9688 3360 9688 0 _003_
rlabel metal2 11144 11032 11144 11032 0 _004_
rlabel metal2 8232 7168 8232 7168 0 _005_
rlabel metal3 16016 10808 16016 10808 0 _006_
rlabel metal2 11928 11200 11928 11200 0 _007_
rlabel metal2 15568 5992 15568 5992 0 _008_
rlabel metal2 12488 7784 12488 7784 0 _009_
rlabel metal2 20552 9464 20552 9464 0 _010_
rlabel metal2 18648 9632 18648 9632 0 _011_
rlabel metal2 21952 7672 21952 7672 0 _012_
rlabel metal2 24248 9184 24248 9184 0 _013_
rlabel metal2 27776 4872 27776 4872 0 _014_
rlabel metal2 24304 4536 24304 4536 0 _015_
rlabel metal2 26824 8792 26824 8792 0 _016_
rlabel metal3 24024 11592 24024 11592 0 _017_
rlabel metal2 20216 11312 20216 11312 0 _018_
rlabel metal2 18648 11200 18648 11200 0 _019_
rlabel metal2 12040 13552 12040 13552 0 _020_
rlabel metal3 8008 11760 8008 11760 0 _021_
rlabel metal2 4984 14168 4984 14168 0 _022_
rlabel metal2 11816 14280 11816 14280 0 _023_
rlabel metal2 2856 15736 2856 15736 0 _024_
rlabel metal2 8680 14056 8680 14056 0 _025_
rlabel metal2 7560 17248 7560 17248 0 _026_
rlabel metal2 5656 17416 5656 17416 0 _027_
rlabel metal2 11256 17472 11256 17472 0 _028_
rlabel metal2 9576 16352 9576 16352 0 _029_
rlabel metal2 16296 18760 16296 18760 0 _030_
rlabel metal2 13608 19264 13608 19264 0 _031_
rlabel metal2 19880 18144 19880 18144 0 _032_
rlabel metal2 17752 18704 17752 18704 0 _033_
rlabel metal2 24136 18816 24136 18816 0 _034_
rlabel metal2 20776 18928 20776 18928 0 _035_
rlabel metal2 27608 19040 27608 19040 0 _036_
rlabel metal2 26152 20608 26152 20608 0 _037_
rlabel metal2 23464 17024 23464 17024 0 _038_
rlabel metal2 27496 10024 27496 10024 0 _039_
rlabel metal2 12936 16576 12936 16576 0 _040_
rlabel metal2 27832 14336 27832 14336 0 _041_
rlabel metal2 18760 15904 18760 15904 0 _042_
rlabel metal3 18424 15848 18424 15848 0 _043_
rlabel metal2 23016 14168 23016 14168 0 _044_
rlabel metal2 21280 15512 21280 15512 0 _045_
rlabel metal2 27608 10472 27608 10472 0 _046_
rlabel metal2 25928 12824 25928 12824 0 _047_
rlabel metal2 26936 13552 26936 13552 0 _048_
rlabel metal2 6552 7336 6552 7336 0 _049_
rlabel metal3 27440 11256 27440 11256 0 _050_
rlabel metal2 6440 14000 6440 14000 0 _051_
rlabel metal2 27328 20440 27328 20440 0 _052_
rlabel metal3 1302 12152 1302 12152 0 ccff_head
rlabel metal2 27720 15512 27720 15512 0 ccff_tail
rlabel metal2 9912 26600 9912 26600 0 chanx_right_in[0]
rlabel metal2 23016 26152 23016 26152 0 chanx_right_in[10]
rlabel metal2 28168 26152 28168 26152 0 chanx_right_in[17]
rlabel metal2 10808 27426 10808 27426 0 chanx_right_in[18]
rlabel metal2 12096 26488 12096 26488 0 chanx_right_in[19]
rlabel metal3 23898 2744 23898 2744 0 chanx_right_in[7]
rlabel metal3 21560 25480 21560 25480 0 chanx_right_in[8]
rlabel metal2 16352 2184 16352 2184 0 chanx_right_in[9]
rlabel metal2 18984 26208 18984 26208 0 chanx_right_out[16]
rlabel metal2 23128 6272 23128 6272 0 chanx_right_out[17]
rlabel metal2 21224 26320 21224 26320 0 chanx_right_out[18]
rlabel metal2 13496 2030 13496 2030 0 chanx_right_out[19]
rlabel metal2 19096 26320 19096 26320 0 chanx_right_out[6]
rlabel metal2 21056 3640 21056 3640 0 chanx_right_out[7]
rlabel metal3 28658 22232 28658 22232 0 chanx_right_out[8]
rlabel metal3 21336 3640 21336 3640 0 chanx_right_out[9]
rlabel metal2 15568 26264 15568 26264 0 chany_top_in[15]
rlabel metal3 28070 5432 28070 5432 0 chany_top_in[16]
rlabel metal2 19656 26208 19656 26208 0 chany_top_in[17]
rlabel metal2 12208 3416 12208 3416 0 chany_top_in[18]
rlabel metal2 16240 26264 16240 26264 0 chany_top_in[5]
rlabel metal3 21280 3528 21280 3528 0 chany_top_in[6]
rlabel metal2 28168 22344 28168 22344 0 chany_top_in[7]
rlabel metal2 19096 2520 19096 2520 0 chany_top_in[8]
rlabel metal2 27720 25872 27720 25872 0 chany_top_out[16]
rlabel metal2 13944 25648 13944 25648 0 chany_top_out[17]
rlabel metal2 14168 26992 14168 26992 0 chany_top_out[18]
rlabel metal2 11144 26656 11144 26656 0 chany_top_out[19]
rlabel metal3 28070 4088 28070 4088 0 chany_top_out[6]
rlabel metal2 22792 26488 22792 26488 0 chany_top_out[7]
rlabel metal2 15512 2058 15512 2058 0 chany_top_out[8]
rlabel metal2 17528 26488 17528 26488 0 chany_top_out[9]
rlabel metal2 14504 13720 14504 13720 0 clknet_0_prog_clk
rlabel metal2 5656 10976 5656 10976 0 clknet_2_0__leaf_prog_clk
rlabel metal3 3584 16856 3584 16856 0 clknet_2_1__leaf_prog_clk
rlabel metal2 28168 11480 28168 11480 0 clknet_2_2__leaf_prog_clk
rlabel metal2 22904 20776 22904 20776 0 clknet_2_3__leaf_prog_clk
rlabel metal2 4200 14672 4200 14672 0 mem_right_track_0.DFFR_0_.D
rlabel metal2 3080 14336 3080 14336 0 mem_right_track_0.DFFR_0_.Q
rlabel metal2 2072 16240 2072 16240 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 23576 17864 23576 17864 0 mem_right_track_10.DFFR_0_.D
rlabel metal3 24864 20104 24864 20104 0 mem_right_track_10.DFFR_0_.Q
rlabel metal3 26096 21672 26096 21672 0 mem_right_track_10.DFFR_1_.Q
rlabel metal3 7224 18536 7224 18536 0 mem_right_track_2.DFFR_0_.Q
rlabel metal2 8344 18032 8344 18032 0 mem_right_track_2.DFFR_1_.Q
rlabel metal2 26712 20356 26712 20356 0 mem_right_track_20.DFFR_0_.Q
rlabel metal2 28280 18200 28280 18200 0 mem_right_track_20.DFFR_1_.Q
rlabel metal2 28280 10080 28280 10080 0 mem_right_track_22.DFFR_0_.Q
rlabel metal3 24696 15400 24696 15400 0 mem_right_track_22.DFFR_1_.Q
rlabel metal2 19992 16464 19992 16464 0 mem_right_track_24.DFFR_0_.Q
rlabel metal3 15288 16968 15288 16968 0 mem_right_track_24.DFFR_1_.Q
rlabel metal3 18200 15960 18200 15960 0 mem_right_track_26.DFFR_0_.Q
rlabel metal3 21504 15400 21504 15400 0 mem_right_track_26.DFFR_1_.Q
rlabel metal2 27496 14560 27496 14560 0 mem_right_track_28.DFFR_0_.Q
rlabel metal2 27272 15848 27272 15848 0 mem_right_track_28.DFFR_1_.Q
rlabel metal2 27384 5992 27384 5992 0 mem_right_track_30.DFFR_0_.Q
rlabel metal2 10360 17248 10360 17248 0 mem_right_track_4.DFFR_0_.Q
rlabel metal2 11816 18480 11816 18480 0 mem_right_track_4.DFFR_1_.Q
rlabel metal2 14168 19264 14168 19264 0 mem_right_track_6.DFFR_0_.Q
rlabel metal3 18200 19096 18200 19096 0 mem_right_track_6.DFFR_1_.Q
rlabel metal2 23240 18592 23240 18592 0 mem_right_track_8.DFFR_0_.Q
rlabel metal2 5320 11032 5320 11032 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 8456 11872 8456 11872 0 mem_top_track_0.DFFR_1_.Q
rlabel metal3 17528 8120 17528 8120 0 mem_top_track_10.DFFR_0_.D
rlabel metal2 23576 9352 23576 9352 0 mem_top_track_10.DFFR_0_.Q
rlabel metal3 22400 8120 22400 8120 0 mem_top_track_10.DFFR_1_.Q
rlabel metal2 1624 7896 1624 7896 0 mem_top_track_2.DFFR_0_.Q
rlabel metal3 6608 7560 6608 7560 0 mem_top_track_2.DFFR_1_.Q
rlabel metal2 27160 9352 27160 9352 0 mem_top_track_20.DFFR_0_.Q
rlabel metal3 21840 5992 21840 5992 0 mem_top_track_20.DFFR_1_.Q
rlabel metal2 24808 4760 24808 4760 0 mem_top_track_22.DFFR_0_.Q
rlabel metal2 27496 3752 27496 3752 0 mem_top_track_22.DFFR_1_.Q
rlabel metal2 24920 6412 24920 6412 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 27496 7896 27496 7896 0 mem_top_track_24.DFFR_1_.Q
rlabel metal3 27272 11424 27272 11424 0 mem_top_track_26.DFFR_0_.Q
rlabel metal3 16800 7560 16800 7560 0 mem_top_track_26.DFFR_1_.Q
rlabel metal2 7224 11760 7224 11760 0 mem_top_track_28.DFFR_0_.Q
rlabel metal2 19432 13496 19432 13496 0 mem_top_track_28.DFFR_1_.Q
rlabel metal2 8792 13160 8792 13160 0 mem_top_track_30.DFFR_0_.Q
rlabel metal2 8904 9352 8904 9352 0 mem_top_track_4.DFFR_0_.Q
rlabel metal2 9520 9800 9520 9800 0 mem_top_track_4.DFFR_1_.Q
rlabel metal2 9352 10360 9352 10360 0 mem_top_track_6.DFFR_0_.Q
rlabel metal2 15848 8456 15848 8456 0 mem_top_track_6.DFFR_1_.Q
rlabel metal3 9744 9128 9744 9128 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 2072 11648 2072 11648 0 net1
rlabel metal2 15400 24024 15400 24024 0 net10
rlabel metal2 4760 7896 4760 7896 0 net100
rlabel metal2 25872 17080 25872 17080 0 net101
rlabel metal3 13496 8232 13496 8232 0 net102
rlabel metal2 20832 16856 20832 16856 0 net103
rlabel metal2 11144 16744 11144 16744 0 net104
rlabel metal2 21448 12152 21448 12152 0 net105
rlabel metal2 16240 11368 16240 11368 0 net106
rlabel metal2 19432 5544 19432 5544 0 net11
rlabel metal2 18928 23912 18928 23912 0 net12
rlabel metal2 12600 4648 12600 4648 0 net13
rlabel metal2 16072 24024 16072 24024 0 net14
rlabel metal2 19936 3416 19936 3416 0 net15
rlabel metal2 27664 23240 27664 23240 0 net16
rlabel metal2 19096 3864 19096 3864 0 net17
rlabel metal2 14392 18032 14392 18032 0 net18
rlabel metal2 28336 9800 28336 9800 0 net19
rlabel metal2 9352 25144 9352 25144 0 net2
rlabel metal3 17192 21784 17192 21784 0 net20
rlabel metal2 19656 5712 19656 5712 0 net21
rlabel metal2 20776 25816 20776 25816 0 net22
rlabel metal2 14280 4760 14280 4760 0 net23
rlabel metal3 17584 21672 17584 21672 0 net24
rlabel metal3 20720 3416 20720 3416 0 net25
rlabel metal2 27160 22792 27160 22792 0 net26
rlabel metal2 22680 3976 22680 3976 0 net27
rlabel metal2 27048 25592 27048 25592 0 net28
rlabel metal2 13160 25088 13160 25088 0 net29
rlabel metal2 22680 25480 22680 25480 0 net3
rlabel metal2 12936 25816 12936 25816 0 net30
rlabel metal2 9576 24528 9576 24528 0 net31
rlabel metal2 21672 6608 21672 6608 0 net32
rlabel metal2 21672 25816 21672 25816 0 net33
rlabel metal2 15176 3976 15176 3976 0 net34
rlabel metal2 16744 25816 16744 25816 0 net35
rlabel metal2 28168 24528 28168 24528 0 net36
rlabel metal2 17808 4424 17808 4424 0 net37
rlabel metal2 20664 26320 20664 26320 0 net38
rlabel metal2 14168 2590 14168 2590 0 net39
rlabel metal2 27496 24808 27496 24808 0 net4
rlabel metal3 27496 25088 27496 25088 0 net40
rlabel metal2 7560 26488 7560 26488 0 net41
rlabel metal2 12824 1190 12824 1190 0 net42
rlabel metal2 28168 6832 28168 6832 0 net43
rlabel metal2 28168 3920 28168 3920 0 net44
rlabel metal2 8792 27874 8792 27874 0 net45
rlabel metal2 25032 26488 25032 26488 0 net46
rlabel metal2 26264 26320 26264 26320 0 net47
rlabel metal2 21560 1582 21560 1582 0 net48
rlabel metal2 24920 2030 24920 2030 0 net49
rlabel metal2 12824 25032 12824 25032 0 net5
rlabel metal2 16856 1246 16856 1246 0 net50
rlabel metal2 8064 26488 8064 26488 0 net51
rlabel metal3 23408 26488 23408 26488 0 net52
rlabel metal2 14840 1862 14840 1862 0 net53
rlabel metal3 28280 23688 28280 23688 0 net54
rlabel metal3 13720 26488 13720 26488 0 net55
rlabel metal2 15064 25928 15064 25928 0 net56
rlabel metal3 1246 24920 1246 24920 0 net57
rlabel metal2 11704 25536 11704 25536 0 net58
rlabel metal2 28224 23688 28224 23688 0 net59
rlabel metal2 12600 25928 12600 25928 0 net6
rlabel metal2 20440 12208 20440 12208 0 net60
rlabel metal2 14280 13664 14280 13664 0 net61
rlabel metal3 17304 16184 17304 16184 0 net62
rlabel metal2 16184 9072 16184 9072 0 net63
rlabel metal2 15512 18480 15512 18480 0 net64
rlabel metal2 4088 12992 4088 12992 0 net65
rlabel metal2 20776 13664 20776 13664 0 net66
rlabel metal2 14056 16408 14056 16408 0 net67
rlabel metal3 12152 10472 12152 10472 0 net68
rlabel metal2 14056 19544 14056 19544 0 net69
rlabel metal2 18760 3332 18760 3332 0 net7
rlabel metal2 6216 8568 6216 8568 0 net70
rlabel metal2 11480 8960 11480 8960 0 net71
rlabel metal2 26208 16744 26208 16744 0 net72
rlabel metal3 24304 5208 24304 5208 0 net73
rlabel metal2 17864 18368 17864 18368 0 net74
rlabel metal2 21896 19544 21896 19544 0 net75
rlabel metal2 11144 18872 11144 18872 0 net76
rlabel metal3 21420 15176 21420 15176 0 net77
rlabel metal3 11760 9800 11760 9800 0 net78
rlabel metal2 7336 13384 7336 13384 0 net79
rlabel metal3 21728 25256 21728 25256 0 net8
rlabel metal2 18200 8960 18200 8960 0 net80
rlabel metal2 7336 16912 7336 16912 0 net81
rlabel metal2 4088 14952 4088 14952 0 net82
rlabel metal2 3864 11928 3864 11928 0 net83
rlabel metal2 20664 9912 20664 9912 0 net84
rlabel metal2 5320 17584 5320 17584 0 net85
rlabel metal2 26432 15176 26432 15176 0 net86
rlabel metal2 8008 15008 8008 15008 0 net87
rlabel metal2 23688 21112 23688 21112 0 net88
rlabel metal3 3248 8344 3248 8344 0 net89
rlabel metal2 16968 3864 16968 3864 0 net9
rlabel metal2 19432 18872 19432 18872 0 net90
rlabel metal2 8792 18760 8792 18760 0 net91
rlabel metal2 24248 7392 24248 7392 0 net92
rlabel metal2 21560 5544 21560 5544 0 net93
rlabel metal2 2968 17584 2968 17584 0 net94
rlabel metal2 6104 9744 6104 9744 0 net95
rlabel metal2 25704 17640 25704 17640 0 net96
rlabel metal2 14784 7336 14784 7336 0 net97
rlabel metal2 24472 5768 24472 5768 0 net98
rlabel metal2 25368 8232 25368 8232 0 net99
rlabel metal2 1736 17136 1736 17136 0 pReset
rlabel metal3 2478 19544 2478 19544 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
