// This is the unpowered netlist.
module sb_0__1_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input [19:0] chanx_right_in;
 output [19:0] chanx_right_out;
 input [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;
 input [19:0] chany_top_in;
 output [19:0] chany_top_out;

 wire net97;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net81;
 wire net78;
 wire net77;
 wire net80;
 wire net79;
 wire net76;
 wire net73;
 wire net72;
 wire net75;
 wire net74;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire clknet_0_prog_clk;
 wire clknet_3_0__leaf_prog_clk;
 wire clknet_3_1__leaf_prog_clk;
 wire clknet_3_2__leaf_prog_clk;
 wire clknet_3_3__leaf_prog_clk;
 wire clknet_3_4__leaf_prog_clk;
 wire clknet_3_5__leaf_prog_clk;
 wire clknet_3_6__leaf_prog_clk;
 wire clknet_3_7__leaf_prog_clk;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_1.DFFR_2_.Q ;
 wire \mem_bottom_track_1.DFFR_3_.Q ;
 wire \mem_bottom_track_1.DFFR_4_.Q ;
 wire \mem_bottom_track_1.DFFR_5_.Q ;
 wire \mem_bottom_track_1.DFFR_6_.Q ;
 wire \mem_bottom_track_1.DFFR_7_.Q ;
 wire \mem_bottom_track_17.DFFR_0_.D ;
 wire \mem_bottom_track_17.DFFR_0_.Q ;
 wire \mem_bottom_track_17.DFFR_1_.Q ;
 wire \mem_bottom_track_17.DFFR_2_.Q ;
 wire \mem_bottom_track_17.DFFR_3_.Q ;
 wire \mem_bottom_track_17.DFFR_4_.Q ;
 wire \mem_bottom_track_17.DFFR_5_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_2_.Q ;
 wire \mem_bottom_track_25.DFFR_3_.Q ;
 wire \mem_bottom_track_25.DFFR_4_.Q ;
 wire \mem_bottom_track_25.DFFR_5_.Q ;
 wire \mem_bottom_track_33.DFFR_0_.Q ;
 wire \mem_bottom_track_33.DFFR_1_.Q ;
 wire \mem_bottom_track_33.DFFR_2_.Q ;
 wire \mem_bottom_track_33.DFFR_3_.Q ;
 wire \mem_bottom_track_33.DFFR_4_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_bottom_track_9.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_2_.Q ;
 wire \mem_bottom_track_9.DFFR_3_.Q ;
 wire \mem_bottom_track_9.DFFR_4_.Q ;
 wire \mem_right_track_0.DFFR_0_.D ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_10.DFFR_0_.D ;
 wire \mem_right_track_10.DFFR_0_.Q ;
 wire \mem_right_track_10.DFFR_1_.Q ;
 wire \mem_right_track_12.DFFR_0_.Q ;
 wire \mem_right_track_12.DFFR_1_.Q ;
 wire \mem_right_track_14.DFFR_0_.Q ;
 wire \mem_right_track_14.DFFR_1_.Q ;
 wire \mem_right_track_16.DFFR_0_.Q ;
 wire \mem_right_track_16.DFFR_1_.Q ;
 wire \mem_right_track_18.DFFR_0_.Q ;
 wire \mem_right_track_18.DFFR_1_.Q ;
 wire \mem_right_track_2.DFFR_0_.Q ;
 wire \mem_right_track_2.DFFR_1_.Q ;
 wire \mem_right_track_2.DFFR_2_.Q ;
 wire \mem_right_track_2.DFFR_3_.Q ;
 wire \mem_right_track_2.DFFR_4_.Q ;
 wire \mem_right_track_2.DFFR_5_.Q ;
 wire \mem_right_track_20.DFFR_0_.Q ;
 wire \mem_right_track_20.DFFR_1_.Q ;
 wire \mem_right_track_22.DFFR_0_.Q ;
 wire \mem_right_track_22.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_26.DFFR_0_.Q ;
 wire \mem_right_track_26.DFFR_1_.Q ;
 wire \mem_right_track_28.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_1_.Q ;
 wire \mem_right_track_4.DFFR_2_.Q ;
 wire \mem_right_track_4.DFFR_3_.Q ;
 wire \mem_right_track_4.DFFR_4_.Q ;
 wire \mem_right_track_4.DFFR_5_.Q ;
 wire \mem_right_track_6.DFFR_0_.Q ;
 wire \mem_right_track_6.DFFR_1_.Q ;
 wire \mem_right_track_6.DFFR_2_.Q ;
 wire \mem_right_track_6.DFFR_3_.Q ;
 wire \mem_right_track_6.DFFR_4_.Q ;
 wire \mem_right_track_6.DFFR_5_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_0.DFFR_2_.Q ;
 wire \mem_top_track_0.DFFR_3_.Q ;
 wire \mem_top_track_0.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_5_.Q ;
 wire \mem_top_track_0.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_7_.Q ;
 wire \mem_top_track_16.DFFR_0_.D ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_2_.Q ;
 wire \mem_top_track_16.DFFR_3_.Q ;
 wire \mem_top_track_16.DFFR_4_.Q ;
 wire \mem_top_track_16.DFFR_5_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_2_.Q ;
 wire \mem_top_track_24.DFFR_3_.Q ;
 wire \mem_top_track_24.DFFR_4_.Q ;
 wire \mem_top_track_24.DFFR_5_.Q ;
 wire \mem_top_track_32.DFFR_0_.Q ;
 wire \mem_top_track_32.DFFR_1_.Q ;
 wire \mem_top_track_32.DFFR_2_.Q ;
 wire \mem_top_track_32.DFFR_3_.Q ;
 wire \mem_top_track_32.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire \mem_top_track_8.DFFR_1_.Q ;
 wire \mem_top_track_8.DFFR_2_.Q ;
 wire \mem_top_track_8.DFFR_3_.Q ;
 wire \mem_top_track_8.DFFR_4_.Q ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net8;
 wire net9;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__122__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__130__I (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__133__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__I (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__I (.I(_113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__I (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__221__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__I (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__RN (.I(_005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__RN (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__244__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__CLK (.I(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__CLK (.I(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__CLK (.I(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__374__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__380__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(chany_bottom_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(chany_bottom_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(chany_bottom_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(chany_bottom_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(chany_bottom_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(chany_bottom_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(chany_bottom_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(chany_bottom_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(chany_bottom_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(chany_bottom_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(chany_bottom_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(chany_top_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(chany_top_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(chany_top_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(chany_top_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(chany_top_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(chany_top_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(chany_top_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(chany_top_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(chany_top_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(chany_bottom_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(chany_top_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(chany_top_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(chany_top_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(chany_top_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(chany_top_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(chany_top_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(chany_bottom_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(chany_bottom_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(chany_bottom_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(chany_bottom_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(chany_bottom_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(chany_bottom_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(chany_bottom_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_108 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _118_ (.I(net36),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _119_ (.I(_106_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _120_ (.I(_107_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _121_ (.I(_108_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _122_ (.I(_108_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _123_ (.I(_108_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _124_ (.I(_108_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _125_ (.I(_108_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _126_ (.I(_108_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _127_ (.I(_108_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _128_ (.I(_108_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _129_ (.I(_108_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _130_ (.I(_108_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _131_ (.I(_107_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _132_ (.I(_109_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _133_ (.I(_109_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _134_ (.I(_109_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _135_ (.I(_109_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _136_ (.I(_109_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _137_ (.I(_109_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _138_ (.I(_109_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _139_ (.I(_109_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _140_ (.I(_109_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _141_ (.I(_109_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _142_ (.I(_107_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _143_ (.I(_110_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _144_ (.I(_110_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _145_ (.I(_110_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _146_ (.I(_110_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _147_ (.I(_110_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _148_ (.I(_110_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _149_ (.I(_110_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _150_ (.I(_110_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _151_ (.I(_110_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _152_ (.I(_110_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _153_ (.I(_107_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _154_ (.I(_111_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _155_ (.I(_111_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _156_ (.I(_111_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _157_ (.I(_111_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _158_ (.I(_111_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _159_ (.I(_111_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _160_ (.I(_111_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _161_ (.I(_111_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _162_ (.I(_111_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _163_ (.I(_111_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _164_ (.I(_106_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _165_ (.I(_112_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _166_ (.I(_112_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _167_ (.I(_112_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _168_ (.I(_112_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _169_ (.I(_112_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _170_ (.I(_112_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _171_ (.I(_112_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _172_ (.I(_112_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _173_ (.I(_112_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _174_ (.I(_112_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _175_ (.I(_106_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _176_ (.I(_113_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _177_ (.I(_113_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _178_ (.I(_113_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _179_ (.I(_113_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _180_ (.I(_113_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _181_ (.I(_113_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _182_ (.I(_113_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _183_ (.I(_113_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _184_ (.I(_113_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _185_ (.I(_113_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _186_ (.I(_106_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _187_ (.I(_114_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _188_ (.I(_114_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _189_ (.I(_114_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _190_ (.I(_114_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _191_ (.I(_114_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _192_ (.I(_114_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _193_ (.I(_114_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _194_ (.I(_114_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _195_ (.I(_114_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _196_ (.I(_114_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _197_ (.I(_106_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _198_ (.I(_115_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _199_ (.I(_115_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _200_ (.I(_115_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _201_ (.I(_115_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _202_ (.I(_115_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _203_ (.I(_115_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _204_ (.I(_115_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _205_ (.I(_115_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _206_ (.I(_115_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _207_ (.I(_115_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _208_ (.I(_106_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _209_ (.I(_116_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _210_ (.I(_116_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _211_ (.I(_116_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _212_ (.I(_116_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _213_ (.I(_116_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _214_ (.I(_116_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _215_ (.I(_116_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _216_ (.I(_116_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _217_ (.I(_116_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _218_ (.I(_116_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _219_ (.I(_106_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _220_ (.I(_117_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _221_ (.I(_117_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _222_ (.I(_117_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _223_ (.I(_117_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _224_ (.I(_117_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _225_ (.I(_117_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _226_ (.I(_117_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _227_ (.I(_117_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _228_ (.I(_117_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _229_ (.I(_117_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _230_ (.I(_107_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _231_ (.I(_107_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _232_ (.I(_107_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _233_ (.I(_107_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _234_ (.I(_107_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _235_ (.I(_107_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _236_ (.D(net146),
    .RN(_000_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _237_ (.D(net161),
    .RN(_001_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _238_ (.D(net119),
    .RN(_002_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _239_ (.D(net166),
    .RN(_003_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _240_ (.D(net138),
    .RN(_004_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _241_ (.D(net169),
    .RN(_005_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _242_ (.D(net198),
    .RN(_006_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _243_ (.D(net1),
    .RN(_007_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _244_ (.D(net139),
    .RN(_008_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _245_ (.D(net123),
    .RN(_009_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _246_ (.D(net148),
    .RN(_010_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _247_ (.D(net136),
    .RN(_011_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _248_ (.D(net193),
    .RN(_012_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _249_ (.D(net151),
    .RN(_013_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _250_ (.D(net155),
    .RN(_014_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _251_ (.D(net129),
    .RN(_015_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _252_ (.D(net174),
    .RN(_016_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _253_ (.D(net145),
    .RN(_017_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _254_ (.D(net105),
    .RN(_018_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _255_ (.D(net189),
    .RN(_019_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _256_ (.D(net181),
    .RN(_020_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _257_ (.D(net116),
    .RN(_021_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _258_ (.D(net128),
    .RN(_022_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _259_ (.D(net117),
    .RN(_023_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _260_ (.D(net137),
    .RN(_024_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _261_ (.D(net162),
    .RN(_025_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _262_ (.D(net120),
    .RN(_026_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _263_ (.D(net143),
    .RN(_027_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _264_ (.D(net122),
    .RN(_028_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _265_ (.D(net199),
    .RN(_029_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _266_ (.D(net147),
    .RN(_030_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _267_ (.D(net184),
    .RN(_031_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _268_ (.D(net104),
    .RN(_032_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _269_ (.D(net163),
    .RN(_033_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _270_ (.D(net164),
    .RN(_034_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _271_ (.D(net194),
    .RN(_035_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _272_ (.D(net187),
    .RN(_036_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _273_ (.D(net171),
    .RN(_037_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _274_ (.D(net112),
    .RN(_038_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _275_ (.D(net130),
    .RN(_039_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _276_ (.D(net102),
    .RN(_040_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _277_ (.D(net182),
    .RN(_041_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _278_ (.D(net132),
    .RN(_042_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _279_ (.D(net121),
    .RN(_043_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _280_ (.D(net177),
    .RN(_044_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _281_ (.D(net170),
    .RN(_045_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _282_ (.D(net131),
    .RN(_046_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _283_ (.D(net150),
    .RN(_047_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _284_ (.D(net101),
    .RN(_048_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _285_ (.D(net190),
    .RN(_049_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _286_ (.D(net167),
    .RN(_050_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _287_ (.D(net173),
    .RN(_051_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _288_ (.D(net195),
    .RN(_052_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _289_ (.D(net197),
    .RN(_053_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _290_ (.D(net124),
    .RN(_054_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _291_ (.D(net108),
    .RN(_055_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _292_ (.D(net157),
    .RN(_056_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _293_ (.D(net115),
    .RN(_057_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _294_ (.D(net192),
    .RN(_058_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _295_ (.D(net183),
    .RN(_059_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _296_ (.D(net134),
    .RN(_060_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _297_ (.D(net118),
    .RN(_061_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _298_ (.D(net127),
    .RN(_062_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _299_ (.D(net201),
    .RN(_063_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _300_ (.D(net159),
    .RN(_064_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _301_ (.D(net202),
    .RN(_065_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _302_ (.D(net107),
    .RN(_066_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_10.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _303_ (.D(net152),
    .RN(_067_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _304_ (.D(net135),
    .RN(_068_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_10.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _305_ (.D(net172),
    .RN(_069_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_10.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _306_ (.D(net142),
    .RN(_070_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_20.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _307_ (.D(net191),
    .RN(_071_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_20.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _308_ (.D(net98),
    .RN(_072_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_right_track_22.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _309_ (.D(net196),
    .RN(_073_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_22.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _310_ (.D(net165),
    .RN(_074_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _311_ (.D(net125),
    .RN(_075_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _312_ (.D(net110),
    .RN(_076_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_26.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _313_ (.D(net144),
    .RN(_077_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_26.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _314_ (.D(net106),
    .RN(_078_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _315_ (.D(net168),
    .RN(_079_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_28.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _316_ (.D(net111),
    .RN(_080_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _317_ (.D(net149),
    .RN(_081_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _318_ (.D(net160),
    .RN(_082_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _319_ (.D(net141),
    .RN(_083_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _320_ (.D(net100),
    .RN(_084_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _321_ (.D(net185),
    .RN(_085_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_2.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _322_ (.D(net113),
    .RN(_086_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _323_ (.D(net99),
    .RN(_087_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _324_ (.D(net178),
    .RN(_088_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _325_ (.D(net126),
    .RN(_089_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _326_ (.D(net153),
    .RN(_090_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _327_ (.D(net188),
    .RN(_091_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_4.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _328_ (.D(net140),
    .RN(_092_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _329_ (.D(net114),
    .RN(_093_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _330_ (.D(net133),
    .RN(_094_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _331_ (.D(net176),
    .RN(_095_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _332_ (.D(net156),
    .RN(_096_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _333_ (.D(net180),
    .RN(_097_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_6.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _334_ (.D(net158),
    .RN(_098_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_12.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _335_ (.D(net200),
    .RN(_099_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_12.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _336_ (.D(net154),
    .RN(_100_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_14.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _337_ (.D(net175),
    .RN(_101_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_right_track_14.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _338_ (.D(net179),
    .RN(_102_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _339_ (.D(net103),
    .RN(_103_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _340_ (.D(net109),
    .RN(_104_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_right_track_18.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _341_ (.D(net186),
    .RN(_105_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_right_track_18.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _368_ (.I(net14),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _369_ (.I(net18),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _370_ (.I(net4),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _371_ (.I(net8),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _372_ (.I(net28),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _373_ (.I(net27),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _374_ (.I(net26),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _375_ (.I(net25),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _376_ (.I(net24),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _377_ (.I(net23),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _378_ (.I(net22),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _379_ (.I(net35),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _380_ (.I(net34),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _381_ (.I(net33),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _382_ (.I(net32),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _383_ (.I(net31),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _384_ (.I(net30),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _385_ (.I(net29),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _386_ (.I(net21),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _387_ (.I(net11),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _388_ (.I(net10),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _389_ (.I(net9),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _390_ (.I(net7),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _391_ (.I(net6),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _392_ (.I(net5),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _393_ (.I(net3),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _394_ (.I(net20),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _395_ (.I(net19),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _396_ (.I(net17),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _397_ (.I(net16),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _398_ (.I(net15),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _399_ (.I(net13),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _400_ (.I(net12),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _401_ (.I(net2),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_4__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\mem_right_track_22.DFFR_0_.Q ),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\mem_right_track_8.DFFR_0_.Q ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(\mem_bottom_track_25.DFFR_3_.Q ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(\mem_top_track_0.DFFR_0_.Q ),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(\mem_top_track_24.DFFR_3_.Q ),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(\mem_right_track_10.DFFR_1_.Q ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(\mem_bottom_track_25.DFFR_5_.Q ),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(\mem_right_track_0.DFFR_0_.D ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\mem_bottom_track_25.DFFR_1_.Q ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\mem_right_track_18.DFFR_0_.Q ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\mem_right_track_26.DFFR_0_.Q ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\mem_right_track_2.DFFR_4_.Q ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\mem_top_track_32.DFFR_0_.Q ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\mem_right_track_4.DFFR_4_.Q ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\mem_right_track_6.DFFR_3_.Q ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\mem_bottom_track_17.DFFR_5_.Q ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\mem_top_track_0.DFFR_7_.Q ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\mem_right_track_4.DFFR_3_.Q ),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\mem_top_track_16.DFFR_3_.Q ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\mem_bottom_track_33.DFFR_1_.Q ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\mem_top_track_0.DFFR_4_.Q ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\mem_top_track_16.DFFR_0_.Q ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\mem_bottom_track_9.DFFR_1_.Q ),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\mem_top_track_24.DFFR_4_.Q ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\mem_bottom_track_1.DFFR_5_.Q ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\mem_bottom_track_25.DFFR_2_.Q ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\mem_right_track_22.DFFR_1_.Q ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\mem_right_track_4.DFFR_1_.Q ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\mem_right_track_2.DFFR_0_.Q ),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\mem_bottom_track_33.DFFR_0_.Q ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\mem_top_track_16.DFFR_4_.Q ),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\mem_bottom_track_1.DFFR_0_.D ),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\mem_top_track_24.DFFR_5_.Q ),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\mem_bottom_track_17.DFFR_4_.Q ),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\mem_bottom_track_9.DFFR_2_.Q ),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\mem_right_track_6.DFFR_2_.Q ),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\mem_bottom_track_33.DFFR_2_.Q ),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\mem_right_track_10.DFFR_0_.Q ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\mem_bottom_track_1.DFFR_3_.Q ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\mem_bottom_track_17.DFFR_2_.Q ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\mem_top_track_16.DFFR_2_.Q ),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\mem_top_track_0.DFFR_2_.Q ),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\mem_bottom_track_1.DFFR_6_.Q ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\mem_right_track_6.DFFR_4_.Q ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\mem_right_track_2.DFFR_1_.Q ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\mem_right_track_20.DFFR_0_.Q ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\mem_top_track_16.DFFR_0_.D ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\mem_right_track_24.DFFR_1_.Q ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(\mem_top_track_8.DFFR_3_.Q ),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\mem_top_track_0.DFFR_6_.Q ),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\mem_bottom_track_9.DFFR_4_.Q ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(\mem_top_track_24.DFFR_2_.Q ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\mem_bottom_track_1.DFFR_4_.Q ),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(\mem_right_track_2.DFFR_3_.Q ),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\mem_bottom_track_17.DFFR_3_.Q ),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(\mem_bottom_track_1.DFFR_1_.Q ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\mem_right_track_6.DFFR_5_.Q ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(\mem_right_track_4.DFFR_0_.Q ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\mem_right_track_14.DFFR_0_.Q ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(\mem_bottom_track_1.DFFR_0_.Q ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\mem_right_track_6.DFFR_0_.Q ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\mem_right_track_14.DFFR_1_.Q ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(\mem_bottom_track_25.DFFR_0_.Q ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\mem_right_track_12.DFFR_0_.Q ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(\mem_right_track_0.DFFR_0_.Q ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\mem_right_track_2.DFFR_2_.Q ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(\mem_top_track_0.DFFR_5_.Q ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\mem_top_track_16.DFFR_1_.Q ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(\mem_top_track_16.DFFR_5_.Q ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\mem_top_track_32.DFFR_4_.Q ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(\mem_right_track_24.DFFR_0_.Q ),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\mem_top_track_0.DFFR_3_.Q ),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\mem_top_track_24.DFFR_0_.Q ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(\mem_bottom_track_17.DFFR_0_.Q ),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\mem_right_track_26.DFFR_1_.Q ),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(\mem_top_track_0.DFFR_1_.Q ),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\mem_bottom_track_1.DFFR_7_.Q ),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(\mem_top_track_32.DFFR_1_.Q ),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\mem_right_track_10.DFFR_0_.D ),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(\mem_bottom_track_17.DFFR_0_.D ),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\mem_top_track_8.DFFR_4_.Q ),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(\mem_right_track_12.DFFR_1_.Q ),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\mem_right_track_6.DFFR_1_.Q ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\mem_top_track_8.DFFR_2_.Q ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(\mem_bottom_track_9.DFFR_0_.Q ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\mem_right_track_4.DFFR_2_.Q ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(\mem_right_track_16.DFFR_0_.Q ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\mem_right_track_4.DFFR_5_.Q ),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(\mem_top_track_8.DFFR_0_.Q ),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\mem_bottom_track_9.DFFR_3_.Q ),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(\mem_bottom_track_33.DFFR_3_.Q ),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\mem_top_track_24.DFFR_1_.Q ),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(\mem_right_track_0.DFFR_1_.Q ),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\mem_right_track_16.DFFR_1_.Q ),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\mem_right_track_28.DFFR_0_.Q ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(\mem_top_track_32.DFFR_2_.Q ),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\mem_right_track_2.DFFR_5_.Q ),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(\mem_top_track_8.DFFR_1_.Q ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\mem_bottom_track_17.DFFR_1_.Q ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(\mem_right_track_18.DFFR_1_.Q ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(\mem_bottom_track_33.DFFR_4_.Q ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(\mem_bottom_track_1.DFFR_2_.Q ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(\mem_top_track_32.DFFR_3_.Q ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(\mem_bottom_track_25.DFFR_4_.Q ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(\mem_right_track_20.DFFR_1_.Q ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(chany_bottom_in[17]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(chany_bottom_in[18]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(chany_bottom_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(chany_bottom_in[2]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(chany_bottom_in[3]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(chany_bottom_in[4]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(chany_bottom_in[5]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(chany_bottom_in[6]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(chany_bottom_in[7]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(chany_bottom_in[8]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(chany_bottom_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(chany_bottom_in[9]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(chany_top_in[0]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(chany_top_in[10]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(chany_top_in[12]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(chany_top_in[13]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(chany_top_in[14]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(chany_top_in[16]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(chany_top_in[17]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(chany_top_in[18]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(chany_top_in[1]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(chany_bottom_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(chany_top_in[2]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(chany_top_in[4]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(chany_top_in[5]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(chany_top_in[6]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(chany_top_in[8]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(chany_top_in[9]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(pReset),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(chany_bottom_in[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(chany_bottom_in[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(chany_bottom_in[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(chany_bottom_in[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(chany_bottom_in[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(chany_bottom_in[16]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(chanx_right_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output39 (.I(net39),
    .Z(chanx_right_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output40 (.I(net40),
    .Z(chanx_right_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output41 (.I(net41),
    .Z(chanx_right_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output42 (.I(net42),
    .Z(chany_bottom_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output43 (.I(net43),
    .Z(chany_bottom_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output44 (.I(net44),
    .Z(chany_bottom_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output45 (.I(net45),
    .Z(chany_bottom_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output46 (.I(net46),
    .Z(chany_bottom_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output47 (.I(net47),
    .Z(chany_bottom_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output48 (.I(net48),
    .Z(chany_bottom_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output49 (.I(net49),
    .Z(chany_bottom_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output50 (.I(net50),
    .Z(chany_bottom_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output51 (.I(net51),
    .Z(chany_bottom_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output52 (.I(net52),
    .Z(chany_bottom_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output53 (.I(net53),
    .Z(chany_bottom_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output54 (.I(net54),
    .Z(chany_bottom_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output55 (.I(net55),
    .Z(chany_bottom_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output56 (.I(net56),
    .Z(chany_bottom_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(chany_top_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output58 (.I(net58),
    .Z(chany_top_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output59 (.I(net59),
    .Z(chany_top_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output60 (.I(net60),
    .Z(chany_top_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output61 (.I(net61),
    .Z(chany_top_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output62 (.I(net62),
    .Z(chany_top_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output63 (.I(net63),
    .Z(chany_top_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(chany_top_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output65 (.I(net65),
    .Z(chany_top_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output66 (.I(net66),
    .Z(chany_top_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output67 (.I(net67),
    .Z(chany_top_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(chany_top_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output69 (.I(net69),
    .Z(chany_top_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output70 (.I(net70),
    .Z(chany_top_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output71 (.I(net71),
    .Z(chany_top_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_0__1__97 (.ZN(net97));
 assign chanx_right_out[0] = net97;
 assign chanx_right_out[10] = net87;
 assign chanx_right_out[11] = net86;
 assign chanx_right_out[12] = net85;
 assign chanx_right_out[13] = net84;
 assign chanx_right_out[14] = net83;
 assign chanx_right_out[19] = net82;
 assign chanx_right_out[1] = net96;
 assign chanx_right_out[2] = net95;
 assign chanx_right_out[3] = net94;
 assign chanx_right_out[4] = net93;
 assign chanx_right_out[5] = net92;
 assign chanx_right_out[6] = net91;
 assign chanx_right_out[7] = net90;
 assign chanx_right_out[8] = net89;
 assign chanx_right_out[9] = net88;
 assign chany_bottom_out[0] = net81;
 assign chany_bottom_out[12] = net78;
 assign chany_bottom_out[16] = net77;
 assign chany_bottom_out[4] = net80;
 assign chany_bottom_out[8] = net79;
 assign chany_top_out[0] = net76;
 assign chany_top_out[12] = net73;
 assign chany_top_out[16] = net72;
 assign chany_top_out[4] = net75;
 assign chany_top_out[8] = net74;
endmodule

