// This is the unpowered netlist.
module sb_2__1_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
    ccff_head,
    ccff_tail,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    pReset,
    prog_clk,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
    chanx_left_in,
    chanx_left_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
 input ccff_head;
 output ccff_tail;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input pReset;
 input prog_clk;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
 input [19:0] chanx_left_in;
 output [19:0] chanx_left_out;
 input [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;
 input [19:0] chany_top_in;
 output [19:0] chany_top_out;

 wire net97;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net81;
 wire net78;
 wire net77;
 wire net80;
 wire net79;
 wire net76;
 wire net73;
 wire net72;
 wire net75;
 wire net74;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire clknet_0_prog_clk;
 wire clknet_3_0__leaf_prog_clk;
 wire clknet_3_1__leaf_prog_clk;
 wire clknet_3_2__leaf_prog_clk;
 wire clknet_3_3__leaf_prog_clk;
 wire clknet_3_4__leaf_prog_clk;
 wire clknet_3_5__leaf_prog_clk;
 wire clknet_3_6__leaf_prog_clk;
 wire clknet_3_7__leaf_prog_clk;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_1.DFFR_2_.Q ;
 wire \mem_bottom_track_1.DFFR_3_.Q ;
 wire \mem_bottom_track_1.DFFR_4_.Q ;
 wire \mem_bottom_track_1.DFFR_5_.Q ;
 wire \mem_bottom_track_1.DFFR_6_.Q ;
 wire \mem_bottom_track_1.DFFR_7_.Q ;
 wire \mem_bottom_track_17.DFFR_0_.D ;
 wire \mem_bottom_track_17.DFFR_0_.Q ;
 wire \mem_bottom_track_17.DFFR_1_.Q ;
 wire \mem_bottom_track_17.DFFR_2_.Q ;
 wire \mem_bottom_track_17.DFFR_3_.Q ;
 wire \mem_bottom_track_17.DFFR_4_.Q ;
 wire \mem_bottom_track_17.DFFR_5_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_2_.Q ;
 wire \mem_bottom_track_25.DFFR_3_.Q ;
 wire \mem_bottom_track_25.DFFR_4_.Q ;
 wire \mem_bottom_track_25.DFFR_5_.Q ;
 wire \mem_bottom_track_33.DFFR_0_.Q ;
 wire \mem_bottom_track_33.DFFR_1_.Q ;
 wire \mem_bottom_track_33.DFFR_2_.Q ;
 wire \mem_bottom_track_33.DFFR_3_.Q ;
 wire \mem_bottom_track_33.DFFR_4_.Q ;
 wire \mem_bottom_track_33.DFFR_5_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_bottom_track_9.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_2_.Q ;
 wire \mem_bottom_track_9.DFFR_3_.Q ;
 wire \mem_bottom_track_9.DFFR_4_.Q ;
 wire \mem_left_track_1.DFFR_0_.Q ;
 wire \mem_left_track_1.DFFR_1_.Q ;
 wire \mem_left_track_1.DFFR_2_.Q ;
 wire \mem_left_track_1.DFFR_3_.Q ;
 wire \mem_left_track_1.DFFR_4_.Q ;
 wire \mem_left_track_1.DFFR_5_.Q ;
 wire \mem_left_track_11.DFFR_0_.D ;
 wire \mem_left_track_11.DFFR_0_.Q ;
 wire \mem_left_track_11.DFFR_1_.Q ;
 wire \mem_left_track_13.DFFR_0_.Q ;
 wire \mem_left_track_13.DFFR_1_.Q ;
 wire \mem_left_track_15.DFFR_0_.Q ;
 wire \mem_left_track_15.DFFR_1_.Q ;
 wire \mem_left_track_17.DFFR_0_.Q ;
 wire \mem_left_track_17.DFFR_1_.Q ;
 wire \mem_left_track_19.DFFR_0_.Q ;
 wire \mem_left_track_19.DFFR_1_.Q ;
 wire \mem_left_track_21.DFFR_0_.Q ;
 wire \mem_left_track_21.DFFR_1_.Q ;
 wire \mem_left_track_23.DFFR_0_.Q ;
 wire \mem_left_track_23.DFFR_1_.Q ;
 wire \mem_left_track_25.DFFR_0_.Q ;
 wire \mem_left_track_25.DFFR_1_.Q ;
 wire \mem_left_track_27.DFFR_0_.Q ;
 wire \mem_left_track_27.DFFR_1_.Q ;
 wire \mem_left_track_29.DFFR_0_.Q ;
 wire \mem_left_track_3.DFFR_0_.Q ;
 wire \mem_left_track_3.DFFR_1_.Q ;
 wire \mem_left_track_3.DFFR_2_.Q ;
 wire \mem_left_track_3.DFFR_3_.Q ;
 wire \mem_left_track_3.DFFR_4_.Q ;
 wire \mem_left_track_3.DFFR_5_.Q ;
 wire \mem_left_track_5.DFFR_0_.Q ;
 wire \mem_left_track_5.DFFR_1_.Q ;
 wire \mem_left_track_5.DFFR_2_.Q ;
 wire \mem_left_track_5.DFFR_3_.Q ;
 wire \mem_left_track_5.DFFR_4_.Q ;
 wire \mem_left_track_5.DFFR_5_.Q ;
 wire \mem_left_track_7.DFFR_0_.Q ;
 wire \mem_left_track_7.DFFR_1_.Q ;
 wire \mem_left_track_7.DFFR_2_.Q ;
 wire \mem_left_track_7.DFFR_3_.Q ;
 wire \mem_left_track_7.DFFR_4_.Q ;
 wire \mem_left_track_7.DFFR_5_.Q ;
 wire \mem_left_track_9.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_0.DFFR_2_.Q ;
 wire \mem_top_track_0.DFFR_3_.Q ;
 wire \mem_top_track_0.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_5_.Q ;
 wire \mem_top_track_0.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_7_.Q ;
 wire \mem_top_track_16.DFFR_0_.D ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_2_.Q ;
 wire \mem_top_track_16.DFFR_3_.Q ;
 wire \mem_top_track_16.DFFR_4_.Q ;
 wire \mem_top_track_16.DFFR_5_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_2_.Q ;
 wire \mem_top_track_24.DFFR_3_.Q ;
 wire \mem_top_track_24.DFFR_4_.Q ;
 wire \mem_top_track_24.DFFR_5_.Q ;
 wire \mem_top_track_32.DFFR_0_.Q ;
 wire \mem_top_track_32.DFFR_1_.Q ;
 wire \mem_top_track_32.DFFR_2_.Q ;
 wire \mem_top_track_32.DFFR_3_.Q ;
 wire \mem_top_track_32.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire \mem_top_track_8.DFFR_1_.Q ;
 wire \mem_top_track_8.DFFR_2_.Q ;
 wire \mem_top_track_8.DFFR_3_.Q ;
 wire \mem_top_track_8.DFFR_4_.Q ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net8;
 wire net9;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__244__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__CLK (.I(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__CLK (.I(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_prog_clk_I (.I(prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_prog_clk_I (.I(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(chany_bottom_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(chany_bottom_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(chany_bottom_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(chany_bottom_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(chany_bottom_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(chany_bottom_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(chany_bottom_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(chany_top_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(chany_top_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(chany_top_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ccff_head));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(chany_top_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(chany_top_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(chany_top_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(chany_top_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(chany_top_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(chany_top_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(chany_top_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(chany_top_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(chany_top_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(chany_top_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(chany_bottom_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(chany_top_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(chany_top_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(chany_top_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(chany_top_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(chany_top_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(chany_top_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(pReset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(chany_bottom_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(chany_bottom_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(chany_bottom_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(chany_bottom_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(chany_bottom_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(chany_bottom_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(chany_bottom_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_134 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _122_ (.I(net36),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _123_ (.I(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _124_ (.I(_111_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _125_ (.I(_111_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _126_ (.I(_111_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _127_ (.I(_111_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _128_ (.I(_111_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _129_ (.I(_111_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _130_ (.I(_111_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _131_ (.I(_111_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _132_ (.I(_111_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _133_ (.I(_111_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _134_ (.I(_110_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _135_ (.I(_112_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _136_ (.I(_112_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _137_ (.I(_112_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _138_ (.I(_112_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _139_ (.I(_112_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _140_ (.I(_112_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _141_ (.I(_112_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _142_ (.I(_112_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _143_ (.I(_112_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _144_ (.I(_112_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _145_ (.I(_110_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _146_ (.I(_113_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _147_ (.I(_113_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _148_ (.I(_113_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _149_ (.I(_113_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _150_ (.I(_113_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _151_ (.I(_113_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _152_ (.I(_113_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _153_ (.I(_113_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _154_ (.I(_113_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _155_ (.I(_113_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _156_ (.I(_110_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _157_ (.I(_114_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _158_ (.I(_114_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _159_ (.I(_114_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _160_ (.I(_114_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _161_ (.I(_114_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _162_ (.I(_114_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _163_ (.I(_114_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _164_ (.I(_114_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _165_ (.I(_114_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _166_ (.I(_114_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _167_ (.I(_110_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _168_ (.I(_115_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _169_ (.I(_115_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _170_ (.I(_115_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _171_ (.I(_115_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _172_ (.I(_115_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _173_ (.I(_115_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _174_ (.I(_115_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _175_ (.I(_115_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _176_ (.I(_115_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _177_ (.I(_115_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _178_ (.I(_110_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _179_ (.I(_116_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _180_ (.I(_116_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _181_ (.I(_116_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _182_ (.I(_116_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _183_ (.I(_116_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _184_ (.I(_116_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _185_ (.I(_116_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _186_ (.I(_116_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _187_ (.I(_116_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _188_ (.I(_116_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _189_ (.I(_110_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _190_ (.I(_117_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _191_ (.I(_117_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _192_ (.I(_117_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _193_ (.I(_117_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _194_ (.I(_117_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _195_ (.I(_117_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _196_ (.I(_117_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _197_ (.I(_117_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _198_ (.I(_117_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _199_ (.I(_117_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _200_ (.I(_110_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _201_ (.I(_118_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _202_ (.I(_118_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _203_ (.I(_118_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _204_ (.I(_118_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _205_ (.I(_118_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _206_ (.I(_118_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _207_ (.I(_118_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _208_ (.I(_118_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _209_ (.I(_118_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _210_ (.I(_118_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _211_ (.I(_110_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _212_ (.I(_119_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _213_ (.I(_119_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _214_ (.I(_119_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _215_ (.I(_119_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _216_ (.I(_119_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _217_ (.I(_119_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _218_ (.I(_119_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _219_ (.I(_119_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _220_ (.I(_119_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _221_ (.I(_119_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _222_ (.I(_110_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _223_ (.I(_120_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _224_ (.I(_120_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _225_ (.I(_120_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _226_ (.I(_120_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _227_ (.I(_120_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _228_ (.I(_120_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _229_ (.I(_120_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _230_ (.I(_120_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _231_ (.I(_120_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _232_ (.I(_120_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _233_ (.I(net36),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _234_ (.I(_121_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _235_ (.I(_121_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _236_ (.I(_121_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _237_ (.I(_121_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _238_ (.I(_121_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _239_ (.I(_121_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _240_ (.I(_121_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _241_ (.I(_121_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _242_ (.I(_121_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _243_ (.I(_121_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _244_ (.D(net135),
    .RN(_000_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _245_ (.D(net183),
    .RN(_001_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _246_ (.D(net168),
    .RN(_002_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _247_ (.D(net154),
    .RN(_003_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _248_ (.D(net201),
    .RN(_004_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _249_ (.D(net206),
    .RN(_005_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _250_ (.D(net203),
    .RN(_006_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _251_ (.D(net1),
    .RN(_007_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _252_ (.D(net193),
    .RN(_008_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_7_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _253_ (.D(net202),
    .RN(_009_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_6_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _254_ (.D(net113),
    .RN(_010_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _255_ (.D(net102),
    .RN(_011_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _256_ (.D(net121),
    .RN(_012_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _257_ (.D(net171),
    .RN(_013_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _258_ (.D(net104),
    .RN(_014_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _259_ (.D(net200),
    .RN(_015_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _260_ (.D(net133),
    .RN(_016_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _261_ (.D(net147),
    .RN(_017_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _262_ (.D(net141),
    .RN(_018_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _263_ (.D(net117),
    .RN(_019_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _264_ (.D(net173),
    .RN(_020_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _265_ (.D(net122),
    .RN(_021_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _266_ (.D(net164),
    .RN(_022_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _267_ (.D(net100),
    .RN(_023_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _268_ (.D(net114),
    .RN(_024_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _269_ (.D(net132),
    .RN(_025_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _270_ (.D(net185),
    .RN(_026_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _271_ (.D(net161),
    .RN(_027_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _272_ (.D(net160),
    .RN(_028_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _273_ (.D(net134),
    .RN(_029_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _274_ (.D(net172),
    .RN(_030_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _275_ (.D(net149),
    .RN(_031_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _276_ (.D(net145),
    .RN(_032_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _277_ (.D(net118),
    .RN(_033_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _278_ (.D(net159),
    .RN(_034_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _279_ (.D(net152),
    .RN(_035_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _280_ (.D(net123),
    .RN(_036_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _281_ (.D(net105),
    .RN(_037_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _282_ (.D(net103),
    .RN(_038_),
    .CLK(clknet_3_1__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _283_ (.D(net116),
    .RN(_039_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_top_track_32.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _284_ (.D(net175),
    .RN(_040_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _285_ (.D(net125),
    .RN(_041_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _286_ (.D(net156),
    .RN(_042_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _287_ (.D(net111),
    .RN(_043_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _288_ (.D(net177),
    .RN(_044_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _289_ (.D(net142),
    .RN(_045_),
    .CLK(clknet_3_0__leaf_prog_clk),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _290_ (.D(net169),
    .RN(_046_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _291_ (.D(net195),
    .RN(_047_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _292_ (.D(net199),
    .RN(_048_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _293_ (.D(net119),
    .RN(_049_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _294_ (.D(net109),
    .RN(_050_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _295_ (.D(net140),
    .RN(_051_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_17.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _296_ (.D(net184),
    .RN(_052_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _297_ (.D(net110),
    .RN(_053_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _298_ (.D(net189),
    .RN(_054_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _299_ (.D(net131),
    .RN(_055_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _300_ (.D(net137),
    .RN(_056_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _301_ (.D(net128),
    .RN(_057_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _302_ (.D(net107),
    .RN(_058_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _303_ (.D(net124),
    .RN(_059_),
    .CLK(clknet_3_2__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _304_ (.D(net115),
    .RN(_060_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _305_ (.D(net180),
    .RN(_061_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _306_ (.D(net194),
    .RN(_062_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _307_ (.D(net143),
    .RN(_063_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_bottom_track_33.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _308_ (.D(net120),
    .RN(_064_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _309_ (.D(net158),
    .RN(_065_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _310_ (.D(net153),
    .RN(_066_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _311_ (.D(net181),
    .RN(_067_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _312_ (.D(net151),
    .RN(_068_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _313_ (.D(net192),
    .RN(_069_),
    .CLK(clknet_3_3__leaf_prog_clk),
    .Q(\mem_left_track_1.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _314_ (.D(net196),
    .RN(_070_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_3.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _315_ (.D(net182),
    .RN(_071_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_3.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _316_ (.D(net144),
    .RN(_072_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_3.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _317_ (.D(net188),
    .RN(_073_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_3.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _318_ (.D(net174),
    .RN(_074_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_3.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _319_ (.D(net139),
    .RN(_075_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_3.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _320_ (.D(net178),
    .RN(_076_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_5.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _321_ (.D(net130),
    .RN(_077_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_5.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _322_ (.D(net165),
    .RN(_078_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_5.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _323_ (.D(net127),
    .RN(_079_),
    .CLK(clknet_3_6__leaf_prog_clk),
    .Q(\mem_left_track_5.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _324_ (.D(net155),
    .RN(_080_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_5.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _325_ (.D(net106),
    .RN(_081_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_5.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _326_ (.D(net162),
    .RN(_082_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_7.DFFR_5_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _327_ (.D(net163),
    .RN(_083_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_7.DFFR_4_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _328_ (.D(net146),
    .RN(_084_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_7.DFFR_3_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _329_ (.D(net138),
    .RN(_085_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_7.DFFR_2_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _330_ (.D(net179),
    .RN(_086_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_7.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _331_ (.D(net108),
    .RN(_087_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_7.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _332_ (.D(net157),
    .RN(_088_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_11.DFFR_0_.D ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _333_ (.D(net197),
    .RN(_089_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_9.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _334_ (.D(net112),
    .RN(_090_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_left_track_11.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _335_ (.D(net167),
    .RN(_091_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_11.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _336_ (.D(net98),
    .RN(_092_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_21.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _337_ (.D(net204),
    .RN(_093_),
    .CLK(clknet_3_4__leaf_prog_clk),
    .Q(\mem_left_track_21.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _338_ (.D(net187),
    .RN(_094_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_23.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _339_ (.D(net150),
    .RN(_095_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_23.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _340_ (.D(net190),
    .RN(_096_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _341_ (.D(net136),
    .RN(_097_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_25.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _342_ (.D(net99),
    .RN(_098_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_27.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _343_ (.D(net126),
    .RN(_099_),
    .CLK(clknet_3_7__leaf_prog_clk),
    .Q(\mem_left_track_27.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _344_ (.D(net186),
    .RN(_100_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_13.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _345_ (.D(net101),
    .RN(_101_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_13.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _346_ (.D(net191),
    .RN(_102_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_15.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _347_ (.D(net148),
    .RN(_103_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_15.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _348_ (.D(net176),
    .RN(_104_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _349_ (.D(net129),
    .RN(_105_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_17.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _350_ (.D(net166),
    .RN(_106_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_19.DFFR_1_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _351_ (.D(net205),
    .RN(_107_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_19.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _352_ (.D(net170),
    .RN(_108_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _353_ (.D(net198),
    .RN(_109_),
    .CLK(clknet_3_5__leaf_prog_clk),
    .Q(\mem_left_track_29.DFFR_0_.Q ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _380_ (.I(net33),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _381_ (.I(net19),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _382_ (.I(net23),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _383_ (.I(net27),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _384_ (.I(net26),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _385_ (.I(net25),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _386_ (.I(net24),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _387_ (.I(net22),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _388_ (.I(net21),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _389_ (.I(net20),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _390_ (.I(net18),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _391_ (.I(net35),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _392_ (.I(net34),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _393_ (.I(net32),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _394_ (.I(net31),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _395_ (.I(net30),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _396_ (.I(net29),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _397_ (.I(net28),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _398_ (.I(net17),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _399_ (.I(net9),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _400_ (.I(net8),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _401_ (.I(net7),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _402_ (.I(net6),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _403_ (.I(net5),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _404_ (.I(net4),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _405_ (.I(net3),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _406_ (.I(net16),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _407_ (.I(net15),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _408_ (.I(net14),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _409_ (.I(net13),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _410_ (.I(net12),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _411_ (.I(net11),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _412_ (.I(net10),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _413_ (.I(net2),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_prog_clk (.I(prog_clk),
    .Z(clknet_0_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_0__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_1__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_2__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_3__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_4__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_5__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_6__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_prog_clk (.I(clknet_0_prog_clk),
    .Z(clknet_3_7__leaf_prog_clk));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(\mem_left_track_21.DFFR_0_.Q ),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\mem_bottom_track_33.DFFR_4_.Q ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(\mem_left_track_7.DFFR_5_.Q ),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(\mem_left_track_27.DFFR_1_.Q ),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(\mem_bottom_track_17.DFFR_2_.Q ),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(\mem_bottom_track_1.DFFR_0_.D ),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(\mem_top_track_0.DFFR_2_.Q ),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(\mem_bottom_track_1.DFFR_5_.Q ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(\mem_top_track_0.DFFR_0_.Q ),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(\mem_left_track_19.DFFR_1_.Q ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold108 (.I(\mem_left_track_17.DFFR_1_.Q ),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(\mem_top_track_0.DFFR_1_.Q ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\mem_left_track_5.DFFR_5_.Q ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\mem_bottom_track_17.DFFR_0_.Q ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\mem_bottom_track_25.DFFR_3_.Q ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\mem_bottom_track_9.DFFR_1_.Q ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\mem_left_track_11.DFFR_0_.Q ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\mem_bottom_track_1.DFFR_4_.Q ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\mem_top_track_16.DFFR_2_.Q ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\mem_bottom_track_33.DFFR_2_.Q ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\mem_top_track_24.DFFR_5_.Q ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\mem_left_track_27.DFFR_0_.Q ),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\mem_top_track_8.DFFR_1_.Q ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\mem_top_track_16.DFFR_5_.Q ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\mem_bottom_track_17.DFFR_1_.Q ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\mem_left_track_1.DFFR_4_.Q ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\mem_bottom_track_1.DFFR_2_.Q ),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\mem_top_track_0.DFFR_7_.Q ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\mem_top_track_32.DFFR_2_.Q ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\mem_bottom_track_33.DFFR_3_.Q ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\mem_bottom_track_9.DFFR_3_.Q ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\mem_left_track_25.DFFR_1_.Q ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\mem_top_track_16.DFFR_3_.Q ),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\mem_left_track_5.DFFR_1_.Q ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\mem_bottom_track_17.DFFR_5_.Q ),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\mem_left_track_15.DFFR_1_.Q ),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\mem_left_track_5.DFFR_3_.Q ),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\mem_bottom_track_25.DFFR_1_.Q ),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\mem_top_track_16.DFFR_1_.Q ),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\mem_top_track_8.DFFR_4_.Q ),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\mem_top_track_24.DFFR_3_.Q ),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\mem_top_track_0.DFFR_6_.Q ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\mem_left_track_23.DFFR_1_.Q ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\mem_left_track_11.DFFR_1_.Q ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\mem_bottom_track_25.DFFR_0_.Q ),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\mem_left_track_7.DFFR_1_.Q ),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\mem_left_track_1.DFFR_5_.Q ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\mem_bottom_track_17.DFFR_0_.D ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\mem_top_track_8.DFFR_2_.Q ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\mem_bottom_track_1.DFFR_7_.Q ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\mem_bottom_track_25.DFFR_5_.Q ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\mem_left_track_3.DFFR_2_.Q ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(\mem_top_track_24.DFFR_0_.Q ),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\mem_left_track_7.DFFR_2_.Q ),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\mem_bottom_track_1.DFFR_3_.Q ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(\mem_top_track_8.DFFR_3_.Q ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\mem_left_track_13.DFFR_1_.Q ),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(\mem_top_track_24.DFFR_1_.Q ),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\mem_left_track_21.DFFR_1_.Q ),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(\mem_left_track_1.DFFR_0_.Q ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\mem_top_track_32.DFFR_3_.Q ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(\mem_left_track_1.DFFR_2_.Q ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\mem_top_track_0.DFFR_3_.Q ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(\mem_left_track_5.DFFR_0_.Q ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\mem_bottom_track_9.DFFR_2_.Q ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\mem_top_track_32.DFFR_0_.Q ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(\mem_left_track_9.DFFR_0_.Q ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\mem_left_track_1.DFFR_3_.Q ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(\mem_top_track_32.DFFR_4_.Q ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\mem_top_track_24.DFFR_4_.Q ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(\mem_top_track_16.DFFR_0_.D ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\mem_left_track_7.DFFR_4_.Q ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(\mem_left_track_7.DFFR_3_.Q ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\mem_top_track_16.DFFR_4_.Q ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(\mem_left_track_5.DFFR_2_.Q ),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\mem_left_track_19.DFFR_0_.Q ),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\mem_bottom_track_1.DFFR_0_.Q ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(\mem_left_track_11.DFFR_0_.D ),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\mem_top_track_0.DFFR_4_.Q ),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(\mem_bottom_track_17.DFFR_4_.Q ),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\mem_left_track_29.DFFR_0_.Q ),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(\mem_bottom_track_1.DFFR_1_.Q ),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\mem_top_track_24.DFFR_2_.Q ),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(\mem_top_track_8.DFFR_0_.Q ),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\mem_left_track_3.DFFR_0_.Q ),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(\mem_bottom_track_9.DFFR_4_.Q ),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\mem_left_track_17.DFFR_0_.Q ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\mem_top_track_32.DFFR_1_.Q ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(\mem_bottom_track_9.DFFR_0_.Q ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\mem_left_track_5.DFFR_4_.Q ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(\mem_left_track_7.DFFR_0_.Q ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\mem_bottom_track_33.DFFR_1_.Q ),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(\mem_left_track_1.DFFR_1_.Q ),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\mem_left_track_3.DFFR_3_.Q ),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(\mem_top_track_0.DFFR_5_.Q ),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\mem_bottom_track_25.DFFR_4_.Q ),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(\mem_top_track_16.DFFR_0_.Q ),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\mem_left_track_13.DFFR_0_.Q ),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\mem_left_track_3.DFFR_5_.Q ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(\mem_left_track_23.DFFR_0_.Q ),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\mem_left_track_3.DFFR_1_.Q ),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(\mem_bottom_track_25.DFFR_2_.Q ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\mem_left_track_25.DFFR_0_.Q ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(\mem_left_track_15.DFFR_0_.Q ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(\mem_bottom_track_33.DFFR_5_.Q ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(\mem_bottom_track_1.DFFR_6_.Q ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(\mem_bottom_track_33.DFFR_0_.Q ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(\mem_bottom_track_17.DFFR_3_.Q ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(\mem_left_track_3.DFFR_4_.Q ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ccff_head),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(chany_bottom_in[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(chany_bottom_in[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(chany_bottom_in[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(chany_bottom_in[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(chany_bottom_in[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(chany_bottom_in[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(chany_bottom_in[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(chany_top_in[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(chany_top_in[10]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(chany_top_in[11]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(chany_bottom_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(chany_top_in[12]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(chany_top_in[13]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(chany_top_in[14]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(chany_top_in[15]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(chany_top_in[16]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(chany_top_in[17]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(chany_top_in[18]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(chany_top_in[19]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(chany_top_in[1]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(chany_top_in[2]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(chany_bottom_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(chany_top_in[4]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(chany_top_in[5]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(chany_top_in[6]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(chany_top_in[7]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(chany_top_in[8]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(chany_top_in[9]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(pReset),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(chany_bottom_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(chany_bottom_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(chany_bottom_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(chany_bottom_in[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(chany_bottom_in[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(chany_bottom_in[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(ccff_tail));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(chanx_left_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(chanx_left_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output40 (.I(net40),
    .Z(chanx_left_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output41 (.I(net41),
    .Z(chanx_left_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output42 (.I(net42),
    .Z(chany_bottom_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output43 (.I(net43),
    .Z(chany_bottom_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output44 (.I(net44),
    .Z(chany_bottom_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output45 (.I(net45),
    .Z(chany_bottom_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output46 (.I(net46),
    .Z(chany_bottom_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output47 (.I(net47),
    .Z(chany_bottom_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output48 (.I(net48),
    .Z(chany_bottom_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(chany_bottom_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output50 (.I(net50),
    .Z(chany_bottom_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output51 (.I(net51),
    .Z(chany_bottom_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output52 (.I(net52),
    .Z(chany_bottom_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output53 (.I(net53),
    .Z(chany_bottom_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output54 (.I(net54),
    .Z(chany_bottom_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output55 (.I(net55),
    .Z(chany_bottom_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output56 (.I(net56),
    .Z(chany_bottom_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output57 (.I(net57),
    .Z(chany_top_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output58 (.I(net58),
    .Z(chany_top_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output59 (.I(net59),
    .Z(chany_top_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(chany_top_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output61 (.I(net61),
    .Z(chany_top_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output62 (.I(net62),
    .Z(chany_top_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output63 (.I(net63),
    .Z(chany_top_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output64 (.I(net64),
    .Z(chany_top_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output65 (.I(net65),
    .Z(chany_top_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output66 (.I(net66),
    .Z(chany_top_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output67 (.I(net67),
    .Z(chany_top_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(chany_top_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output69 (.I(net69),
    .Z(chany_top_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output70 (.I(net70),
    .Z(chany_top_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output71 (.I(net71),
    .Z(chany_top_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel sb_2__1__97 (.ZN(net97));
 assign chanx_left_out[0] = net97;
 assign chanx_left_out[10] = net87;
 assign chanx_left_out[11] = net86;
 assign chanx_left_out[12] = net85;
 assign chanx_left_out[13] = net84;
 assign chanx_left_out[14] = net83;
 assign chanx_left_out[15] = net82;
 assign chanx_left_out[1] = net96;
 assign chanx_left_out[2] = net95;
 assign chanx_left_out[3] = net94;
 assign chanx_left_out[4] = net93;
 assign chanx_left_out[5] = net92;
 assign chanx_left_out[6] = net91;
 assign chanx_left_out[7] = net90;
 assign chanx_left_out[8] = net89;
 assign chanx_left_out[9] = net88;
 assign chany_bottom_out[0] = net81;
 assign chany_bottom_out[12] = net78;
 assign chany_bottom_out[16] = net77;
 assign chany_bottom_out[4] = net80;
 assign chany_bottom_out[8] = net79;
 assign chany_top_out[0] = net76;
 assign chany_top_out[12] = net73;
 assign chany_top_out[16] = net72;
 assign chany_top_out[4] = net75;
 assign chany_top_out[8] = net74;
endmodule

