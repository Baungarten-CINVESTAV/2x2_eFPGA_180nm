magic
tech gf180mcuD
magscale 1 10
timestamp 1702149352
<< metal1 >>
rect 10098 41806 10110 41858
rect 10162 41855 10174 41858
rect 11218 41855 11230 41858
rect 10162 41809 11230 41855
rect 10162 41806 10174 41809
rect 11218 41806 11230 41809
rect 11282 41806 11294 41858
rect 15474 41246 15486 41298
rect 15538 41295 15550 41298
rect 16034 41295 16046 41298
rect 15538 41249 16046 41295
rect 15538 41246 15550 41249
rect 16034 41246 16046 41249
rect 16098 41246 16110 41298
rect 5394 41022 5406 41074
rect 5458 41071 5470 41074
rect 5954 41071 5966 41074
rect 5458 41025 5966 41071
rect 5458 41022 5470 41025
rect 5954 41022 5966 41025
rect 6018 41022 6030 41074
rect 22194 41022 22206 41074
rect 22258 41071 22270 41074
rect 23314 41071 23326 41074
rect 22258 41025 23326 41071
rect 22258 41022 22270 41025
rect 23314 41022 23326 41025
rect 23378 41022 23390 41074
rect 20178 40910 20190 40962
rect 20242 40959 20254 40962
rect 20850 40959 20862 40962
rect 20242 40913 20862 40959
rect 20242 40910 20254 40913
rect 20850 40910 20862 40913
rect 20914 40910 20926 40962
rect 1344 40794 42560 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 42560 40794
rect 1344 40708 42560 40742
rect 1822 40626 1874 40638
rect 1822 40562 1874 40574
rect 11902 40626 11954 40638
rect 11902 40562 11954 40574
rect 12350 40626 12402 40638
rect 12350 40562 12402 40574
rect 13134 40626 13186 40638
rect 13134 40562 13186 40574
rect 13694 40626 13746 40638
rect 13694 40562 13746 40574
rect 14254 40626 14306 40638
rect 14254 40562 14306 40574
rect 14814 40626 14866 40638
rect 14814 40562 14866 40574
rect 17726 40626 17778 40638
rect 17726 40562 17778 40574
rect 19182 40626 19234 40638
rect 19182 40562 19234 40574
rect 19854 40626 19906 40638
rect 19854 40562 19906 40574
rect 20190 40626 20242 40638
rect 20190 40562 20242 40574
rect 9326 40514 9378 40526
rect 17054 40514 17106 40526
rect 4050 40462 4062 40514
rect 4114 40462 4126 40514
rect 5954 40462 5966 40514
rect 6018 40462 6030 40514
rect 7858 40462 7870 40514
rect 7922 40462 7934 40514
rect 11218 40462 11230 40514
rect 11282 40462 11294 40514
rect 16034 40462 16046 40514
rect 16098 40462 16110 40514
rect 9326 40450 9378 40462
rect 17054 40450 17106 40462
rect 20750 40514 20802 40526
rect 20750 40450 20802 40462
rect 21758 40514 21810 40526
rect 23314 40462 23326 40514
rect 23378 40462 23390 40514
rect 21758 40450 21810 40462
rect 24558 40402 24610 40414
rect 3266 40350 3278 40402
rect 3330 40350 3342 40402
rect 4946 40350 4958 40402
rect 5010 40350 5022 40402
rect 6626 40350 6638 40402
rect 6690 40350 6702 40402
rect 8754 40350 8766 40402
rect 8818 40350 8830 40402
rect 9538 40350 9550 40402
rect 9602 40350 9614 40402
rect 10322 40350 10334 40402
rect 10386 40350 10398 40402
rect 15138 40350 15150 40402
rect 15202 40350 15214 40402
rect 17266 40350 17278 40402
rect 17330 40350 17342 40402
rect 18498 40350 18510 40402
rect 18562 40350 18574 40402
rect 20962 40350 20974 40402
rect 21026 40350 21038 40402
rect 21970 40350 21982 40402
rect 22034 40350 22046 40402
rect 22418 40350 22430 40402
rect 22482 40350 22494 40402
rect 24558 40338 24610 40350
rect 25790 40402 25842 40414
rect 25790 40338 25842 40350
rect 26126 40402 26178 40414
rect 26126 40338 26178 40350
rect 2706 40238 2718 40290
rect 2770 40238 2782 40290
rect 24994 40238 25006 40290
rect 25058 40238 25070 40290
rect 26562 40238 26574 40290
rect 26626 40238 26638 40290
rect 1344 40010 42560 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 42560 40010
rect 1344 39924 42560 39958
rect 2494 39842 2546 39854
rect 2494 39778 2546 39790
rect 4062 39842 4114 39854
rect 4062 39778 4114 39790
rect 10222 39730 10274 39742
rect 17614 39730 17666 39742
rect 9426 39678 9438 39730
rect 9490 39678 9502 39730
rect 16818 39678 16830 39730
rect 16882 39678 16894 39730
rect 10222 39666 10274 39678
rect 17614 39666 17666 39678
rect 18846 39730 18898 39742
rect 18846 39666 18898 39678
rect 21534 39730 21586 39742
rect 21534 39666 21586 39678
rect 22878 39730 22930 39742
rect 22878 39666 22930 39678
rect 25566 39730 25618 39742
rect 27570 39678 27582 39730
rect 27634 39678 27646 39730
rect 25566 39666 25618 39678
rect 6974 39618 7026 39630
rect 7858 39566 7870 39618
rect 7922 39566 7934 39618
rect 8418 39566 8430 39618
rect 8482 39566 8494 39618
rect 19282 39566 19294 39618
rect 19346 39566 19358 39618
rect 23986 39566 23998 39618
rect 24050 39566 24062 39618
rect 26002 39566 26014 39618
rect 26066 39566 26078 39618
rect 26674 39566 26686 39618
rect 26738 39566 26750 39618
rect 6974 39554 7026 39566
rect 5630 39506 5682 39518
rect 5630 39442 5682 39454
rect 5966 39506 6018 39518
rect 5966 39442 6018 39454
rect 6638 39506 6690 39518
rect 6638 39442 6690 39454
rect 10558 39506 10610 39518
rect 10558 39442 10610 39454
rect 11006 39506 11058 39518
rect 11006 39442 11058 39454
rect 20414 39506 20466 39518
rect 20414 39442 20466 39454
rect 23102 39506 23154 39518
rect 23102 39442 23154 39454
rect 3278 39394 3330 39406
rect 3278 39330 3330 39342
rect 4846 39394 4898 39406
rect 4846 39330 4898 39342
rect 6302 39394 6354 39406
rect 6302 39330 6354 39342
rect 7310 39394 7362 39406
rect 7310 39330 7362 39342
rect 7646 39394 7698 39406
rect 7646 39330 7698 39342
rect 8654 39394 8706 39406
rect 8654 39330 8706 39342
rect 8990 39394 9042 39406
rect 8990 39330 9042 39342
rect 16382 39394 16434 39406
rect 16382 39330 16434 39342
rect 19070 39394 19122 39406
rect 19070 39330 19122 39342
rect 23774 39394 23826 39406
rect 23774 39330 23826 39342
rect 25790 39394 25842 39406
rect 25790 39330 25842 39342
rect 26462 39394 26514 39406
rect 26462 39330 26514 39342
rect 27134 39394 27186 39406
rect 27134 39330 27186 39342
rect 1344 39226 42560 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 42560 39226
rect 1344 39140 42560 39174
rect 2158 39058 2210 39070
rect 2158 38994 2210 39006
rect 3726 39058 3778 39070
rect 3726 38994 3778 39006
rect 5518 39058 5570 39070
rect 5518 38994 5570 39006
rect 6862 39058 6914 39070
rect 6862 38994 6914 39006
rect 7534 39058 7586 39070
rect 7534 38994 7586 39006
rect 8654 39058 8706 39070
rect 8654 38994 8706 39006
rect 9662 39058 9714 39070
rect 9662 38994 9714 39006
rect 26238 39058 26290 39070
rect 26238 38994 26290 39006
rect 2942 38946 2994 38958
rect 2942 38882 2994 38894
rect 4846 38946 4898 38958
rect 4846 38882 4898 38894
rect 6190 38946 6242 38958
rect 6190 38882 6242 38894
rect 8318 38946 8370 38958
rect 8318 38882 8370 38894
rect 6526 38834 6578 38846
rect 4386 38782 4398 38834
rect 4450 38782 4462 38834
rect 5058 38782 5070 38834
rect 5122 38782 5134 38834
rect 5730 38782 5742 38834
rect 5794 38782 5806 38834
rect 6526 38770 6578 38782
rect 7198 38834 7250 38846
rect 8082 38782 8094 38834
rect 8146 38782 8158 38834
rect 8866 38782 8878 38834
rect 8930 38782 8942 38834
rect 7198 38770 7250 38782
rect 1822 38722 1874 38734
rect 1822 38658 1874 38670
rect 10222 38722 10274 38734
rect 10222 38658 10274 38670
rect 26798 38722 26850 38734
rect 26798 38658 26850 38670
rect 1344 38442 42560 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 42560 38442
rect 1344 38356 42560 38390
rect 2158 38274 2210 38286
rect 2158 38210 2210 38222
rect 8318 38050 8370 38062
rect 10670 38050 10722 38062
rect 7074 37998 7086 38050
rect 7138 37998 7150 38050
rect 9090 37998 9102 38050
rect 9154 37998 9166 38050
rect 9762 37998 9774 38050
rect 9826 37998 9838 38050
rect 8318 37986 8370 37998
rect 10670 37986 10722 37998
rect 3614 37938 3666 37950
rect 3614 37874 3666 37886
rect 3950 37938 4002 37950
rect 3950 37874 4002 37886
rect 4734 37938 4786 37950
rect 4734 37874 4786 37886
rect 5966 37938 6018 37950
rect 5966 37874 6018 37886
rect 6302 37938 6354 37950
rect 6302 37874 6354 37886
rect 6638 37938 6690 37950
rect 6638 37874 6690 37886
rect 7310 37938 7362 37950
rect 7310 37874 7362 37886
rect 7646 37938 7698 37950
rect 7646 37874 7698 37886
rect 7982 37938 8034 37950
rect 7982 37874 8034 37886
rect 9326 37938 9378 37950
rect 9326 37874 9378 37886
rect 9998 37938 10050 37950
rect 9998 37874 10050 37886
rect 10334 37938 10386 37950
rect 10334 37874 10386 37886
rect 1934 37826 1986 37838
rect 1934 37762 1986 37774
rect 2942 37826 2994 37838
rect 2942 37762 2994 37774
rect 3278 37826 3330 37838
rect 3278 37762 3330 37774
rect 4398 37826 4450 37838
rect 4398 37762 4450 37774
rect 5630 37826 5682 37838
rect 5630 37762 5682 37774
rect 8654 37826 8706 37838
rect 8654 37762 8706 37774
rect 1344 37658 42560 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 42560 37658
rect 1344 37572 42560 37606
rect 2158 37490 2210 37502
rect 2158 37426 2210 37438
rect 2942 37490 2994 37502
rect 2942 37426 2994 37438
rect 4622 37490 4674 37502
rect 4622 37426 4674 37438
rect 5294 37490 5346 37502
rect 5294 37426 5346 37438
rect 6302 37490 6354 37502
rect 6302 37426 6354 37438
rect 6974 37490 7026 37502
rect 6974 37426 7026 37438
rect 7422 37490 7474 37502
rect 7422 37426 7474 37438
rect 8430 37490 8482 37502
rect 8430 37426 8482 37438
rect 3278 37378 3330 37390
rect 3278 37314 3330 37326
rect 3950 37378 4002 37390
rect 3950 37314 4002 37326
rect 4958 37378 5010 37390
rect 4958 37314 5010 37326
rect 3614 37266 3666 37278
rect 3614 37202 3666 37214
rect 4286 37266 4338 37278
rect 5506 37214 5518 37266
rect 5570 37214 5582 37266
rect 8194 37214 8206 37266
rect 8258 37214 8270 37266
rect 4286 37202 4338 37214
rect 1822 37154 1874 37166
rect 1822 37090 1874 37102
rect 8990 37154 9042 37166
rect 8990 37090 9042 37102
rect 1344 36874 42560 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 42560 36874
rect 1344 36788 42560 36822
rect 5742 36594 5794 36606
rect 40674 36542 40686 36594
rect 40738 36542 40750 36594
rect 5742 36530 5794 36542
rect 1710 36482 1762 36494
rect 4398 36482 4450 36494
rect 3266 36430 3278 36482
rect 3330 36430 3342 36482
rect 1710 36418 1762 36430
rect 4398 36418 4450 36430
rect 2046 36370 2098 36382
rect 2046 36306 2098 36318
rect 2382 36370 2434 36382
rect 2382 36306 2434 36318
rect 2718 36370 2770 36382
rect 2718 36306 2770 36318
rect 4062 36370 4114 36382
rect 4062 36306 4114 36318
rect 4734 36370 4786 36382
rect 41682 36318 41694 36370
rect 41746 36318 41758 36370
rect 4734 36306 4786 36318
rect 3054 36258 3106 36270
rect 3054 36194 3106 36206
rect 3726 36258 3778 36270
rect 3726 36194 3778 36206
rect 1344 36090 42560 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 42560 36090
rect 1344 36004 42560 36038
rect 2046 35922 2098 35934
rect 2046 35858 2098 35870
rect 2942 35922 2994 35934
rect 2942 35858 2994 35870
rect 3950 35922 4002 35934
rect 3950 35858 4002 35870
rect 4398 35922 4450 35934
rect 4398 35858 4450 35870
rect 2382 35810 2434 35822
rect 2382 35746 2434 35758
rect 3278 35810 3330 35822
rect 3278 35746 3330 35758
rect 3614 35810 3666 35822
rect 3614 35746 3666 35758
rect 1710 35698 1762 35710
rect 1710 35634 1762 35646
rect 1344 35306 42560 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 42560 35306
rect 1344 35220 42560 35254
rect 3602 35086 3614 35138
rect 3666 35135 3678 35138
rect 3826 35135 3838 35138
rect 3666 35089 3838 35135
rect 3666 35086 3678 35089
rect 3826 35086 3838 35089
rect 3890 35086 3902 35138
rect 3838 35026 3890 35038
rect 40338 34974 40350 35026
rect 40402 34974 40414 35026
rect 3838 34962 3890 34974
rect 2706 34862 2718 34914
rect 2770 34862 2782 34914
rect 3278 34802 3330 34814
rect 2034 34750 2046 34802
rect 2098 34750 2110 34802
rect 39106 34750 39118 34802
rect 39170 34750 39182 34802
rect 3278 34738 3330 34750
rect 1344 34522 42560 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 42560 34522
rect 1344 34436 42560 34470
rect 2158 34354 2210 34366
rect 2158 34290 2210 34302
rect 1710 34242 1762 34254
rect 16258 34190 16270 34242
rect 16322 34190 16334 34242
rect 19730 34190 19742 34242
rect 19794 34190 19806 34242
rect 27234 34190 27246 34242
rect 27298 34190 27310 34242
rect 35634 34190 35646 34242
rect 35698 34190 35710 34242
rect 37314 34190 37326 34242
rect 37378 34190 37390 34242
rect 1710 34178 1762 34190
rect 15026 33966 15038 34018
rect 15090 33966 15102 34018
rect 18722 33966 18734 34018
rect 18786 33966 18798 34018
rect 26226 33966 26238 34018
rect 26290 33966 26302 34018
rect 34402 33966 34414 34018
rect 34466 33966 34478 34018
rect 38434 33966 38446 34018
rect 38498 33966 38510 34018
rect 1344 33738 42560 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 42560 33738
rect 1344 33652 42560 33686
rect 8754 33406 8766 33458
rect 8818 33406 8830 33458
rect 15138 33406 15150 33458
rect 15202 33406 15214 33458
rect 18386 33406 18398 33458
rect 18450 33406 18462 33458
rect 24546 33406 24558 33458
rect 24610 33406 24622 33458
rect 27122 33406 27134 33458
rect 27186 33406 27198 33458
rect 30146 33406 30158 33458
rect 30210 33406 30222 33458
rect 32946 33406 32958 33458
rect 33010 33406 33022 33458
rect 38434 33406 38446 33458
rect 38498 33406 38510 33458
rect 1710 33234 1762 33246
rect 1710 33170 1762 33182
rect 2046 33234 2098 33246
rect 9762 33182 9774 33234
rect 9826 33182 9838 33234
rect 16146 33182 16158 33234
rect 16210 33182 16222 33234
rect 17042 33182 17054 33234
rect 17106 33182 17118 33234
rect 25666 33182 25678 33234
rect 25730 33182 25742 33234
rect 28130 33182 28142 33234
rect 28194 33182 28206 33234
rect 31154 33182 31166 33234
rect 31218 33182 31230 33234
rect 33954 33182 33966 33234
rect 34018 33182 34030 33234
rect 39442 33182 39454 33234
rect 39506 33182 39518 33234
rect 2046 33170 2098 33182
rect 2494 33122 2546 33134
rect 2494 33058 2546 33070
rect 29374 33122 29426 33134
rect 29374 33058 29426 33070
rect 29822 33122 29874 33134
rect 29822 33058 29874 33070
rect 32734 33122 32786 33134
rect 32734 33058 32786 33070
rect 37214 33122 37266 33134
rect 37214 33058 37266 33070
rect 37662 33122 37714 33134
rect 37662 33058 37714 33070
rect 1344 32954 42560 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 42560 32954
rect 1344 32868 42560 32902
rect 30494 32786 30546 32798
rect 30494 32722 30546 32734
rect 32398 32786 32450 32798
rect 35074 32734 35086 32786
rect 35138 32734 35150 32786
rect 32398 32722 32450 32734
rect 1710 32674 1762 32686
rect 29710 32674 29762 32686
rect 5730 32622 5742 32674
rect 5794 32622 5806 32674
rect 9874 32622 9886 32674
rect 9938 32622 9950 32674
rect 15922 32622 15934 32674
rect 15986 32622 15998 32674
rect 20066 32622 20078 32674
rect 20130 32622 20142 32674
rect 1710 32610 1762 32622
rect 29710 32610 29762 32622
rect 31950 32562 32002 32574
rect 38110 32562 38162 32574
rect 39902 32562 39954 32574
rect 26898 32510 26910 32562
rect 26962 32510 26974 32562
rect 27458 32510 27470 32562
rect 27522 32510 27534 32562
rect 31154 32510 31166 32562
rect 31218 32510 31230 32562
rect 33506 32510 33518 32562
rect 33570 32510 33582 32562
rect 37538 32510 37550 32562
rect 37602 32510 37614 32562
rect 39106 32510 39118 32562
rect 39170 32510 39182 32562
rect 31950 32498 32002 32510
rect 38110 32498 38162 32510
rect 39902 32498 39954 32510
rect 40350 32562 40402 32574
rect 40350 32498 40402 32510
rect 19406 32450 19458 32462
rect 24670 32450 24722 32462
rect 6850 32398 6862 32450
rect 6914 32398 6926 32450
rect 10882 32398 10894 32450
rect 10946 32398 10958 32450
rect 14914 32398 14926 32450
rect 14978 32398 14990 32450
rect 21186 32398 21198 32450
rect 21250 32398 21262 32450
rect 24322 32398 24334 32450
rect 24386 32398 24398 32450
rect 19406 32386 19458 32398
rect 24670 32386 24722 32398
rect 26014 32450 26066 32462
rect 26226 32398 26238 32450
rect 26290 32398 26302 32450
rect 33394 32398 33406 32450
rect 33458 32398 33470 32450
rect 26014 32386 26066 32398
rect 31390 32338 31442 32350
rect 31390 32274 31442 32286
rect 34414 32338 34466 32350
rect 34414 32274 34466 32286
rect 39342 32338 39394 32350
rect 39342 32274 39394 32286
rect 1344 32170 42560 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 42560 32170
rect 1344 32084 42560 32118
rect 27022 32002 27074 32014
rect 27022 31938 27074 31950
rect 19182 31890 19234 31902
rect 8642 31838 8654 31890
rect 8706 31838 8718 31890
rect 11666 31838 11678 31890
rect 11730 31838 11742 31890
rect 19182 31826 19234 31838
rect 36542 31890 36594 31902
rect 37090 31838 37102 31890
rect 37154 31838 37166 31890
rect 40338 31838 40350 31890
rect 40402 31838 40414 31890
rect 36542 31826 36594 31838
rect 15710 31778 15762 31790
rect 23326 31778 23378 31790
rect 29038 31778 29090 31790
rect 33070 31778 33122 31790
rect 38222 31778 38274 31790
rect 2706 31726 2718 31778
rect 2770 31726 2782 31778
rect 16146 31726 16158 31778
rect 16210 31726 16222 31778
rect 20290 31726 20302 31778
rect 20354 31726 20366 31778
rect 23986 31726 23998 31778
rect 24050 31726 24062 31778
rect 28578 31726 28590 31778
rect 28642 31726 28654 31778
rect 29586 31726 29598 31778
rect 29650 31726 29662 31778
rect 33394 31726 33406 31778
rect 33458 31726 33470 31778
rect 37314 31726 37326 31778
rect 37378 31726 37390 31778
rect 15710 31714 15762 31726
rect 23326 31714 23378 31726
rect 29038 31714 29090 31726
rect 33070 31714 33122 31726
rect 38222 31714 38274 31726
rect 19742 31666 19794 31678
rect 2034 31614 2046 31666
rect 2098 31614 2110 31666
rect 9762 31614 9774 31666
rect 9826 31614 9838 31666
rect 12786 31614 12798 31666
rect 12850 31614 12862 31666
rect 19394 31614 19406 31666
rect 19458 31614 19470 31666
rect 19742 31602 19794 31614
rect 26238 31666 26290 31678
rect 39218 31614 39230 31666
rect 39282 31614 39294 31666
rect 26238 31602 26290 31614
rect 8430 31554 8482 31566
rect 8430 31490 8482 31502
rect 11230 31554 11282 31566
rect 11230 31490 11282 31502
rect 14590 31554 14642 31566
rect 20302 31554 20354 31566
rect 18386 31502 18398 31554
rect 18450 31502 18462 31554
rect 14590 31490 14642 31502
rect 20302 31490 20354 31502
rect 21422 31554 21474 31566
rect 21422 31490 21474 31502
rect 27358 31554 27410 31566
rect 27358 31490 27410 31502
rect 28478 31554 28530 31566
rect 32734 31554 32786 31566
rect 31938 31502 31950 31554
rect 32002 31502 32014 31554
rect 35746 31502 35758 31554
rect 35810 31502 35822 31554
rect 28478 31490 28530 31502
rect 32734 31490 32786 31502
rect 1344 31386 42560 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 42560 31386
rect 1344 31300 42560 31334
rect 4958 31218 5010 31230
rect 4958 31154 5010 31166
rect 8990 31218 9042 31230
rect 8990 31154 9042 31166
rect 9662 31218 9714 31230
rect 15262 31218 15314 31230
rect 14690 31166 14702 31218
rect 14754 31166 14766 31218
rect 9662 31154 9714 31166
rect 15262 31154 15314 31166
rect 15598 31218 15650 31230
rect 15598 31154 15650 31166
rect 17278 31218 17330 31230
rect 24782 31218 24834 31230
rect 29374 31218 29426 31230
rect 24210 31166 24222 31218
rect 24274 31166 24286 31218
rect 28578 31166 28590 31218
rect 28642 31166 28654 31218
rect 17278 31154 17330 31166
rect 24782 31154 24834 31166
rect 29374 31154 29426 31166
rect 30158 31218 30210 31230
rect 30158 31154 30210 31166
rect 32958 31218 33010 31230
rect 33618 31166 33630 31218
rect 33682 31166 33694 31218
rect 32958 31154 33010 31166
rect 5742 31106 5794 31118
rect 5742 31042 5794 31054
rect 18062 31106 18114 31118
rect 31826 31054 31838 31106
rect 31890 31054 31902 31106
rect 38882 31054 38894 31106
rect 38946 31054 38958 31106
rect 18062 31042 18114 31054
rect 8654 30994 8706 31006
rect 20750 30994 20802 31006
rect 2930 30942 2942 30994
rect 2994 30942 3006 30994
rect 8082 30942 8094 30994
rect 8146 30942 8158 30994
rect 10322 30942 10334 30994
rect 10386 30942 10398 30994
rect 10994 30942 11006 30994
rect 11058 30942 11070 30994
rect 11666 30942 11678 30994
rect 11730 30942 11742 30994
rect 12114 30942 12126 30994
rect 12178 30942 12190 30994
rect 20402 30942 20414 30994
rect 20466 30942 20478 30994
rect 8654 30930 8706 30942
rect 20750 30930 20802 30942
rect 21086 30994 21138 31006
rect 25678 30994 25730 31006
rect 36654 30994 36706 31006
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 26338 30942 26350 30994
rect 26402 30942 26414 30994
rect 36082 30942 36094 30994
rect 36146 30942 36158 30994
rect 21086 30930 21138 30942
rect 25678 30930 25730 30942
rect 36654 30930 36706 30942
rect 37438 30994 37490 31006
rect 37438 30930 37490 30942
rect 25342 30882 25394 30894
rect 1922 30830 1934 30882
rect 1986 30830 1998 30882
rect 10098 30830 10110 30882
rect 10162 30830 10174 30882
rect 10770 30830 10782 30882
rect 10834 30830 10846 30882
rect 25342 30818 25394 30830
rect 29710 30882 29762 30894
rect 36990 30882 37042 30894
rect 30594 30830 30606 30882
rect 30658 30830 30670 30882
rect 37874 30830 37886 30882
rect 37938 30830 37950 30882
rect 29710 30818 29762 30830
rect 36990 30818 37042 30830
rect 9426 30718 9438 30770
rect 9490 30767 9502 30770
rect 9762 30767 9774 30770
rect 9490 30721 9774 30767
rect 9490 30718 9502 30721
rect 9762 30718 9774 30721
rect 9826 30718 9838 30770
rect 36978 30718 36990 30770
rect 37042 30767 37054 30770
rect 37538 30767 37550 30770
rect 37042 30721 37550 30767
rect 37042 30718 37054 30721
rect 37538 30718 37550 30721
rect 37602 30718 37614 30770
rect 1344 30602 42560 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 42560 30602
rect 1344 30516 42560 30550
rect 29822 30434 29874 30446
rect 29822 30370 29874 30382
rect 27010 30270 27022 30322
rect 27074 30270 27086 30322
rect 35746 30270 35758 30322
rect 35810 30270 35822 30322
rect 2382 30210 2434 30222
rect 2382 30146 2434 30158
rect 3166 30210 3218 30222
rect 3166 30146 3218 30158
rect 7758 30210 7810 30222
rect 17054 30210 17106 30222
rect 8194 30158 8206 30210
rect 8258 30158 8270 30210
rect 11666 30158 11678 30210
rect 11730 30158 11742 30210
rect 12562 30158 12574 30210
rect 12626 30158 12638 30210
rect 13458 30158 13470 30210
rect 13522 30158 13534 30210
rect 14018 30158 14030 30210
rect 14082 30158 14094 30210
rect 7758 30146 7810 30158
rect 17054 30146 17106 30158
rect 17390 30210 17442 30222
rect 30270 30210 30322 30222
rect 33966 30210 34018 30222
rect 36990 30210 37042 30222
rect 40686 30210 40738 30222
rect 17826 30158 17838 30210
rect 17890 30158 17902 30210
rect 21746 30158 21758 30210
rect 21810 30158 21822 30210
rect 22194 30158 22206 30210
rect 22258 30158 22270 30210
rect 22754 30158 22766 30210
rect 22818 30158 22830 30210
rect 29586 30158 29598 30210
rect 29650 30158 29662 30210
rect 33394 30158 33406 30210
rect 33458 30158 33470 30210
rect 34738 30158 34750 30210
rect 34802 30158 34814 30210
rect 35858 30158 35870 30210
rect 35922 30158 35934 30210
rect 37650 30158 37662 30210
rect 37714 30158 37726 30210
rect 40898 30158 40910 30210
rect 40962 30158 40974 30210
rect 17390 30146 17442 30158
rect 30270 30146 30322 30158
rect 33966 30146 34018 30158
rect 36990 30146 37042 30158
rect 40686 30146 40738 30158
rect 1710 30098 1762 30110
rect 1710 30034 1762 30046
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 2718 30098 2770 30110
rect 25790 30098 25842 30110
rect 39902 30098 39954 30110
rect 11442 30046 11454 30098
rect 11506 30046 11518 30098
rect 12338 30046 12350 30098
rect 12402 30046 12414 30098
rect 21522 30046 21534 30098
rect 21586 30046 21598 30098
rect 28018 30046 28030 30098
rect 28082 30046 28094 30098
rect 2718 30034 2770 30046
rect 25790 30034 25842 30046
rect 39902 30034 39954 30046
rect 3614 29986 3666 29998
rect 11230 29986 11282 29998
rect 20862 29986 20914 29998
rect 26126 29986 26178 29998
rect 41022 29986 41074 29998
rect 10658 29934 10670 29986
rect 10722 29934 10734 29986
rect 16482 29934 16494 29986
rect 16546 29934 16558 29986
rect 20290 29934 20302 29986
rect 20354 29934 20366 29986
rect 25106 29934 25118 29986
rect 25170 29934 25182 29986
rect 31042 29934 31054 29986
rect 31106 29934 31118 29986
rect 34514 29934 34526 29986
rect 34578 29934 34590 29986
rect 3614 29922 3666 29934
rect 11230 29922 11282 29934
rect 20862 29922 20914 29934
rect 26126 29922 26178 29934
rect 41022 29922 41074 29934
rect 1344 29818 42560 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 42560 29818
rect 1344 29732 42560 29766
rect 2046 29650 2098 29662
rect 9102 29650 9154 29662
rect 8306 29598 8318 29650
rect 8370 29598 8382 29650
rect 2046 29586 2098 29598
rect 9102 29586 9154 29598
rect 9662 29650 9714 29662
rect 14366 29650 14418 29662
rect 13682 29598 13694 29650
rect 13746 29598 13758 29650
rect 9662 29586 9714 29598
rect 14366 29586 14418 29598
rect 15038 29650 15090 29662
rect 31390 29650 31442 29662
rect 23538 29598 23550 29650
rect 23602 29598 23614 29650
rect 15038 29586 15090 29598
rect 31390 29586 31442 29598
rect 31838 29650 31890 29662
rect 31838 29586 31890 29598
rect 33854 29650 33906 29662
rect 33854 29586 33906 29598
rect 36094 29650 36146 29662
rect 36094 29586 36146 29598
rect 36766 29650 36818 29662
rect 41022 29650 41074 29662
rect 37538 29598 37550 29650
rect 37602 29598 37614 29650
rect 36766 29586 36818 29598
rect 41022 29586 41074 29598
rect 19394 29486 19406 29538
rect 19458 29486 19470 29538
rect 24322 29486 24334 29538
rect 24386 29486 24398 29538
rect 27234 29486 27246 29538
rect 27298 29486 27310 29538
rect 30258 29486 30270 29538
rect 30322 29486 30334 29538
rect 35298 29486 35310 29538
rect 35362 29486 35374 29538
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 5630 29426 5682 29438
rect 10670 29426 10722 29438
rect 24110 29426 24162 29438
rect 40462 29426 40514 29438
rect 6066 29374 6078 29426
rect 6130 29374 6142 29426
rect 10322 29374 10334 29426
rect 10386 29374 10398 29426
rect 11330 29374 11342 29426
rect 11394 29374 11406 29426
rect 16594 29374 16606 29426
rect 16658 29374 16670 29426
rect 20514 29374 20526 29426
rect 20578 29374 20590 29426
rect 21074 29374 21086 29426
rect 21138 29374 21150 29426
rect 31714 29374 31726 29426
rect 31778 29374 31790 29426
rect 39890 29374 39902 29426
rect 39954 29374 39966 29426
rect 5630 29362 5682 29374
rect 10670 29362 10722 29374
rect 24110 29362 24162 29374
rect 40462 29362 40514 29374
rect 2494 29314 2546 29326
rect 14926 29314 14978 29326
rect 10098 29262 10110 29314
rect 10162 29262 10174 29314
rect 2494 29250 2546 29262
rect 14926 29250 14978 29262
rect 17502 29314 17554 29326
rect 17502 29250 17554 29262
rect 17950 29314 18002 29326
rect 24670 29314 24722 29326
rect 18386 29262 18398 29314
rect 18450 29262 18462 29314
rect 17950 29250 18002 29262
rect 24670 29250 24722 29262
rect 25342 29314 25394 29326
rect 28142 29314 28194 29326
rect 33406 29314 33458 29326
rect 36542 29314 36594 29326
rect 26226 29262 26238 29314
rect 26290 29262 26302 29314
rect 29026 29262 29038 29314
rect 29090 29262 29102 29314
rect 34178 29262 34190 29314
rect 34242 29262 34254 29314
rect 25342 29250 25394 29262
rect 28142 29250 28194 29262
rect 33406 29250 33458 29262
rect 36542 29250 36594 29262
rect 15822 29202 15874 29214
rect 15822 29138 15874 29150
rect 1344 29034 42560 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 42560 29034
rect 1344 28948 42560 28982
rect 9214 28866 9266 28878
rect 9214 28802 9266 28814
rect 13022 28866 13074 28878
rect 13022 28802 13074 28814
rect 15934 28866 15986 28878
rect 15934 28802 15986 28814
rect 36878 28866 36930 28878
rect 36878 28802 36930 28814
rect 13682 28702 13694 28754
rect 13746 28702 13758 28754
rect 19842 28702 19854 28754
rect 19906 28702 19918 28754
rect 22306 28702 22318 28754
rect 22370 28702 22382 28754
rect 30482 28702 30494 28754
rect 30546 28702 30558 28754
rect 33282 28702 33294 28754
rect 33346 28702 33358 28754
rect 35298 28702 35310 28754
rect 35362 28702 35374 28754
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 2494 28642 2546 28654
rect 2494 28578 2546 28590
rect 5742 28642 5794 28654
rect 9550 28642 9602 28654
rect 20638 28642 20690 28654
rect 6178 28590 6190 28642
rect 6242 28590 6254 28642
rect 9874 28590 9886 28642
rect 9938 28590 9950 28642
rect 13570 28590 13582 28642
rect 13634 28590 13646 28642
rect 18946 28590 18958 28642
rect 19010 28590 19022 28642
rect 19506 28590 19518 28642
rect 19570 28590 19582 28642
rect 5742 28578 5794 28590
rect 9550 28578 9602 28590
rect 20638 28578 20690 28590
rect 24334 28642 24386 28654
rect 28030 28642 28082 28654
rect 36318 28642 36370 28654
rect 24770 28590 24782 28642
rect 24834 28590 24846 28642
rect 35074 28590 35086 28642
rect 35138 28590 35150 28642
rect 40002 28590 40014 28642
rect 40066 28590 40078 28642
rect 40450 28590 40462 28642
rect 40514 28590 40526 28642
rect 24334 28578 24386 28590
rect 28030 28578 28082 28590
rect 36318 28578 36370 28590
rect 2046 28530 2098 28542
rect 16718 28530 16770 28542
rect 14466 28478 14478 28530
rect 14530 28478 14542 28530
rect 2046 28466 2098 28478
rect 16718 28466 16770 28478
rect 20190 28530 20242 28542
rect 23538 28478 23550 28530
rect 23602 28478 23614 28530
rect 31490 28478 31502 28530
rect 31554 28478 31566 28530
rect 34290 28478 34302 28530
rect 34354 28478 34366 28530
rect 20190 28466 20242 28478
rect 15038 28418 15090 28430
rect 27806 28418 27858 28430
rect 8642 28366 8654 28418
rect 8706 28366 8718 28418
rect 12338 28366 12350 28418
rect 12402 28366 12414 28418
rect 27234 28366 27246 28418
rect 27298 28366 27310 28418
rect 15038 28354 15090 28366
rect 27806 28354 27858 28366
rect 28142 28418 28194 28430
rect 28142 28354 28194 28366
rect 29262 28418 29314 28430
rect 37650 28366 37662 28418
rect 37714 28366 37726 28418
rect 29262 28354 29314 28366
rect 1344 28250 42560 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 42560 28250
rect 1344 28164 42560 28198
rect 9102 28082 9154 28094
rect 9102 28018 9154 28030
rect 12238 28082 12290 28094
rect 16158 28082 16210 28094
rect 15586 28030 15598 28082
rect 15650 28030 15662 28082
rect 12238 28018 12290 28030
rect 16158 28018 16210 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 29598 28082 29650 28094
rect 29598 28018 29650 28030
rect 37662 28082 37714 28094
rect 37662 28018 37714 28030
rect 39790 28082 39842 28094
rect 39790 28018 39842 28030
rect 40238 28082 40290 28094
rect 40238 28018 40290 28030
rect 2046 27970 2098 27982
rect 2046 27906 2098 27918
rect 8318 27970 8370 27982
rect 16830 27970 16882 27982
rect 25566 27970 25618 27982
rect 9874 27918 9886 27970
rect 9938 27918 9950 27970
rect 16482 27918 16494 27970
rect 16546 27918 16558 27970
rect 19730 27918 19742 27970
rect 19794 27918 19806 27970
rect 25218 27918 25230 27970
rect 25282 27918 25294 27970
rect 8318 27906 8370 27918
rect 16830 27906 16882 27918
rect 25566 27906 25618 27918
rect 36878 27970 36930 27982
rect 38882 27918 38894 27970
rect 38946 27918 38958 27970
rect 36878 27906 36930 27918
rect 1710 27858 1762 27870
rect 1710 27794 1762 27806
rect 5630 27858 5682 27870
rect 12686 27858 12738 27870
rect 33966 27858 34018 27870
rect 6066 27806 6078 27858
rect 6130 27806 6142 27858
rect 13122 27806 13134 27858
rect 13186 27806 13198 27858
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 34626 27806 34638 27858
rect 34690 27806 34702 27858
rect 5630 27794 5682 27806
rect 12686 27794 12738 27806
rect 33966 27794 34018 27806
rect 2494 27746 2546 27758
rect 21198 27746 21250 27758
rect 11218 27694 11230 27746
rect 11282 27694 11294 27746
rect 18386 27694 18398 27746
rect 18450 27694 18462 27746
rect 2494 27682 2546 27694
rect 21198 27682 21250 27694
rect 26126 27746 26178 27758
rect 37874 27694 37886 27746
rect 37938 27694 37950 27746
rect 26126 27682 26178 27694
rect 1344 27466 42560 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 42560 27466
rect 1344 27380 42560 27414
rect 25006 27298 25058 27310
rect 25006 27234 25058 27246
rect 29038 27298 29090 27310
rect 39902 27298 39954 27310
rect 32834 27246 32846 27298
rect 32898 27295 32910 27298
rect 33506 27295 33518 27298
rect 32898 27249 33518 27295
rect 32898 27246 32910 27249
rect 33506 27246 33518 27249
rect 33570 27246 33582 27298
rect 29038 27234 29090 27246
rect 39902 27234 39954 27246
rect 6850 27134 6862 27186
rect 6914 27134 6926 27186
rect 14130 27134 14142 27186
rect 14194 27134 14206 27186
rect 18274 27134 18286 27186
rect 18338 27134 18350 27186
rect 34962 27134 34974 27186
rect 35026 27134 35038 27186
rect 37986 27134 37998 27186
rect 38050 27134 38062 27186
rect 12686 27074 12738 27086
rect 28702 27074 28754 27086
rect 32734 27074 32786 27086
rect 2818 27022 2830 27074
rect 2882 27022 2894 27074
rect 8866 27022 8878 27074
rect 8930 27022 8942 27074
rect 12226 27022 12238 27074
rect 12290 27022 12302 27074
rect 14914 27022 14926 27074
rect 14978 27022 14990 27074
rect 16146 27022 16158 27074
rect 16210 27022 16222 27074
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 28130 27022 28142 27074
rect 28194 27022 28206 27074
rect 32162 27022 32174 27074
rect 32226 27022 32238 27074
rect 40114 27022 40126 27074
rect 40178 27022 40190 27074
rect 12686 27010 12738 27022
rect 28702 27010 28754 27022
rect 32734 27010 32786 27022
rect 9998 26962 10050 26974
rect 7858 26910 7870 26962
rect 7922 26910 7934 26962
rect 8642 26910 8654 26962
rect 8706 26910 8718 26962
rect 9998 26898 10050 26910
rect 29822 26962 29874 26974
rect 29822 26898 29874 26910
rect 33182 26962 33234 26974
rect 33182 26898 33234 26910
rect 33518 26962 33570 26974
rect 35970 26910 35982 26962
rect 36034 26910 36046 26962
rect 39330 26910 39342 26962
rect 39394 26910 39406 26962
rect 33518 26898 33570 26910
rect 2158 26850 2210 26862
rect 2158 26786 2210 26798
rect 9214 26850 9266 26862
rect 9214 26786 9266 26798
rect 21982 26850 22034 26862
rect 25778 26798 25790 26850
rect 25842 26798 25854 26850
rect 21982 26786 22034 26798
rect 1344 26682 42560 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 42560 26682
rect 1344 26596 42560 26630
rect 2942 26514 2994 26526
rect 2942 26450 2994 26462
rect 3614 26514 3666 26526
rect 3614 26450 3666 26462
rect 5406 26514 5458 26526
rect 17502 26514 17554 26526
rect 6178 26462 6190 26514
rect 6242 26462 6254 26514
rect 16370 26462 16382 26514
rect 16434 26462 16446 26514
rect 5406 26450 5458 26462
rect 17502 26450 17554 26462
rect 25902 26514 25954 26526
rect 25902 26450 25954 26462
rect 38782 26514 38834 26526
rect 38782 26450 38834 26462
rect 10110 26402 10162 26414
rect 16942 26402 16994 26414
rect 23774 26402 23826 26414
rect 9762 26350 9774 26402
rect 9826 26350 9838 26402
rect 10546 26350 10558 26402
rect 10610 26350 10622 26402
rect 19394 26350 19406 26402
rect 19458 26350 19470 26402
rect 20178 26350 20190 26402
rect 20242 26350 20254 26402
rect 10110 26338 10162 26350
rect 16942 26338 16994 26350
rect 23774 26338 23826 26350
rect 3278 26290 3330 26302
rect 9102 26290 9154 26302
rect 8530 26238 8542 26290
rect 8594 26238 8606 26290
rect 3278 26226 3330 26238
rect 9102 26226 9154 26238
rect 13022 26290 13074 26302
rect 21086 26290 21138 26302
rect 13346 26238 13358 26290
rect 13410 26238 13422 26290
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 20402 26238 20414 26290
rect 20466 26238 20478 26290
rect 21522 26238 21534 26290
rect 21586 26238 21598 26290
rect 25778 26238 25790 26290
rect 25842 26238 25854 26290
rect 28354 26238 28366 26290
rect 28418 26238 28430 26290
rect 33170 26238 33182 26290
rect 33234 26238 33246 26290
rect 38658 26238 38670 26290
rect 38722 26238 38734 26290
rect 13022 26226 13074 26238
rect 21086 26226 21138 26238
rect 1822 26178 1874 26190
rect 25342 26178 25394 26190
rect 39902 26178 39954 26190
rect 2258 26126 2270 26178
rect 2322 26126 2334 26178
rect 11778 26126 11790 26178
rect 11842 26126 11854 26178
rect 18386 26126 18398 26178
rect 18450 26126 18462 26178
rect 28914 26126 28926 26178
rect 28978 26126 28990 26178
rect 35634 26126 35646 26178
rect 35698 26126 35710 26178
rect 1822 26114 1874 26126
rect 25342 26114 25394 26126
rect 39902 26114 39954 26126
rect 24558 26066 24610 26078
rect 17266 26014 17278 26066
rect 17330 26063 17342 26066
rect 17602 26063 17614 26066
rect 17330 26017 17614 26063
rect 17330 26014 17342 26017
rect 17602 26014 17614 26017
rect 17666 26014 17678 26066
rect 24558 26002 24610 26014
rect 1344 25898 42560 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 42560 25898
rect 1344 25812 42560 25846
rect 22430 25730 22482 25742
rect 9314 25678 9326 25730
rect 9378 25727 9390 25730
rect 9650 25727 9662 25730
rect 9378 25681 9662 25727
rect 9378 25678 9390 25681
rect 9650 25678 9662 25681
rect 9714 25678 9726 25730
rect 22430 25666 22482 25678
rect 26462 25730 26514 25742
rect 26462 25666 26514 25678
rect 40798 25730 40850 25742
rect 40798 25666 40850 25678
rect 7310 25618 7362 25630
rect 9550 25618 9602 25630
rect 20526 25618 20578 25630
rect 6962 25566 6974 25618
rect 7026 25566 7038 25618
rect 9090 25566 9102 25618
rect 9154 25566 9166 25618
rect 11442 25566 11454 25618
rect 11506 25566 11518 25618
rect 17490 25566 17502 25618
rect 17554 25566 17566 25618
rect 7310 25554 7362 25566
rect 9550 25554 9602 25566
rect 20526 25554 20578 25566
rect 26798 25618 26850 25630
rect 26798 25554 26850 25566
rect 27246 25618 27298 25630
rect 27246 25554 27298 25566
rect 2942 25506 2994 25518
rect 22990 25506 23042 25518
rect 29262 25506 29314 25518
rect 36318 25506 36370 25518
rect 16258 25454 16270 25506
rect 16322 25454 16334 25506
rect 22194 25454 22206 25506
rect 22258 25454 22270 25506
rect 23314 25454 23326 25506
rect 23378 25454 23390 25506
rect 29698 25454 29710 25506
rect 29762 25454 29774 25506
rect 35970 25454 35982 25506
rect 36034 25454 36046 25506
rect 2942 25442 2994 25454
rect 22990 25442 23042 25454
rect 29262 25442 29314 25454
rect 36318 25442 36370 25454
rect 37102 25506 37154 25518
rect 37762 25454 37774 25506
rect 37826 25454 37838 25506
rect 37102 25442 37154 25454
rect 33630 25394 33682 25406
rect 8082 25342 8094 25394
rect 8146 25342 8158 25394
rect 12786 25342 12798 25394
rect 12850 25342 12862 25394
rect 33630 25330 33682 25342
rect 2158 25282 2210 25294
rect 32734 25282 32786 25294
rect 25890 25230 25902 25282
rect 25954 25230 25966 25282
rect 32162 25230 32174 25282
rect 32226 25230 32238 25282
rect 2158 25218 2210 25230
rect 32734 25218 32786 25230
rect 32846 25282 32898 25294
rect 40002 25230 40014 25282
rect 40066 25230 40078 25282
rect 32846 25218 32898 25230
rect 1344 25114 42560 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 42560 25114
rect 1344 25028 42560 25062
rect 16606 24946 16658 24958
rect 23438 24946 23490 24958
rect 22306 24894 22318 24946
rect 22370 24894 22382 24946
rect 16606 24882 16658 24894
rect 23438 24882 23490 24894
rect 25902 24946 25954 24958
rect 25902 24882 25954 24894
rect 30718 24946 30770 24958
rect 30718 24882 30770 24894
rect 33182 24946 33234 24958
rect 33182 24882 33234 24894
rect 36094 24946 36146 24958
rect 36094 24882 36146 24894
rect 36542 24946 36594 24958
rect 36542 24882 36594 24894
rect 39342 24946 39394 24958
rect 39342 24882 39394 24894
rect 15822 24834 15874 24846
rect 18846 24834 18898 24846
rect 7522 24782 7534 24834
rect 7586 24782 7598 24834
rect 10434 24782 10446 24834
rect 10498 24782 10510 24834
rect 17378 24782 17390 24834
rect 17442 24782 17454 24834
rect 30146 24782 30158 24834
rect 30210 24782 30222 24834
rect 32162 24782 32174 24834
rect 32226 24782 32238 24834
rect 35298 24782 35310 24834
rect 35362 24782 35374 24834
rect 37874 24782 37886 24834
rect 37938 24782 37950 24834
rect 15822 24770 15874 24782
rect 18846 24770 18898 24782
rect 19630 24722 19682 24734
rect 39902 24722 39954 24734
rect 2930 24670 2942 24722
rect 2994 24670 3006 24722
rect 15474 24670 15486 24722
rect 15538 24670 15550 24722
rect 17602 24670 17614 24722
rect 17666 24670 17678 24722
rect 18274 24670 18286 24722
rect 18338 24670 18350 24722
rect 20066 24670 20078 24722
rect 20130 24670 20142 24722
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 30594 24670 30606 24722
rect 30658 24670 30670 24722
rect 31714 24670 31726 24722
rect 31778 24670 31790 24722
rect 39106 24670 39118 24722
rect 39170 24670 39182 24722
rect 19630 24658 19682 24670
rect 39902 24658 39954 24670
rect 33630 24610 33682 24622
rect 1922 24558 1934 24610
rect 1986 24558 1998 24610
rect 6178 24558 6190 24610
rect 6242 24558 6254 24610
rect 16146 24558 16158 24610
rect 16210 24558 16222 24610
rect 18050 24558 18062 24610
rect 18114 24558 18126 24610
rect 19170 24558 19182 24610
rect 19234 24558 19246 24610
rect 28802 24558 28814 24610
rect 28866 24558 28878 24610
rect 34066 24558 34078 24610
rect 34130 24558 34142 24610
rect 36866 24558 36878 24610
rect 36930 24558 36942 24610
rect 33630 24546 33682 24558
rect 23102 24498 23154 24510
rect 35970 24446 35982 24498
rect 36034 24495 36046 24498
rect 36642 24495 36654 24498
rect 36034 24449 36654 24495
rect 36034 24446 36046 24449
rect 36642 24446 36654 24449
rect 36706 24446 36718 24498
rect 23102 24434 23154 24446
rect 1344 24330 42560 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 42560 24330
rect 1344 24244 42560 24278
rect 34302 24162 34354 24174
rect 34302 24098 34354 24110
rect 36990 24162 37042 24174
rect 36990 24098 37042 24110
rect 20414 24050 20466 24062
rect 35758 24050 35810 24062
rect 15250 23998 15262 24050
rect 15314 23998 15326 24050
rect 22306 23998 22318 24050
rect 22370 23998 22382 24050
rect 25106 23998 25118 24050
rect 25170 23998 25182 24050
rect 20414 23986 20466 23998
rect 35758 23986 35810 23998
rect 36206 24050 36258 24062
rect 36206 23986 36258 23998
rect 10894 23938 10946 23950
rect 10546 23886 10558 23938
rect 10610 23886 10622 23938
rect 10894 23874 10946 23886
rect 16494 23938 16546 23950
rect 30830 23938 30882 23950
rect 40462 23938 40514 23950
rect 17154 23886 17166 23938
rect 17218 23886 17230 23938
rect 31266 23886 31278 23938
rect 31330 23886 31342 23938
rect 35074 23886 35086 23938
rect 35138 23886 35150 23938
rect 40114 23886 40126 23938
rect 40178 23886 40190 23938
rect 16494 23874 16546 23886
rect 30830 23874 30882 23886
rect 40462 23874 40514 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 11902 23826 11954 23838
rect 11554 23774 11566 23826
rect 11618 23774 11630 23826
rect 2046 23762 2098 23774
rect 11902 23762 11954 23774
rect 12350 23826 12402 23838
rect 19406 23826 19458 23838
rect 33518 23826 33570 23838
rect 14242 23774 14254 23826
rect 14306 23774 14318 23826
rect 20738 23774 20750 23826
rect 20802 23774 20814 23826
rect 23314 23774 23326 23826
rect 23378 23774 23390 23826
rect 26114 23774 26126 23826
rect 26178 23774 26190 23826
rect 12350 23762 12402 23774
rect 19406 23762 19458 23774
rect 33518 23762 33570 23774
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 7422 23714 7474 23726
rect 15710 23714 15762 23726
rect 8194 23662 8206 23714
rect 8258 23662 8270 23714
rect 7422 23650 7474 23662
rect 15710 23650 15762 23662
rect 20190 23714 20242 23726
rect 20190 23650 20242 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 30270 23714 30322 23726
rect 30270 23650 30322 23662
rect 35198 23714 35250 23726
rect 37762 23662 37774 23714
rect 37826 23662 37838 23714
rect 35198 23650 35250 23662
rect 1344 23546 42560 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 42560 23546
rect 1344 23460 42560 23494
rect 11230 23378 11282 23390
rect 11230 23314 11282 23326
rect 17502 23378 17554 23390
rect 21422 23378 21474 23390
rect 20738 23326 20750 23378
rect 20802 23326 20814 23378
rect 17502 23314 17554 23326
rect 21422 23314 21474 23326
rect 26462 23378 26514 23390
rect 26462 23314 26514 23326
rect 26910 23378 26962 23390
rect 39790 23378 39842 23390
rect 39218 23326 39230 23378
rect 39282 23326 39294 23378
rect 26910 23314 26962 23326
rect 39790 23314 39842 23326
rect 2382 23266 2434 23278
rect 12574 23266 12626 23278
rect 6962 23214 6974 23266
rect 7026 23214 7038 23266
rect 2382 23202 2434 23214
rect 12574 23202 12626 23214
rect 15934 23266 15986 23278
rect 22306 23214 22318 23266
rect 22370 23214 22382 23266
rect 35074 23214 35086 23266
rect 35138 23214 35150 23266
rect 15934 23202 15986 23214
rect 5294 23154 5346 23166
rect 15486 23154 15538 23166
rect 36094 23154 36146 23166
rect 40126 23154 40178 23166
rect 4722 23102 4734 23154
rect 4786 23102 4798 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 17826 23102 17838 23154
rect 17890 23102 17902 23154
rect 18274 23102 18286 23154
rect 18338 23102 18350 23154
rect 27234 23102 27246 23154
rect 27298 23102 27310 23154
rect 36754 23102 36766 23154
rect 36818 23102 36830 23154
rect 5294 23090 5346 23102
rect 15486 23090 15538 23102
rect 36094 23090 36146 23102
rect 40126 23090 40178 23102
rect 5630 23042 5682 23054
rect 33182 23042 33234 23054
rect 7970 22990 7982 23042
rect 8034 22990 8046 23042
rect 16258 22990 16270 23042
rect 16322 22990 16334 23042
rect 23426 22990 23438 23042
rect 23490 22990 23502 23042
rect 30146 22990 30158 23042
rect 30210 22990 30222 23042
rect 5630 22978 5682 22990
rect 33182 22978 33234 22990
rect 33742 23042 33794 23054
rect 34066 22990 34078 23042
rect 34130 22990 34142 23042
rect 33742 22978 33794 22990
rect 1598 22930 1650 22942
rect 1598 22866 1650 22878
rect 11790 22930 11842 22942
rect 33170 22878 33182 22930
rect 33234 22927 33246 22930
rect 33618 22927 33630 22930
rect 33234 22881 33630 22927
rect 33234 22878 33246 22881
rect 33618 22878 33630 22881
rect 33682 22878 33694 22930
rect 11790 22866 11842 22878
rect 1344 22762 42560 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 42560 22762
rect 1344 22676 42560 22710
rect 15710 22594 15762 22606
rect 15710 22530 15762 22542
rect 39902 22594 39954 22606
rect 39902 22530 39954 22542
rect 2494 22482 2546 22494
rect 13582 22482 13634 22494
rect 14926 22482 14978 22494
rect 8082 22430 8094 22482
rect 8146 22430 8158 22482
rect 14578 22430 14590 22482
rect 14642 22430 14654 22482
rect 2494 22418 2546 22430
rect 13582 22418 13634 22430
rect 14926 22418 14978 22430
rect 37102 22482 37154 22494
rect 37102 22418 37154 22430
rect 37550 22482 37602 22494
rect 41022 22482 41074 22494
rect 37986 22430 37998 22482
rect 38050 22430 38062 22482
rect 37550 22418 37602 22430
rect 41022 22418 41074 22430
rect 1710 22370 1762 22382
rect 1710 22306 1762 22318
rect 9550 22370 9602 22382
rect 19182 22370 19234 22382
rect 22878 22370 22930 22382
rect 32510 22370 32562 22382
rect 9874 22318 9886 22370
rect 9938 22318 9950 22370
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 20402 22318 20414 22370
rect 20466 22318 20478 22370
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 23314 22318 23326 22370
rect 23378 22318 23390 22370
rect 27010 22318 27022 22370
rect 27074 22318 27086 22370
rect 27682 22318 27694 22370
rect 27746 22318 27758 22370
rect 32162 22318 32174 22370
rect 32226 22318 32238 22370
rect 9550 22306 9602 22318
rect 19182 22306 19234 22318
rect 22878 22306 22930 22318
rect 32510 22306 32562 22318
rect 32846 22370 32898 22382
rect 33506 22318 33518 22370
rect 33570 22318 33582 22370
rect 40002 22318 40014 22370
rect 40066 22318 40078 22370
rect 32846 22306 32898 22318
rect 2046 22258 2098 22270
rect 14254 22258 14306 22270
rect 7074 22206 7086 22258
rect 7138 22206 7150 22258
rect 13906 22206 13918 22258
rect 13970 22206 13982 22258
rect 2046 22194 2098 22206
rect 14254 22194 14306 22206
rect 26350 22258 26402 22270
rect 26350 22194 26402 22206
rect 35758 22258 35810 22270
rect 38994 22206 39006 22258
rect 39058 22206 39070 22258
rect 35758 22194 35810 22206
rect 13022 22146 13074 22158
rect 20638 22146 20690 22158
rect 12450 22094 12462 22146
rect 12514 22094 12526 22146
rect 16482 22094 16494 22146
rect 16546 22094 16558 22146
rect 13022 22082 13074 22094
rect 20638 22082 20690 22094
rect 21758 22146 21810 22158
rect 27246 22146 27298 22158
rect 29038 22146 29090 22158
rect 36542 22146 36594 22158
rect 25554 22094 25566 22146
rect 25618 22094 25630 22146
rect 28242 22094 28254 22146
rect 28306 22094 28318 22146
rect 29586 22094 29598 22146
rect 29650 22094 29662 22146
rect 21758 22082 21810 22094
rect 27246 22082 27298 22094
rect 29038 22082 29090 22094
rect 36542 22082 36594 22094
rect 1344 21978 42560 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 42560 21978
rect 1344 21892 42560 21926
rect 5294 21810 5346 21822
rect 5294 21746 5346 21758
rect 9438 21810 9490 21822
rect 17502 21810 17554 21822
rect 10210 21758 10222 21810
rect 10274 21758 10286 21810
rect 16146 21758 16158 21810
rect 16210 21758 16222 21810
rect 9438 21746 9490 21758
rect 17502 21746 17554 21758
rect 20974 21810 21026 21822
rect 33182 21810 33234 21822
rect 38446 21810 38498 21822
rect 21746 21758 21758 21810
rect 21810 21758 21822 21810
rect 28018 21758 28030 21810
rect 28082 21758 28094 21810
rect 32050 21758 32062 21810
rect 32114 21758 32126 21810
rect 37426 21758 37438 21810
rect 37490 21758 37502 21810
rect 20974 21746 21026 21758
rect 33182 21746 33234 21758
rect 38446 21746 38498 21758
rect 39566 21810 39618 21822
rect 39566 21746 39618 21758
rect 4510 21698 4562 21710
rect 6962 21646 6974 21698
rect 7026 21646 7038 21698
rect 20066 21646 20078 21698
rect 20130 21646 20142 21698
rect 4510 21634 4562 21646
rect 1822 21586 1874 21598
rect 5630 21586 5682 21598
rect 13134 21586 13186 21598
rect 2146 21534 2158 21586
rect 2210 21534 2222 21586
rect 12450 21534 12462 21586
rect 12514 21534 12526 21586
rect 1822 21522 1874 21534
rect 5630 21522 5682 21534
rect 13134 21522 13186 21534
rect 13470 21586 13522 21598
rect 24446 21586 24498 21598
rect 13794 21534 13806 21586
rect 13858 21534 13870 21586
rect 23986 21534 23998 21586
rect 24050 21534 24062 21586
rect 13470 21522 13522 21534
rect 24446 21522 24498 21534
rect 25118 21586 25170 21598
rect 29150 21586 29202 21598
rect 34638 21586 34690 21598
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 29586 21534 29598 21586
rect 29650 21534 29662 21586
rect 33394 21534 33406 21586
rect 33458 21534 33470 21586
rect 35074 21534 35086 21586
rect 35138 21534 35150 21586
rect 38658 21534 38670 21586
rect 38722 21534 38734 21586
rect 39778 21534 39790 21586
rect 39842 21534 39854 21586
rect 25118 21522 25170 21534
rect 29150 21522 29202 21534
rect 34638 21522 34690 21534
rect 7970 21422 7982 21474
rect 8034 21422 8046 21474
rect 18722 21422 18734 21474
rect 18786 21422 18798 21474
rect 16942 21362 16994 21374
rect 16942 21298 16994 21310
rect 28814 21362 28866 21374
rect 28814 21298 28866 21310
rect 32622 21362 32674 21374
rect 32622 21298 32674 21310
rect 38110 21362 38162 21374
rect 38110 21298 38162 21310
rect 1344 21194 42560 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 42560 21194
rect 1344 21108 42560 21142
rect 17054 21026 17106 21038
rect 17054 20962 17106 20974
rect 34414 21026 34466 21038
rect 34626 20974 34638 21026
rect 34690 21023 34702 21026
rect 35186 21023 35198 21026
rect 34690 20977 35198 21023
rect 34690 20974 34702 20977
rect 35186 20974 35198 20977
rect 35250 20974 35262 21026
rect 34414 20962 34466 20974
rect 11006 20914 11058 20926
rect 3826 20862 3838 20914
rect 3890 20862 3902 20914
rect 10770 20862 10782 20914
rect 10834 20862 10846 20914
rect 11006 20850 11058 20862
rect 11454 20914 11506 20926
rect 11454 20850 11506 20862
rect 12910 20914 12962 20926
rect 12910 20850 12962 20862
rect 17390 20914 17442 20926
rect 19742 20914 19794 20926
rect 34862 20914 34914 20926
rect 19058 20862 19070 20914
rect 19122 20862 19134 20914
rect 24882 20862 24894 20914
rect 24946 20862 24958 20914
rect 17390 20850 17442 20862
rect 19742 20850 19794 20862
rect 34862 20850 34914 20862
rect 35198 20914 35250 20926
rect 35198 20850 35250 20862
rect 37214 20914 37266 20926
rect 37214 20850 37266 20862
rect 37774 20914 37826 20926
rect 40014 20914 40066 20926
rect 37986 20862 37998 20914
rect 38050 20862 38062 20914
rect 37774 20850 37826 20862
rect 40014 20850 40066 20862
rect 1710 20802 1762 20814
rect 6750 20802 6802 20814
rect 13582 20802 13634 20814
rect 20862 20802 20914 20814
rect 30942 20802 30994 20814
rect 6178 20750 6190 20802
rect 6242 20750 6254 20802
rect 7298 20750 7310 20802
rect 7362 20750 7374 20802
rect 13906 20750 13918 20802
rect 13970 20750 13982 20802
rect 21410 20750 21422 20802
rect 21474 20750 21486 20802
rect 27570 20750 27582 20802
rect 27634 20750 27646 20802
rect 31378 20750 31390 20802
rect 31442 20750 31454 20802
rect 1710 20738 1762 20750
rect 6750 20738 6802 20750
rect 13582 20738 13634 20750
rect 20862 20738 20914 20750
rect 30942 20738 30994 20750
rect 2046 20690 2098 20702
rect 16270 20690 16322 20702
rect 2706 20638 2718 20690
rect 2770 20638 2782 20690
rect 17938 20638 17950 20690
rect 18002 20638 18014 20690
rect 38994 20638 39006 20690
rect 39058 20638 39070 20690
rect 2046 20626 2098 20638
rect 16270 20626 16322 20638
rect 10446 20578 10498 20590
rect 5954 20526 5966 20578
rect 6018 20526 6030 20578
rect 9650 20526 9662 20578
rect 9714 20526 9726 20578
rect 10446 20514 10498 20526
rect 27694 20578 27746 20590
rect 33730 20526 33742 20578
rect 33794 20526 33806 20578
rect 27694 20514 27746 20526
rect 1344 20410 42560 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 42560 20410
rect 1344 20324 42560 20358
rect 1822 20242 1874 20254
rect 1822 20178 1874 20190
rect 3614 20242 3666 20254
rect 16606 20242 16658 20254
rect 5842 20190 5854 20242
rect 5906 20190 5918 20242
rect 3614 20178 3666 20190
rect 16606 20178 16658 20190
rect 33742 20242 33794 20254
rect 33742 20178 33794 20190
rect 10670 20130 10722 20142
rect 30046 20130 30098 20142
rect 25554 20078 25566 20130
rect 25618 20078 25630 20130
rect 10670 20066 10722 20078
rect 30046 20066 30098 20078
rect 35870 20130 35922 20142
rect 35870 20066 35922 20078
rect 8766 20018 8818 20030
rect 32510 20018 32562 20030
rect 38782 20018 38834 20030
rect 3378 19966 3390 20018
rect 3442 19966 3454 20018
rect 4050 19966 4062 20018
rect 4114 19966 4126 20018
rect 8082 19966 8094 20018
rect 8146 19966 8158 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 27234 19966 27246 20018
rect 27298 19966 27310 20018
rect 27794 19966 27806 20018
rect 27858 19966 27870 20018
rect 33506 19966 33518 20018
rect 33570 19966 33582 20018
rect 38098 19966 38110 20018
rect 38162 19966 38174 20018
rect 8766 19954 8818 19966
rect 32510 19954 32562 19966
rect 38782 19954 38834 19966
rect 39118 20018 39170 20030
rect 39118 19954 39170 19966
rect 9774 19906 9826 19918
rect 15262 19906 15314 19918
rect 21758 19906 21810 19918
rect 11890 19854 11902 19906
rect 11954 19854 11966 19906
rect 20066 19854 20078 19906
rect 20130 19854 20142 19906
rect 9774 19842 9826 19854
rect 15262 19842 15314 19854
rect 21758 19842 21810 19854
rect 26686 19906 26738 19918
rect 26686 19842 26738 19854
rect 4174 19794 4226 19806
rect 4174 19730 4226 19742
rect 5070 19794 5122 19806
rect 5070 19730 5122 19742
rect 30830 19794 30882 19806
rect 30830 19730 30882 19742
rect 35086 19794 35138 19806
rect 35086 19730 35138 19742
rect 1344 19626 42560 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 42560 19626
rect 1344 19540 42560 19574
rect 4050 19294 4062 19346
rect 4114 19294 4126 19346
rect 7298 19294 7310 19346
rect 7362 19294 7374 19346
rect 26114 19294 26126 19346
rect 26178 19294 26190 19346
rect 33954 19294 33966 19346
rect 34018 19294 34030 19346
rect 37986 19294 37998 19346
rect 38050 19294 38062 19346
rect 12462 19234 12514 19246
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 12462 19170 12514 19182
rect 13582 19234 13634 19246
rect 20862 19234 20914 19246
rect 13906 19182 13918 19234
rect 13970 19182 13982 19234
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 13582 19170 13634 19182
rect 20862 19170 20914 19182
rect 21198 19234 21250 19246
rect 33070 19234 33122 19246
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 32162 19182 32174 19234
rect 32226 19182 32238 19234
rect 32610 19182 32622 19234
rect 32674 19182 32686 19234
rect 21198 19170 21250 19182
rect 33070 19170 33122 19182
rect 24110 19122 24162 19134
rect 3042 19070 3054 19122
rect 3106 19070 3118 19122
rect 6178 19070 6190 19122
rect 6242 19070 6254 19122
rect 24110 19058 24162 19070
rect 24894 19122 24946 19134
rect 27122 19070 27134 19122
rect 27186 19070 27198 19122
rect 34962 19070 34974 19122
rect 35026 19070 35038 19122
rect 38994 19070 39006 19122
rect 39058 19070 39070 19122
rect 24894 19058 24946 19070
rect 8766 19010 8818 19022
rect 12798 19010 12850 19022
rect 17054 19010 17106 19022
rect 9314 18958 9326 19010
rect 9378 18958 9390 19010
rect 16370 18958 16382 19010
rect 16434 18958 16446 19010
rect 8766 18946 8818 18958
rect 12798 18946 12850 18958
rect 17054 18946 17106 18958
rect 17166 19010 17218 19022
rect 25790 19010 25842 19022
rect 17826 18958 17838 19010
rect 17890 18958 17902 19010
rect 17166 18946 17218 18958
rect 25790 18946 25842 18958
rect 29038 19010 29090 19022
rect 29810 18958 29822 19010
rect 29874 18958 29886 19010
rect 29038 18946 29090 18958
rect 1344 18842 42560 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 42560 18842
rect 1344 18756 42560 18790
rect 3054 18674 3106 18686
rect 8878 18674 8930 18686
rect 3826 18622 3838 18674
rect 3890 18622 3902 18674
rect 13234 18622 13246 18674
rect 13298 18622 13310 18674
rect 3054 18610 3106 18622
rect 8878 18610 8930 18622
rect 10322 18510 10334 18562
rect 10386 18510 10398 18562
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 24546 18510 24558 18562
rect 24610 18510 24622 18562
rect 27234 18510 27246 18562
rect 27298 18510 27310 18562
rect 6526 18450 6578 18462
rect 16270 18450 16322 18462
rect 2370 18398 2382 18450
rect 2434 18398 2446 18450
rect 6066 18398 6078 18450
rect 6130 18398 6142 18450
rect 7522 18398 7534 18450
rect 7586 18398 7598 18450
rect 8978 18398 8990 18450
rect 9042 18398 9054 18450
rect 15586 18398 15598 18450
rect 15650 18398 15662 18450
rect 6526 18386 6578 18398
rect 16270 18386 16322 18398
rect 17614 18450 17666 18462
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 19058 18398 19070 18450
rect 19122 18398 19134 18450
rect 26338 18398 26350 18450
rect 26402 18398 26414 18450
rect 30706 18398 30718 18450
rect 30770 18398 30782 18450
rect 33506 18398 33518 18450
rect 33570 18398 33582 18450
rect 38658 18398 38670 18450
rect 38722 18398 38734 18450
rect 17614 18386 17666 18398
rect 16606 18338 16658 18350
rect 2258 18286 2270 18338
rect 2322 18286 2334 18338
rect 7746 18286 7758 18338
rect 7810 18286 7822 18338
rect 11330 18286 11342 18338
rect 11394 18286 11406 18338
rect 16606 18274 16658 18286
rect 17950 18338 18002 18350
rect 39902 18338 39954 18350
rect 20738 18286 20750 18338
rect 20802 18286 20814 18338
rect 23202 18286 23214 18338
rect 23266 18286 23278 18338
rect 35298 18286 35310 18338
rect 35362 18286 35374 18338
rect 38770 18286 38782 18338
rect 38834 18286 38846 18338
rect 17950 18274 18002 18286
rect 39902 18274 39954 18286
rect 12574 18226 12626 18238
rect 12574 18162 12626 18174
rect 26238 18226 26290 18238
rect 26238 18162 26290 18174
rect 1344 18058 42560 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 42560 18058
rect 1344 17972 42560 18006
rect 13022 17890 13074 17902
rect 13022 17826 13074 17838
rect 14030 17890 14082 17902
rect 14030 17826 14082 17838
rect 6302 17778 6354 17790
rect 20750 17778 20802 17790
rect 3490 17726 3502 17778
rect 3554 17726 3566 17778
rect 8082 17726 8094 17778
rect 8146 17726 8158 17778
rect 16818 17726 16830 17778
rect 16882 17726 16894 17778
rect 6302 17714 6354 17726
rect 20750 17714 20802 17726
rect 22878 17778 22930 17790
rect 33518 17778 33570 17790
rect 32498 17726 32510 17778
rect 32562 17726 32574 17778
rect 22878 17714 22930 17726
rect 33518 17714 33570 17726
rect 34638 17778 34690 17790
rect 37986 17726 37998 17778
rect 38050 17726 38062 17778
rect 34638 17714 34690 17726
rect 9550 17666 9602 17678
rect 28590 17666 28642 17678
rect 41022 17666 41074 17678
rect 2370 17614 2382 17666
rect 2434 17614 2446 17666
rect 3378 17614 3390 17666
rect 3442 17614 3454 17666
rect 4722 17614 4734 17666
rect 4786 17614 4798 17666
rect 9874 17614 9886 17666
rect 9938 17614 9950 17666
rect 13906 17614 13918 17666
rect 13970 17614 13982 17666
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 29138 17614 29150 17666
rect 29202 17614 29214 17666
rect 35410 17614 35422 17666
rect 35474 17614 35486 17666
rect 39778 17614 39790 17666
rect 39842 17614 39854 17666
rect 9550 17602 9602 17614
rect 28590 17602 28642 17614
rect 41022 17602 41074 17614
rect 7074 17502 7086 17554
rect 7138 17502 7150 17554
rect 38994 17502 39006 17554
rect 39058 17502 39070 17554
rect 2158 17442 2210 17454
rect 2158 17378 2210 17390
rect 4958 17442 5010 17454
rect 13582 17442 13634 17454
rect 12450 17390 12462 17442
rect 12514 17390 12526 17442
rect 4958 17378 5010 17390
rect 13582 17378 13634 17390
rect 26910 17442 26962 17454
rect 26910 17378 26962 17390
rect 27582 17442 27634 17454
rect 27582 17378 27634 17390
rect 35646 17442 35698 17454
rect 35646 17378 35698 17390
rect 39902 17442 39954 17454
rect 39902 17378 39954 17390
rect 1344 17274 42560 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 42560 17274
rect 1344 17188 42560 17222
rect 5630 17106 5682 17118
rect 2146 17054 2158 17106
rect 2210 17054 2222 17106
rect 28018 17054 28030 17106
rect 28082 17054 28094 17106
rect 36082 17054 36094 17106
rect 36146 17054 36158 17106
rect 5630 17042 5682 17054
rect 22094 16994 22146 17006
rect 8866 16942 8878 16994
rect 8930 16942 8942 16994
rect 10546 16942 10558 16994
rect 10610 16942 10622 16994
rect 22094 16930 22146 16942
rect 28814 16994 28866 17006
rect 31042 16942 31054 16994
rect 31106 16942 31118 16994
rect 39554 16942 39566 16994
rect 39618 16942 39630 16994
rect 28814 16930 28866 16942
rect 5294 16882 5346 16894
rect 18958 16882 19010 16894
rect 4722 16830 4734 16882
rect 4786 16830 4798 16882
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 5294 16818 5346 16830
rect 18958 16818 19010 16830
rect 19406 16882 19458 16894
rect 25342 16882 25394 16894
rect 33182 16882 33234 16894
rect 37214 16882 37266 16894
rect 19730 16830 19742 16882
rect 19794 16830 19806 16882
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 33842 16830 33854 16882
rect 33906 16830 33918 16882
rect 19406 16818 19458 16830
rect 25342 16818 25394 16830
rect 33182 16818 33234 16830
rect 37214 16818 37266 16830
rect 37662 16882 37714 16894
rect 37662 16818 37714 16830
rect 15934 16770 15986 16782
rect 7522 16718 7534 16770
rect 7586 16718 7598 16770
rect 30034 16718 30046 16770
rect 30098 16718 30110 16770
rect 38546 16718 38558 16770
rect 38610 16718 38622 16770
rect 15934 16706 15986 16718
rect 1598 16658 1650 16670
rect 1598 16594 1650 16606
rect 22878 16658 22930 16670
rect 22878 16594 22930 16606
rect 36878 16658 36930 16670
rect 36878 16594 36930 16606
rect 1344 16490 42560 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 42560 16490
rect 1344 16404 42560 16438
rect 13582 16322 13634 16334
rect 13582 16258 13634 16270
rect 21982 16322 22034 16334
rect 21982 16258 22034 16270
rect 30382 16322 30434 16334
rect 30382 16258 30434 16270
rect 36430 16210 36482 16222
rect 4050 16158 4062 16210
rect 4114 16158 4126 16210
rect 11778 16158 11790 16210
rect 11842 16158 11854 16210
rect 18386 16158 18398 16210
rect 18450 16158 18462 16210
rect 29698 16158 29710 16210
rect 29762 16158 29774 16210
rect 36430 16146 36482 16158
rect 9214 16098 9266 16110
rect 23550 16098 23602 16110
rect 31502 16098 31554 16110
rect 40574 16098 40626 16110
rect 8530 16046 8542 16098
rect 8594 16046 8606 16098
rect 13794 16046 13806 16098
rect 13858 16046 13870 16098
rect 16146 16046 16158 16098
rect 16210 16046 16222 16098
rect 22082 16046 22094 16098
rect 22146 16046 22158 16098
rect 23986 16046 23998 16098
rect 24050 16046 24062 16098
rect 29922 16046 29934 16098
rect 29986 16046 29998 16098
rect 30258 16046 30270 16098
rect 30322 16046 30334 16098
rect 31938 16046 31950 16098
rect 32002 16046 32014 16098
rect 35522 16046 35534 16098
rect 35586 16046 35598 16098
rect 40114 16046 40126 16098
rect 40178 16046 40190 16098
rect 9214 16034 9266 16046
rect 23550 16034 23602 16046
rect 31502 16034 31554 16046
rect 40574 16034 40626 16046
rect 5518 15986 5570 15998
rect 26238 15986 26290 15998
rect 3042 15934 3054 15986
rect 3106 15934 3118 15986
rect 10546 15934 10558 15986
rect 10610 15934 10622 15986
rect 5518 15922 5570 15934
rect 26238 15922 26290 15934
rect 37886 15986 37938 15998
rect 37886 15922 37938 15934
rect 9550 15874 9602 15886
rect 6066 15822 6078 15874
rect 6130 15822 6142 15874
rect 9550 15810 9602 15822
rect 20526 15874 20578 15886
rect 20526 15810 20578 15822
rect 27022 15874 27074 15886
rect 27022 15810 27074 15822
rect 28590 15874 28642 15886
rect 34974 15874 35026 15886
rect 34402 15822 34414 15874
rect 34466 15822 34478 15874
rect 28590 15810 28642 15822
rect 34974 15810 35026 15822
rect 35310 15874 35362 15886
rect 35310 15810 35362 15822
rect 37102 15874 37154 15886
rect 37102 15810 37154 15822
rect 1344 15706 42560 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 42560 15706
rect 1344 15620 42560 15654
rect 13246 15538 13298 15550
rect 7410 15486 7422 15538
rect 7474 15486 7486 15538
rect 13246 15474 13298 15486
rect 35982 15538 36034 15550
rect 35982 15474 36034 15486
rect 36542 15538 36594 15550
rect 36542 15474 36594 15486
rect 21310 15426 21362 15438
rect 39678 15426 39730 15438
rect 1922 15374 1934 15426
rect 1986 15374 1998 15426
rect 19394 15374 19406 15426
rect 19458 15374 19470 15426
rect 28690 15374 28702 15426
rect 28754 15374 28766 15426
rect 32050 15374 32062 15426
rect 32114 15374 32126 15426
rect 35074 15374 35086 15426
rect 35138 15374 35150 15426
rect 21310 15362 21362 15374
rect 39678 15362 39730 15374
rect 4734 15314 4786 15326
rect 15598 15314 15650 15326
rect 24222 15314 24274 15326
rect 5058 15262 5070 15314
rect 5122 15262 5134 15314
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 16706 15262 16718 15314
rect 16770 15262 16782 15314
rect 23650 15262 23662 15314
rect 23714 15262 23726 15314
rect 4734 15250 4786 15262
rect 15598 15250 15650 15262
rect 24222 15250 24274 15262
rect 29934 15314 29986 15326
rect 29934 15250 29986 15262
rect 36766 15314 36818 15326
rect 37426 15262 37438 15314
rect 37490 15262 37502 15314
rect 36766 15250 36818 15262
rect 8542 15202 8594 15214
rect 20526 15202 20578 15214
rect 3266 15150 3278 15202
rect 3330 15150 3342 15202
rect 18386 15150 18398 15202
rect 18450 15150 18462 15202
rect 27570 15150 27582 15202
rect 27634 15150 27646 15202
rect 30706 15150 30718 15202
rect 30770 15150 30782 15202
rect 34066 15150 34078 15202
rect 34130 15150 34142 15202
rect 8542 15138 8594 15150
rect 20526 15138 20578 15150
rect 8206 15090 8258 15102
rect 8206 15026 8258 15038
rect 16718 15090 16770 15102
rect 16718 15026 16770 15038
rect 40462 15090 40514 15102
rect 40462 15026 40514 15038
rect 1344 14922 42560 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 42560 14922
rect 1344 14836 42560 14870
rect 22318 14754 22370 14766
rect 22318 14690 22370 14702
rect 20750 14642 20802 14654
rect 3938 14590 3950 14642
rect 4002 14590 4014 14642
rect 11330 14590 11342 14642
rect 11394 14590 11406 14642
rect 20750 14578 20802 14590
rect 21422 14642 21474 14654
rect 24434 14590 24446 14642
rect 24498 14590 24510 14642
rect 29922 14590 29934 14642
rect 29986 14590 29998 14642
rect 34962 14590 34974 14642
rect 35026 14590 35038 14642
rect 21422 14578 21474 14590
rect 6414 14530 6466 14542
rect 15822 14530 15874 14542
rect 32398 14530 32450 14542
rect 40350 14530 40402 14542
rect 7074 14478 7086 14530
rect 7138 14478 7150 14530
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 20290 14478 20302 14530
rect 20354 14478 20366 14530
rect 22194 14478 22206 14530
rect 22258 14478 22270 14530
rect 32722 14478 32734 14530
rect 32786 14478 32798 14530
rect 40002 14478 40014 14530
rect 40066 14478 40078 14530
rect 6414 14466 6466 14478
rect 15822 14466 15874 14478
rect 32398 14466 32450 14478
rect 40350 14466 40402 14478
rect 10110 14418 10162 14430
rect 18510 14418 18562 14430
rect 2706 14366 2718 14418
rect 2770 14366 2782 14418
rect 12338 14366 12350 14418
rect 12402 14366 12414 14418
rect 25442 14366 25454 14418
rect 25506 14366 25518 14418
rect 30930 14366 30942 14418
rect 30994 14366 31006 14418
rect 36306 14366 36318 14418
rect 36370 14366 36382 14418
rect 10110 14354 10162 14366
rect 18510 14354 18562 14366
rect 10446 14306 10498 14318
rect 9538 14254 9550 14306
rect 9602 14254 9614 14306
rect 10446 14242 10498 14254
rect 19294 14306 19346 14318
rect 19294 14242 19346 14254
rect 20190 14306 20242 14318
rect 20190 14242 20242 14254
rect 27246 14306 27298 14318
rect 27246 14242 27298 14254
rect 32846 14306 32898 14318
rect 32846 14242 32898 14254
rect 36878 14306 36930 14318
rect 37650 14254 37662 14306
rect 37714 14254 37726 14306
rect 36878 14242 36930 14254
rect 1344 14138 42560 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 42560 14138
rect 1344 14052 42560 14086
rect 1598 13970 1650 13982
rect 5630 13970 5682 13982
rect 29822 13970 29874 13982
rect 2258 13918 2270 13970
rect 2322 13918 2334 13970
rect 16370 13918 16382 13970
rect 16434 13918 16446 13970
rect 20178 13918 20190 13970
rect 20242 13918 20254 13970
rect 1598 13906 1650 13918
rect 5630 13906 5682 13918
rect 29822 13906 29874 13918
rect 36990 13970 37042 13982
rect 36990 13906 37042 13918
rect 39790 13970 39842 13982
rect 39790 13906 39842 13918
rect 23998 13858 24050 13870
rect 8530 13806 8542 13858
rect 8594 13806 8606 13858
rect 10658 13806 10670 13858
rect 10722 13806 10734 13858
rect 23998 13794 24050 13806
rect 29038 13858 29090 13870
rect 35870 13858 35922 13870
rect 32050 13806 32062 13858
rect 32114 13806 32126 13858
rect 37762 13806 37774 13858
rect 37826 13806 37838 13858
rect 29038 13794 29090 13806
rect 35870 13794 35922 13806
rect 17502 13746 17554 13758
rect 21310 13746 21362 13758
rect 26126 13746 26178 13758
rect 33182 13746 33234 13758
rect 4610 13694 4622 13746
rect 4674 13694 4686 13746
rect 5170 13694 5182 13746
rect 5234 13694 5246 13746
rect 13346 13694 13358 13746
rect 13410 13694 13422 13746
rect 13906 13694 13918 13746
rect 13970 13694 13982 13746
rect 17938 13694 17950 13746
rect 18002 13694 18014 13746
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 26786 13694 26798 13746
rect 26850 13694 26862 13746
rect 33618 13694 33630 13746
rect 33682 13694 33694 13746
rect 17502 13682 17554 13694
rect 21310 13682 21362 13694
rect 26126 13682 26178 13694
rect 33182 13682 33234 13694
rect 7522 13582 7534 13634
rect 7586 13582 7598 13634
rect 12002 13582 12014 13634
rect 12066 13582 12078 13634
rect 31042 13582 31054 13634
rect 31106 13582 31118 13634
rect 38882 13582 38894 13634
rect 38946 13582 38958 13634
rect 16942 13522 16994 13534
rect 16942 13458 16994 13470
rect 20974 13522 21026 13534
rect 20974 13458 21026 13470
rect 24782 13522 24834 13534
rect 24782 13458 24834 13470
rect 36654 13522 36706 13534
rect 36654 13458 36706 13470
rect 1344 13354 42560 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 42560 13354
rect 1344 13268 42560 13302
rect 4174 13186 4226 13198
rect 27358 13186 27410 13198
rect 23202 13134 23214 13186
rect 23266 13134 23278 13186
rect 4174 13122 4226 13134
rect 27358 13122 27410 13134
rect 33070 13074 33122 13086
rect 16482 13022 16494 13074
rect 16546 13022 16558 13074
rect 19506 13022 19518 13074
rect 19570 13022 19582 13074
rect 33070 13010 33122 13022
rect 33518 13074 33570 13086
rect 37102 13074 37154 13086
rect 33954 13022 33966 13074
rect 34018 13022 34030 13074
rect 38322 13022 38334 13074
rect 38386 13022 38398 13074
rect 40338 13022 40350 13074
rect 40402 13022 40414 13074
rect 33518 13010 33570 13022
rect 37102 13010 37154 13022
rect 10670 12962 10722 12974
rect 29262 12962 29314 12974
rect 3938 12910 3950 12962
rect 4002 12910 4014 12962
rect 6962 12910 6974 12962
rect 7026 12910 7038 12962
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 12450 12910 12462 12962
rect 12514 12910 12526 12962
rect 13570 12910 13582 12962
rect 13634 12910 13646 12962
rect 21634 12910 21646 12962
rect 21698 12910 21710 12962
rect 22642 12910 22654 12962
rect 22706 12910 22718 12962
rect 23762 12910 23774 12962
rect 23826 12910 23838 12962
rect 24322 12910 24334 12962
rect 24386 12910 24398 12962
rect 27794 12910 27806 12962
rect 27858 12910 27870 12962
rect 29698 12910 29710 12962
rect 29762 12910 29774 12962
rect 40114 12910 40126 12962
rect 40178 12910 40190 12962
rect 10670 12898 10722 12910
rect 29262 12898 29314 12910
rect 32734 12850 32786 12862
rect 17490 12798 17502 12850
rect 17554 12798 17566 12850
rect 20626 12798 20638 12850
rect 20690 12798 20702 12850
rect 21522 12798 21534 12850
rect 21586 12798 21598 12850
rect 34962 12798 34974 12850
rect 35026 12798 35038 12850
rect 39330 12798 39342 12850
rect 39394 12798 39406 12850
rect 32734 12786 32786 12798
rect 6862 12738 6914 12750
rect 6862 12674 6914 12686
rect 7198 12738 7250 12750
rect 11230 12738 11282 12750
rect 7746 12686 7758 12738
rect 7810 12686 7822 12738
rect 7198 12674 7250 12686
rect 11230 12674 11282 12686
rect 12238 12738 12290 12750
rect 16158 12738 16210 12750
rect 27694 12738 27746 12750
rect 14130 12686 14142 12738
rect 14194 12686 14206 12738
rect 26786 12686 26798 12738
rect 26850 12686 26862 12738
rect 32162 12686 32174 12738
rect 32226 12686 32238 12738
rect 12238 12674 12290 12686
rect 16158 12674 16210 12686
rect 27694 12674 27746 12686
rect 1344 12570 42560 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 42560 12570
rect 1344 12484 42560 12518
rect 9662 12402 9714 12414
rect 17502 12402 17554 12414
rect 14914 12350 14926 12402
rect 14978 12350 14990 12402
rect 9662 12338 9714 12350
rect 17502 12338 17554 12350
rect 17950 12402 18002 12414
rect 38110 12402 38162 12414
rect 29474 12350 29486 12402
rect 29538 12350 29550 12402
rect 33282 12350 33294 12402
rect 33346 12350 33358 12402
rect 37090 12350 37102 12402
rect 37154 12350 37166 12402
rect 17950 12338 18002 12350
rect 38110 12338 38162 12350
rect 39342 12402 39394 12414
rect 39342 12338 39394 12350
rect 8318 12290 8370 12302
rect 21198 12290 21250 12302
rect 19730 12238 19742 12290
rect 19794 12238 19806 12290
rect 8318 12226 8370 12238
rect 21198 12226 21250 12238
rect 25902 12290 25954 12302
rect 25902 12226 25954 12238
rect 5630 12178 5682 12190
rect 12238 12178 12290 12190
rect 23886 12178 23938 12190
rect 28590 12178 28642 12190
rect 32622 12178 32674 12190
rect 34078 12178 34130 12190
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 9874 12126 9886 12178
rect 9938 12126 9950 12178
rect 11778 12126 11790 12178
rect 11842 12126 11854 12178
rect 12562 12126 12574 12178
rect 12626 12126 12638 12178
rect 16706 12126 16718 12178
rect 16770 12126 16782 12178
rect 23426 12126 23438 12178
rect 23490 12126 23502 12178
rect 28242 12126 28254 12178
rect 28306 12126 28318 12178
rect 32050 12126 32062 12178
rect 32114 12126 32126 12178
rect 33506 12126 33518 12178
rect 33570 12126 33582 12178
rect 34738 12126 34750 12178
rect 34802 12126 34814 12178
rect 39218 12126 39230 12178
rect 39282 12126 39294 12178
rect 5630 12114 5682 12126
rect 12238 12114 12290 12126
rect 23886 12114 23938 12126
rect 28590 12114 28642 12126
rect 32622 12114 32674 12126
rect 34078 12114 34130 12126
rect 18722 12014 18734 12066
rect 18786 12014 18798 12066
rect 9102 11954 9154 11966
rect 9102 11890 9154 11902
rect 11678 11954 11730 11966
rect 11678 11890 11730 11902
rect 15710 11954 15762 11966
rect 15710 11890 15762 11902
rect 16718 11954 16770 11966
rect 16718 11890 16770 11902
rect 20414 11954 20466 11966
rect 20414 11890 20466 11902
rect 25118 11954 25170 11966
rect 25118 11890 25170 11902
rect 28926 11954 28978 11966
rect 28926 11890 28978 11902
rect 37774 11954 37826 11966
rect 37774 11890 37826 11902
rect 1344 11786 42560 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 42560 11786
rect 1344 11700 42560 11734
rect 9326 11618 9378 11630
rect 9326 11554 9378 11566
rect 27582 11618 27634 11630
rect 27582 11554 27634 11566
rect 37102 11618 37154 11630
rect 37102 11554 37154 11566
rect 36542 11506 36594 11518
rect 7634 11454 7646 11506
rect 7698 11454 7710 11506
rect 14914 11454 14926 11506
rect 14978 11454 14990 11506
rect 22306 11454 22318 11506
rect 22370 11454 22382 11506
rect 25666 11454 25678 11506
rect 25730 11454 25742 11506
rect 33954 11454 33966 11506
rect 34018 11454 34030 11506
rect 36542 11442 36594 11454
rect 38446 11506 38498 11518
rect 40674 11454 40686 11506
rect 40738 11454 40750 11506
rect 38446 11442 38498 11454
rect 13022 11394 13074 11406
rect 20078 11394 20130 11406
rect 30046 11394 30098 11406
rect 12338 11342 12350 11394
rect 12402 11342 12414 11394
rect 19618 11342 19630 11394
rect 19682 11342 19694 11394
rect 27570 11342 27582 11394
rect 27634 11342 27646 11394
rect 30706 11342 30718 11394
rect 30770 11342 30782 11394
rect 36978 11342 36990 11394
rect 37042 11342 37054 11394
rect 13022 11330 13074 11342
rect 20078 11330 20130 11342
rect 30046 11330 30098 11342
rect 10110 11282 10162 11294
rect 8642 11230 8654 11282
rect 8706 11230 8718 11282
rect 15922 11230 15934 11282
rect 15986 11230 15998 11282
rect 23538 11230 23550 11282
rect 23602 11230 23614 11282
rect 27010 11230 27022 11282
rect 27074 11230 27086 11282
rect 34962 11230 34974 11282
rect 35026 11230 35038 11282
rect 41682 11230 41694 11282
rect 41746 11230 41758 11282
rect 10110 11218 10162 11230
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 14590 11170 14642 11182
rect 14590 11106 14642 11118
rect 16606 11170 16658 11182
rect 33742 11170 33794 11182
rect 17154 11118 17166 11170
rect 17218 11118 17230 11170
rect 33170 11118 33182 11170
rect 33234 11118 33246 11170
rect 16606 11106 16658 11118
rect 33742 11106 33794 11118
rect 1344 11002 42560 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 42560 11002
rect 1344 10916 42560 10950
rect 8318 10834 8370 10846
rect 8318 10770 8370 10782
rect 16494 10834 16546 10846
rect 16494 10770 16546 10782
rect 17502 10834 17554 10846
rect 22654 10834 22706 10846
rect 21522 10782 21534 10834
rect 21586 10782 21598 10834
rect 17502 10770 17554 10782
rect 22654 10770 22706 10782
rect 32622 10834 32674 10846
rect 32622 10770 32674 10782
rect 33182 10834 33234 10846
rect 33182 10770 33234 10782
rect 34414 10834 34466 10846
rect 34414 10770 34466 10782
rect 15374 10722 15426 10734
rect 11554 10670 11566 10722
rect 11618 10670 11630 10722
rect 26226 10670 26238 10722
rect 26290 10670 26302 10722
rect 30034 10670 30046 10722
rect 30098 10670 30110 10722
rect 37874 10670 37886 10722
rect 37938 10670 37950 10722
rect 15374 10658 15426 10670
rect 12686 10610 12738 10622
rect 18622 10610 18674 10622
rect 8530 10558 8542 10610
rect 8594 10558 8606 10610
rect 13122 10558 13134 10610
rect 13186 10558 13198 10610
rect 17714 10558 17726 10610
rect 17778 10558 17790 10610
rect 19282 10558 19294 10610
rect 19346 10558 19358 10610
rect 22530 10558 22542 10610
rect 22594 10558 22606 10610
rect 33058 10558 33070 10610
rect 33122 10558 33134 10610
rect 12686 10546 12738 10558
rect 18622 10546 18674 10558
rect 9662 10498 9714 10510
rect 28030 10498 28082 10510
rect 32062 10498 32114 10510
rect 10546 10446 10558 10498
rect 10610 10446 10622 10498
rect 27346 10446 27358 10498
rect 27410 10446 27422 10498
rect 31154 10446 31166 10498
rect 31218 10446 31230 10498
rect 36866 10446 36878 10498
rect 36930 10446 36942 10498
rect 9662 10434 9714 10446
rect 28030 10434 28082 10446
rect 32062 10434 32114 10446
rect 16158 10386 16210 10398
rect 16158 10322 16210 10334
rect 22318 10386 22370 10398
rect 22318 10322 22370 10334
rect 1344 10218 42560 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 42560 10218
rect 1344 10132 42560 10166
rect 28478 10050 28530 10062
rect 14354 9998 14366 10050
rect 14418 9998 14430 10050
rect 28478 9986 28530 9998
rect 18958 9938 19010 9950
rect 18958 9874 19010 9886
rect 19406 9938 19458 9950
rect 24322 9886 24334 9938
rect 24386 9886 24398 9938
rect 30034 9886 30046 9938
rect 30098 9886 30110 9938
rect 40226 9886 40238 9938
rect 40290 9886 40302 9938
rect 19406 9874 19458 9886
rect 9550 9826 9602 9838
rect 15038 9826 15090 9838
rect 27582 9826 27634 9838
rect 29486 9826 29538 9838
rect 2930 9774 2942 9826
rect 2994 9774 3006 9826
rect 9986 9774 9998 9826
rect 10050 9774 10062 9826
rect 13794 9774 13806 9826
rect 13858 9774 13870 9826
rect 15474 9774 15486 9826
rect 15538 9774 15550 9826
rect 28578 9774 28590 9826
rect 28642 9774 28654 9826
rect 30482 9774 30494 9826
rect 30546 9774 30558 9826
rect 9550 9762 9602 9774
rect 15038 9762 15090 9774
rect 27582 9762 27634 9774
rect 29486 9762 29538 9774
rect 12238 9714 12290 9726
rect 2034 9662 2046 9714
rect 2098 9662 2110 9714
rect 23202 9662 23214 9714
rect 23266 9662 23278 9714
rect 39106 9662 39118 9714
rect 39170 9662 39182 9714
rect 12238 9650 12290 9662
rect 13022 9602 13074 9614
rect 18510 9602 18562 9614
rect 17714 9550 17726 9602
rect 17778 9550 17790 9602
rect 13022 9538 13074 9550
rect 18510 9538 18562 9550
rect 1344 9434 42560 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 42560 9434
rect 1344 9348 42560 9382
rect 13010 9102 13022 9154
rect 13074 9102 13086 9154
rect 16706 9102 16718 9154
rect 16770 9102 16782 9154
rect 17714 9102 17726 9154
rect 17778 9102 17790 9154
rect 21970 9102 21982 9154
rect 22034 9102 22046 9154
rect 2930 8990 2942 9042
rect 2994 8990 3006 9042
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 17826 8990 17838 9042
rect 17890 8990 17902 9042
rect 13918 8930 13970 8942
rect 1922 8878 1934 8930
rect 1986 8878 1998 8930
rect 12002 8878 12014 8930
rect 12066 8878 12078 8930
rect 15362 8878 15374 8930
rect 15426 8878 15438 8930
rect 20962 8878 20974 8930
rect 21026 8878 21038 8930
rect 13918 8866 13970 8878
rect 10334 8818 10386 8830
rect 10334 8754 10386 8766
rect 1344 8650 42560 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 42560 8650
rect 1344 8564 42560 8598
rect 11678 8370 11730 8382
rect 11678 8306 11730 8318
rect 12126 8370 12178 8382
rect 16258 8318 16270 8370
rect 16322 8318 16334 8370
rect 19506 8318 19518 8370
rect 19570 8318 19582 8370
rect 12126 8306 12178 8318
rect 8206 8258 8258 8270
rect 2706 8206 2718 8258
rect 2770 8206 2782 8258
rect 8642 8206 8654 8258
rect 8706 8206 8718 8258
rect 8206 8194 8258 8206
rect 10894 8146 10946 8158
rect 2034 8094 2046 8146
rect 2098 8094 2110 8146
rect 17266 8094 17278 8146
rect 17330 8094 17342 8146
rect 18386 8094 18398 8146
rect 18450 8094 18462 8146
rect 10894 8082 10946 8094
rect 3278 8034 3330 8046
rect 3278 7970 3330 7982
rect 1344 7866 42560 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 42560 7866
rect 1344 7780 42560 7814
rect 14242 7534 14254 7586
rect 14306 7534 14318 7586
rect 2930 7422 2942 7474
rect 2994 7422 3006 7474
rect 1922 7310 1934 7362
rect 1986 7310 1998 7362
rect 13234 7310 13246 7362
rect 13298 7310 13310 7362
rect 1344 7082 42560 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 42560 7082
rect 1344 6996 42560 7030
rect 2818 6638 2830 6690
rect 2882 6638 2894 6690
rect 2034 6526 2046 6578
rect 2098 6526 2110 6578
rect 1344 6298 42560 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 42560 6298
rect 1344 6212 42560 6246
rect 3278 6130 3330 6142
rect 3278 6066 3330 6078
rect 2706 5854 2718 5906
rect 2770 5854 2782 5906
rect 3490 5854 3502 5906
rect 3554 5854 3566 5906
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 1344 5514 42560 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 42560 5514
rect 1344 5428 42560 5462
rect 6974 5122 7026 5134
rect 3826 5070 3838 5122
rect 3890 5070 3902 5122
rect 4498 5070 4510 5122
rect 4562 5070 4574 5122
rect 10434 5070 10446 5122
rect 10498 5070 10510 5122
rect 6974 5058 7026 5070
rect 2270 5010 2322 5022
rect 2270 4946 2322 4958
rect 2606 5010 2658 5022
rect 2606 4946 2658 4958
rect 2942 5010 2994 5022
rect 2942 4946 2994 4958
rect 3278 5010 3330 5022
rect 3278 4946 3330 4958
rect 3614 5010 3666 5022
rect 3614 4946 3666 4958
rect 4286 5010 4338 5022
rect 4286 4946 4338 4958
rect 1710 4898 1762 4910
rect 1710 4834 1762 4846
rect 7310 4898 7362 4910
rect 7310 4834 7362 4846
rect 10670 4898 10722 4910
rect 10670 4834 10722 4846
rect 1344 4730 42560 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 42560 4730
rect 1344 4644 42560 4678
rect 2046 4562 2098 4574
rect 2046 4498 2098 4510
rect 2942 4562 2994 4574
rect 2942 4498 2994 4510
rect 3614 4562 3666 4574
rect 3614 4498 3666 4510
rect 1710 4450 1762 4462
rect 1710 4386 1762 4398
rect 2382 4450 2434 4462
rect 2382 4386 2434 4398
rect 3278 4450 3330 4462
rect 3278 4386 3330 4398
rect 4846 4450 4898 4462
rect 4846 4386 4898 4398
rect 3826 4286 3838 4338
rect 3890 4286 3902 4338
rect 4398 4226 4450 4238
rect 4398 4162 4450 4174
rect 5294 4226 5346 4238
rect 5294 4162 5346 4174
rect 5742 4226 5794 4238
rect 5742 4162 5794 4174
rect 1344 3946 42560 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 42560 3946
rect 1344 3860 42560 3894
rect 7970 3614 7982 3666
rect 8034 3614 8046 3666
rect 11442 3614 11454 3666
rect 11506 3614 11518 3666
rect 1710 3554 1762 3566
rect 7534 3554 7586 3566
rect 3938 3502 3950 3554
rect 4002 3502 4014 3554
rect 1710 3490 1762 3502
rect 7534 3490 7586 3502
rect 11006 3554 11058 3566
rect 11006 3490 11058 3502
rect 2046 3442 2098 3454
rect 2046 3378 2098 3390
rect 2382 3442 2434 3454
rect 2382 3378 2434 3390
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 3054 3442 3106 3454
rect 3054 3378 3106 3390
rect 3390 3442 3442 3454
rect 3390 3378 3442 3390
rect 3726 3442 3778 3454
rect 3726 3378 3778 3390
rect 4510 3442 4562 3454
rect 4510 3378 4562 3390
rect 4958 3442 5010 3454
rect 4958 3378 5010 3390
rect 6078 3442 6130 3454
rect 6078 3378 6130 3390
rect 6302 3442 6354 3454
rect 6302 3378 6354 3390
rect 6638 3442 6690 3454
rect 6638 3378 6690 3390
rect 10110 3442 10162 3454
rect 10110 3378 10162 3390
rect 10334 3442 10386 3454
rect 10334 3378 10386 3390
rect 10670 3442 10722 3454
rect 10670 3378 10722 3390
rect 6974 3330 7026 3342
rect 6974 3266 7026 3278
rect 9326 3330 9378 3342
rect 9326 3266 9378 3278
rect 13134 3330 13186 3342
rect 13134 3266 13186 3278
rect 1344 3162 42560 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 42560 3162
rect 1344 3076 42560 3110
rect 12114 1710 12126 1762
rect 12178 1759 12190 1762
rect 13122 1759 13134 1762
rect 12178 1713 13134 1759
rect 12178 1710 12190 1713
rect 13122 1710 13134 1713
rect 13186 1710 13198 1762
<< via1 >>
rect 10110 41806 10162 41858
rect 11230 41806 11282 41858
rect 15486 41246 15538 41298
rect 16046 41246 16098 41298
rect 5406 41022 5458 41074
rect 5966 41022 6018 41074
rect 22206 41022 22258 41074
rect 23326 41022 23378 41074
rect 20190 40910 20242 40962
rect 20862 40910 20914 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 1822 40574 1874 40626
rect 11902 40574 11954 40626
rect 12350 40574 12402 40626
rect 13134 40574 13186 40626
rect 13694 40574 13746 40626
rect 14254 40574 14306 40626
rect 14814 40574 14866 40626
rect 17726 40574 17778 40626
rect 19182 40574 19234 40626
rect 19854 40574 19906 40626
rect 20190 40574 20242 40626
rect 4062 40462 4114 40514
rect 5966 40462 6018 40514
rect 7870 40462 7922 40514
rect 9326 40462 9378 40514
rect 11230 40462 11282 40514
rect 16046 40462 16098 40514
rect 17054 40462 17106 40514
rect 20750 40462 20802 40514
rect 21758 40462 21810 40514
rect 23326 40462 23378 40514
rect 3278 40350 3330 40402
rect 4958 40350 5010 40402
rect 6638 40350 6690 40402
rect 8766 40350 8818 40402
rect 9550 40350 9602 40402
rect 10334 40350 10386 40402
rect 15150 40350 15202 40402
rect 17278 40350 17330 40402
rect 18510 40350 18562 40402
rect 20974 40350 21026 40402
rect 21982 40350 22034 40402
rect 22430 40350 22482 40402
rect 24558 40350 24610 40402
rect 25790 40350 25842 40402
rect 26126 40350 26178 40402
rect 2718 40238 2770 40290
rect 25006 40238 25058 40290
rect 26574 40238 26626 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 2494 39790 2546 39842
rect 4062 39790 4114 39842
rect 9438 39678 9490 39730
rect 10222 39678 10274 39730
rect 16830 39678 16882 39730
rect 17614 39678 17666 39730
rect 18846 39678 18898 39730
rect 21534 39678 21586 39730
rect 22878 39678 22930 39730
rect 25566 39678 25618 39730
rect 27582 39678 27634 39730
rect 6974 39566 7026 39618
rect 7870 39566 7922 39618
rect 8430 39566 8482 39618
rect 19294 39566 19346 39618
rect 23998 39566 24050 39618
rect 26014 39566 26066 39618
rect 26686 39566 26738 39618
rect 5630 39454 5682 39506
rect 5966 39454 6018 39506
rect 6638 39454 6690 39506
rect 10558 39454 10610 39506
rect 11006 39454 11058 39506
rect 20414 39454 20466 39506
rect 23102 39454 23154 39506
rect 3278 39342 3330 39394
rect 4846 39342 4898 39394
rect 6302 39342 6354 39394
rect 7310 39342 7362 39394
rect 7646 39342 7698 39394
rect 8654 39342 8706 39394
rect 8990 39342 9042 39394
rect 16382 39342 16434 39394
rect 19070 39342 19122 39394
rect 23774 39342 23826 39394
rect 25790 39342 25842 39394
rect 26462 39342 26514 39394
rect 27134 39342 27186 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 2158 39006 2210 39058
rect 3726 39006 3778 39058
rect 5518 39006 5570 39058
rect 6862 39006 6914 39058
rect 7534 39006 7586 39058
rect 8654 39006 8706 39058
rect 9662 39006 9714 39058
rect 26238 39006 26290 39058
rect 2942 38894 2994 38946
rect 4846 38894 4898 38946
rect 6190 38894 6242 38946
rect 8318 38894 8370 38946
rect 4398 38782 4450 38834
rect 5070 38782 5122 38834
rect 5742 38782 5794 38834
rect 6526 38782 6578 38834
rect 7198 38782 7250 38834
rect 8094 38782 8146 38834
rect 8878 38782 8930 38834
rect 1822 38670 1874 38722
rect 10222 38670 10274 38722
rect 26798 38670 26850 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 2158 38222 2210 38274
rect 7086 37998 7138 38050
rect 8318 37998 8370 38050
rect 9102 37998 9154 38050
rect 9774 37998 9826 38050
rect 10670 37998 10722 38050
rect 3614 37886 3666 37938
rect 3950 37886 4002 37938
rect 4734 37886 4786 37938
rect 5966 37886 6018 37938
rect 6302 37886 6354 37938
rect 6638 37886 6690 37938
rect 7310 37886 7362 37938
rect 7646 37886 7698 37938
rect 7982 37886 8034 37938
rect 9326 37886 9378 37938
rect 9998 37886 10050 37938
rect 10334 37886 10386 37938
rect 1934 37774 1986 37826
rect 2942 37774 2994 37826
rect 3278 37774 3330 37826
rect 4398 37774 4450 37826
rect 5630 37774 5682 37826
rect 8654 37774 8706 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 2158 37438 2210 37490
rect 2942 37438 2994 37490
rect 4622 37438 4674 37490
rect 5294 37438 5346 37490
rect 6302 37438 6354 37490
rect 6974 37438 7026 37490
rect 7422 37438 7474 37490
rect 8430 37438 8482 37490
rect 3278 37326 3330 37378
rect 3950 37326 4002 37378
rect 4958 37326 5010 37378
rect 3614 37214 3666 37266
rect 4286 37214 4338 37266
rect 5518 37214 5570 37266
rect 8206 37214 8258 37266
rect 1822 37102 1874 37154
rect 8990 37102 9042 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 5742 36542 5794 36594
rect 40686 36542 40738 36594
rect 1710 36430 1762 36482
rect 3278 36430 3330 36482
rect 4398 36430 4450 36482
rect 2046 36318 2098 36370
rect 2382 36318 2434 36370
rect 2718 36318 2770 36370
rect 4062 36318 4114 36370
rect 4734 36318 4786 36370
rect 41694 36318 41746 36370
rect 3054 36206 3106 36258
rect 3726 36206 3778 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 2046 35870 2098 35922
rect 2942 35870 2994 35922
rect 3950 35870 4002 35922
rect 4398 35870 4450 35922
rect 2382 35758 2434 35810
rect 3278 35758 3330 35810
rect 3614 35758 3666 35810
rect 1710 35646 1762 35698
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 3614 35086 3666 35138
rect 3838 35086 3890 35138
rect 3838 34974 3890 35026
rect 40350 34974 40402 35026
rect 2718 34862 2770 34914
rect 2046 34750 2098 34802
rect 3278 34750 3330 34802
rect 39118 34750 39170 34802
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2158 34302 2210 34354
rect 1710 34190 1762 34242
rect 16270 34190 16322 34242
rect 19742 34190 19794 34242
rect 27246 34190 27298 34242
rect 35646 34190 35698 34242
rect 37326 34190 37378 34242
rect 15038 33966 15090 34018
rect 18734 33966 18786 34018
rect 26238 33966 26290 34018
rect 34414 33966 34466 34018
rect 38446 33966 38498 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 8766 33406 8818 33458
rect 15150 33406 15202 33458
rect 18398 33406 18450 33458
rect 24558 33406 24610 33458
rect 27134 33406 27186 33458
rect 30158 33406 30210 33458
rect 32958 33406 33010 33458
rect 38446 33406 38498 33458
rect 1710 33182 1762 33234
rect 2046 33182 2098 33234
rect 9774 33182 9826 33234
rect 16158 33182 16210 33234
rect 17054 33182 17106 33234
rect 25678 33182 25730 33234
rect 28142 33182 28194 33234
rect 31166 33182 31218 33234
rect 33966 33182 34018 33234
rect 39454 33182 39506 33234
rect 2494 33070 2546 33122
rect 29374 33070 29426 33122
rect 29822 33070 29874 33122
rect 32734 33070 32786 33122
rect 37214 33070 37266 33122
rect 37662 33070 37714 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 30494 32734 30546 32786
rect 32398 32734 32450 32786
rect 35086 32734 35138 32786
rect 1710 32622 1762 32674
rect 5742 32622 5794 32674
rect 9886 32622 9938 32674
rect 15934 32622 15986 32674
rect 20078 32622 20130 32674
rect 29710 32622 29762 32674
rect 26910 32510 26962 32562
rect 27470 32510 27522 32562
rect 31166 32510 31218 32562
rect 31950 32510 32002 32562
rect 33518 32510 33570 32562
rect 37550 32510 37602 32562
rect 38110 32510 38162 32562
rect 39118 32510 39170 32562
rect 39902 32510 39954 32562
rect 40350 32510 40402 32562
rect 6862 32398 6914 32450
rect 10894 32398 10946 32450
rect 14926 32398 14978 32450
rect 19406 32398 19458 32450
rect 21198 32398 21250 32450
rect 24334 32398 24386 32450
rect 24670 32398 24722 32450
rect 26014 32398 26066 32450
rect 26238 32398 26290 32450
rect 33406 32398 33458 32450
rect 31390 32286 31442 32338
rect 34414 32286 34466 32338
rect 39342 32286 39394 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 27022 31950 27074 32002
rect 8654 31838 8706 31890
rect 11678 31838 11730 31890
rect 19182 31838 19234 31890
rect 36542 31838 36594 31890
rect 37102 31838 37154 31890
rect 40350 31838 40402 31890
rect 2718 31726 2770 31778
rect 15710 31726 15762 31778
rect 16158 31726 16210 31778
rect 20302 31726 20354 31778
rect 23326 31726 23378 31778
rect 23998 31726 24050 31778
rect 28590 31726 28642 31778
rect 29038 31726 29090 31778
rect 29598 31726 29650 31778
rect 33070 31726 33122 31778
rect 33406 31726 33458 31778
rect 37326 31726 37378 31778
rect 38222 31726 38274 31778
rect 2046 31614 2098 31666
rect 9774 31614 9826 31666
rect 12798 31614 12850 31666
rect 19406 31614 19458 31666
rect 19742 31614 19794 31666
rect 26238 31614 26290 31666
rect 39230 31614 39282 31666
rect 8430 31502 8482 31554
rect 11230 31502 11282 31554
rect 14590 31502 14642 31554
rect 18398 31502 18450 31554
rect 20302 31502 20354 31554
rect 21422 31502 21474 31554
rect 27358 31502 27410 31554
rect 28478 31502 28530 31554
rect 31950 31502 32002 31554
rect 32734 31502 32786 31554
rect 35758 31502 35810 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4958 31166 5010 31218
rect 8990 31166 9042 31218
rect 9662 31166 9714 31218
rect 14702 31166 14754 31218
rect 15262 31166 15314 31218
rect 15598 31166 15650 31218
rect 17278 31166 17330 31218
rect 24222 31166 24274 31218
rect 24782 31166 24834 31218
rect 28590 31166 28642 31218
rect 29374 31166 29426 31218
rect 30158 31166 30210 31218
rect 32958 31166 33010 31218
rect 33630 31166 33682 31218
rect 5742 31054 5794 31106
rect 18062 31054 18114 31106
rect 31838 31054 31890 31106
rect 38894 31054 38946 31106
rect 2942 30942 2994 30994
rect 8094 30942 8146 30994
rect 8654 30942 8706 30994
rect 10334 30942 10386 30994
rect 11006 30942 11058 30994
rect 11678 30942 11730 30994
rect 12126 30942 12178 30994
rect 20414 30942 20466 30994
rect 20750 30942 20802 30994
rect 21086 30942 21138 30994
rect 21758 30942 21810 30994
rect 25678 30942 25730 30994
rect 26350 30942 26402 30994
rect 36094 30942 36146 30994
rect 36654 30942 36706 30994
rect 37438 30942 37490 30994
rect 1934 30830 1986 30882
rect 10110 30830 10162 30882
rect 10782 30830 10834 30882
rect 25342 30830 25394 30882
rect 29710 30830 29762 30882
rect 30606 30830 30658 30882
rect 36990 30830 37042 30882
rect 37886 30830 37938 30882
rect 9438 30718 9490 30770
rect 9774 30718 9826 30770
rect 36990 30718 37042 30770
rect 37550 30718 37602 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 29822 30382 29874 30434
rect 27022 30270 27074 30322
rect 35758 30270 35810 30322
rect 2382 30158 2434 30210
rect 3166 30158 3218 30210
rect 7758 30158 7810 30210
rect 8206 30158 8258 30210
rect 11678 30158 11730 30210
rect 12574 30158 12626 30210
rect 13470 30158 13522 30210
rect 14030 30158 14082 30210
rect 17054 30158 17106 30210
rect 17390 30158 17442 30210
rect 17838 30158 17890 30210
rect 21758 30158 21810 30210
rect 22206 30158 22258 30210
rect 22766 30158 22818 30210
rect 29598 30158 29650 30210
rect 30270 30158 30322 30210
rect 33406 30158 33458 30210
rect 33966 30158 34018 30210
rect 34750 30158 34802 30210
rect 35870 30158 35922 30210
rect 36990 30158 37042 30210
rect 37662 30158 37714 30210
rect 40686 30158 40738 30210
rect 40910 30158 40962 30210
rect 1710 30046 1762 30098
rect 2046 30046 2098 30098
rect 2718 30046 2770 30098
rect 11454 30046 11506 30098
rect 12350 30046 12402 30098
rect 21534 30046 21586 30098
rect 25790 30046 25842 30098
rect 28030 30046 28082 30098
rect 39902 30046 39954 30098
rect 3614 29934 3666 29986
rect 10670 29934 10722 29986
rect 11230 29934 11282 29986
rect 16494 29934 16546 29986
rect 20302 29934 20354 29986
rect 20862 29934 20914 29986
rect 25118 29934 25170 29986
rect 26126 29934 26178 29986
rect 31054 29934 31106 29986
rect 34526 29934 34578 29986
rect 41022 29934 41074 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 2046 29598 2098 29650
rect 8318 29598 8370 29650
rect 9102 29598 9154 29650
rect 9662 29598 9714 29650
rect 13694 29598 13746 29650
rect 14366 29598 14418 29650
rect 15038 29598 15090 29650
rect 23550 29598 23602 29650
rect 31390 29598 31442 29650
rect 31838 29598 31890 29650
rect 33854 29598 33906 29650
rect 36094 29598 36146 29650
rect 36766 29598 36818 29650
rect 37550 29598 37602 29650
rect 41022 29598 41074 29650
rect 19406 29486 19458 29538
rect 24334 29486 24386 29538
rect 27246 29486 27298 29538
rect 30270 29486 30322 29538
rect 35310 29486 35362 29538
rect 1710 29374 1762 29426
rect 5630 29374 5682 29426
rect 6078 29374 6130 29426
rect 10334 29374 10386 29426
rect 10670 29374 10722 29426
rect 11342 29374 11394 29426
rect 16606 29374 16658 29426
rect 20526 29374 20578 29426
rect 21086 29374 21138 29426
rect 24110 29374 24162 29426
rect 31726 29374 31778 29426
rect 39902 29374 39954 29426
rect 40462 29374 40514 29426
rect 2494 29262 2546 29314
rect 10110 29262 10162 29314
rect 14926 29262 14978 29314
rect 17502 29262 17554 29314
rect 17950 29262 18002 29314
rect 18398 29262 18450 29314
rect 24670 29262 24722 29314
rect 25342 29262 25394 29314
rect 26238 29262 26290 29314
rect 28142 29262 28194 29314
rect 29038 29262 29090 29314
rect 33406 29262 33458 29314
rect 34190 29262 34242 29314
rect 36542 29262 36594 29314
rect 15822 29150 15874 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 9214 28814 9266 28866
rect 13022 28814 13074 28866
rect 15934 28814 15986 28866
rect 36878 28814 36930 28866
rect 13694 28702 13746 28754
rect 19854 28702 19906 28754
rect 22318 28702 22370 28754
rect 30494 28702 30546 28754
rect 33294 28702 33346 28754
rect 35310 28702 35362 28754
rect 1710 28590 1762 28642
rect 2494 28590 2546 28642
rect 5742 28590 5794 28642
rect 6190 28590 6242 28642
rect 9550 28590 9602 28642
rect 9886 28590 9938 28642
rect 13582 28590 13634 28642
rect 18958 28590 19010 28642
rect 19518 28590 19570 28642
rect 20638 28590 20690 28642
rect 24334 28590 24386 28642
rect 24782 28590 24834 28642
rect 28030 28590 28082 28642
rect 35086 28590 35138 28642
rect 36318 28590 36370 28642
rect 40014 28590 40066 28642
rect 40462 28590 40514 28642
rect 2046 28478 2098 28530
rect 14478 28478 14530 28530
rect 16718 28478 16770 28530
rect 20190 28478 20242 28530
rect 23550 28478 23602 28530
rect 31502 28478 31554 28530
rect 34302 28478 34354 28530
rect 8654 28366 8706 28418
rect 12350 28366 12402 28418
rect 15038 28366 15090 28418
rect 27246 28366 27298 28418
rect 27806 28366 27858 28418
rect 28142 28366 28194 28418
rect 29262 28366 29314 28418
rect 37662 28366 37714 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 9102 28030 9154 28082
rect 12238 28030 12290 28082
rect 15598 28030 15650 28082
rect 16158 28030 16210 28082
rect 17502 28030 17554 28082
rect 29598 28030 29650 28082
rect 37662 28030 37714 28082
rect 39790 28030 39842 28082
rect 40238 28030 40290 28082
rect 2046 27918 2098 27970
rect 8318 27918 8370 27970
rect 9886 27918 9938 27970
rect 16494 27918 16546 27970
rect 16830 27918 16882 27970
rect 19742 27918 19794 27970
rect 25230 27918 25282 27970
rect 25566 27918 25618 27970
rect 36878 27918 36930 27970
rect 38894 27918 38946 27970
rect 1710 27806 1762 27858
rect 5630 27806 5682 27858
rect 6078 27806 6130 27858
rect 12686 27806 12738 27858
rect 13134 27806 13186 27858
rect 20190 27806 20242 27858
rect 26350 27806 26402 27858
rect 33966 27806 34018 27858
rect 34638 27806 34690 27858
rect 2494 27694 2546 27746
rect 11230 27694 11282 27746
rect 18398 27694 18450 27746
rect 21198 27694 21250 27746
rect 26126 27694 26178 27746
rect 37886 27694 37938 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 25006 27246 25058 27298
rect 29038 27246 29090 27298
rect 32846 27246 32898 27298
rect 33518 27246 33570 27298
rect 39902 27246 39954 27298
rect 6862 27134 6914 27186
rect 14142 27134 14194 27186
rect 18286 27134 18338 27186
rect 34974 27134 35026 27186
rect 37998 27134 38050 27186
rect 2830 27022 2882 27074
rect 8878 27022 8930 27074
rect 12238 27022 12290 27074
rect 12686 27022 12738 27074
rect 14926 27022 14978 27074
rect 16158 27022 16210 27074
rect 21870 27022 21922 27074
rect 28142 27022 28194 27074
rect 28702 27022 28754 27074
rect 32174 27022 32226 27074
rect 32734 27022 32786 27074
rect 40126 27022 40178 27074
rect 7870 26910 7922 26962
rect 8654 26910 8706 26962
rect 9998 26910 10050 26962
rect 29822 26910 29874 26962
rect 33182 26910 33234 26962
rect 33518 26910 33570 26962
rect 35982 26910 36034 26962
rect 39342 26910 39394 26962
rect 2158 26798 2210 26850
rect 9214 26798 9266 26850
rect 21982 26798 22034 26850
rect 25790 26798 25842 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 2942 26462 2994 26514
rect 3614 26462 3666 26514
rect 5406 26462 5458 26514
rect 6190 26462 6242 26514
rect 16382 26462 16434 26514
rect 17502 26462 17554 26514
rect 25902 26462 25954 26514
rect 38782 26462 38834 26514
rect 9774 26350 9826 26402
rect 10110 26350 10162 26402
rect 10558 26350 10610 26402
rect 16942 26350 16994 26402
rect 19406 26350 19458 26402
rect 20190 26350 20242 26402
rect 23774 26350 23826 26402
rect 3278 26238 3330 26290
rect 8542 26238 8594 26290
rect 9102 26238 9154 26290
rect 13022 26238 13074 26290
rect 13358 26238 13410 26290
rect 13918 26238 13970 26290
rect 20414 26238 20466 26290
rect 21086 26238 21138 26290
rect 21534 26238 21586 26290
rect 25790 26238 25842 26290
rect 28366 26238 28418 26290
rect 33182 26238 33234 26290
rect 38670 26238 38722 26290
rect 1822 26126 1874 26178
rect 2270 26126 2322 26178
rect 11790 26126 11842 26178
rect 18398 26126 18450 26178
rect 25342 26126 25394 26178
rect 28926 26126 28978 26178
rect 35646 26126 35698 26178
rect 39902 26126 39954 26178
rect 17278 26014 17330 26066
rect 17614 26014 17666 26066
rect 24558 26014 24610 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 9326 25678 9378 25730
rect 9662 25678 9714 25730
rect 22430 25678 22482 25730
rect 26462 25678 26514 25730
rect 40798 25678 40850 25730
rect 6974 25566 7026 25618
rect 7310 25566 7362 25618
rect 9102 25566 9154 25618
rect 9550 25566 9602 25618
rect 11454 25566 11506 25618
rect 17502 25566 17554 25618
rect 20526 25566 20578 25618
rect 26798 25566 26850 25618
rect 27246 25566 27298 25618
rect 2942 25454 2994 25506
rect 16270 25454 16322 25506
rect 22206 25454 22258 25506
rect 22990 25454 23042 25506
rect 23326 25454 23378 25506
rect 29262 25454 29314 25506
rect 29710 25454 29762 25506
rect 35982 25454 36034 25506
rect 36318 25454 36370 25506
rect 37102 25454 37154 25506
rect 37774 25454 37826 25506
rect 8094 25342 8146 25394
rect 12798 25342 12850 25394
rect 33630 25342 33682 25394
rect 2158 25230 2210 25282
rect 25902 25230 25954 25282
rect 32174 25230 32226 25282
rect 32734 25230 32786 25282
rect 32846 25230 32898 25282
rect 40014 25230 40066 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16606 24894 16658 24946
rect 22318 24894 22370 24946
rect 23438 24894 23490 24946
rect 25902 24894 25954 24946
rect 30718 24894 30770 24946
rect 33182 24894 33234 24946
rect 36094 24894 36146 24946
rect 36542 24894 36594 24946
rect 39342 24894 39394 24946
rect 7534 24782 7586 24834
rect 10446 24782 10498 24834
rect 15822 24782 15874 24834
rect 17390 24782 17442 24834
rect 18846 24782 18898 24834
rect 30158 24782 30210 24834
rect 32174 24782 32226 24834
rect 35310 24782 35362 24834
rect 37886 24782 37938 24834
rect 2942 24670 2994 24722
rect 15486 24670 15538 24722
rect 17614 24670 17666 24722
rect 18286 24670 18338 24722
rect 19630 24670 19682 24722
rect 20078 24670 20130 24722
rect 25678 24670 25730 24722
rect 30606 24670 30658 24722
rect 31726 24670 31778 24722
rect 39118 24670 39170 24722
rect 39902 24670 39954 24722
rect 1934 24558 1986 24610
rect 6190 24558 6242 24610
rect 16158 24558 16210 24610
rect 18062 24558 18114 24610
rect 19182 24558 19234 24610
rect 28814 24558 28866 24610
rect 33630 24558 33682 24610
rect 34078 24558 34130 24610
rect 36878 24558 36930 24610
rect 23102 24446 23154 24498
rect 35982 24446 36034 24498
rect 36654 24446 36706 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 34302 24110 34354 24162
rect 36990 24110 37042 24162
rect 15262 23998 15314 24050
rect 20414 23998 20466 24050
rect 22318 23998 22370 24050
rect 25118 23998 25170 24050
rect 35758 23998 35810 24050
rect 36206 23998 36258 24050
rect 10558 23886 10610 23938
rect 10894 23886 10946 23938
rect 16494 23886 16546 23938
rect 17166 23886 17218 23938
rect 30830 23886 30882 23938
rect 31278 23886 31330 23938
rect 35086 23886 35138 23938
rect 40126 23886 40178 23938
rect 40462 23886 40514 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 11566 23774 11618 23826
rect 11902 23774 11954 23826
rect 12350 23774 12402 23826
rect 14254 23774 14306 23826
rect 19406 23774 19458 23826
rect 20750 23774 20802 23826
rect 23326 23774 23378 23826
rect 26126 23774 26178 23826
rect 33518 23774 33570 23826
rect 2494 23662 2546 23714
rect 7422 23662 7474 23714
rect 8206 23662 8258 23714
rect 15710 23662 15762 23714
rect 20190 23662 20242 23714
rect 21422 23662 21474 23714
rect 30270 23662 30322 23714
rect 35198 23662 35250 23714
rect 37774 23662 37826 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 11230 23326 11282 23378
rect 17502 23326 17554 23378
rect 20750 23326 20802 23378
rect 21422 23326 21474 23378
rect 26462 23326 26514 23378
rect 26910 23326 26962 23378
rect 39230 23326 39282 23378
rect 39790 23326 39842 23378
rect 2382 23214 2434 23266
rect 6974 23214 7026 23266
rect 12574 23214 12626 23266
rect 15934 23214 15986 23266
rect 22318 23214 22370 23266
rect 35086 23214 35138 23266
rect 4734 23102 4786 23154
rect 5294 23102 5346 23154
rect 14926 23102 14978 23154
rect 15486 23102 15538 23154
rect 17838 23102 17890 23154
rect 18286 23102 18338 23154
rect 27246 23102 27298 23154
rect 36094 23102 36146 23154
rect 36766 23102 36818 23154
rect 40126 23102 40178 23154
rect 5630 22990 5682 23042
rect 7982 22990 8034 23042
rect 16270 22990 16322 23042
rect 23438 22990 23490 23042
rect 30158 22990 30210 23042
rect 33182 22990 33234 23042
rect 33742 22990 33794 23042
rect 34078 22990 34130 23042
rect 1598 22878 1650 22930
rect 11790 22878 11842 22930
rect 33182 22878 33234 22930
rect 33630 22878 33682 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 15710 22542 15762 22594
rect 39902 22542 39954 22594
rect 2494 22430 2546 22482
rect 8094 22430 8146 22482
rect 13582 22430 13634 22482
rect 14590 22430 14642 22482
rect 14926 22430 14978 22482
rect 37102 22430 37154 22482
rect 37550 22430 37602 22482
rect 37998 22430 38050 22482
rect 41022 22430 41074 22482
rect 1710 22318 1762 22370
rect 9550 22318 9602 22370
rect 9886 22318 9938 22370
rect 18734 22318 18786 22370
rect 19182 22318 19234 22370
rect 20414 22318 20466 22370
rect 21646 22318 21698 22370
rect 22878 22318 22930 22370
rect 23326 22318 23378 22370
rect 27022 22318 27074 22370
rect 27694 22318 27746 22370
rect 32174 22318 32226 22370
rect 32510 22318 32562 22370
rect 32846 22318 32898 22370
rect 33518 22318 33570 22370
rect 40014 22318 40066 22370
rect 2046 22206 2098 22258
rect 7086 22206 7138 22258
rect 13918 22206 13970 22258
rect 14254 22206 14306 22258
rect 26350 22206 26402 22258
rect 35758 22206 35810 22258
rect 39006 22206 39058 22258
rect 12462 22094 12514 22146
rect 13022 22094 13074 22146
rect 16494 22094 16546 22146
rect 20638 22094 20690 22146
rect 21758 22094 21810 22146
rect 25566 22094 25618 22146
rect 27246 22094 27298 22146
rect 28254 22094 28306 22146
rect 29038 22094 29090 22146
rect 29598 22094 29650 22146
rect 36542 22094 36594 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 5294 21758 5346 21810
rect 9438 21758 9490 21810
rect 10222 21758 10274 21810
rect 16158 21758 16210 21810
rect 17502 21758 17554 21810
rect 20974 21758 21026 21810
rect 21758 21758 21810 21810
rect 28030 21758 28082 21810
rect 32062 21758 32114 21810
rect 33182 21758 33234 21810
rect 37438 21758 37490 21810
rect 38446 21758 38498 21810
rect 39566 21758 39618 21810
rect 4510 21646 4562 21698
rect 6974 21646 7026 21698
rect 20078 21646 20130 21698
rect 1822 21534 1874 21586
rect 2158 21534 2210 21586
rect 5630 21534 5682 21586
rect 12462 21534 12514 21586
rect 13134 21534 13186 21586
rect 13470 21534 13522 21586
rect 13806 21534 13858 21586
rect 23998 21534 24050 21586
rect 24446 21534 24498 21586
rect 25118 21534 25170 21586
rect 25790 21534 25842 21586
rect 29150 21534 29202 21586
rect 29598 21534 29650 21586
rect 33406 21534 33458 21586
rect 34638 21534 34690 21586
rect 35086 21534 35138 21586
rect 38670 21534 38722 21586
rect 39790 21534 39842 21586
rect 7982 21422 8034 21474
rect 18734 21422 18786 21474
rect 16942 21310 16994 21362
rect 28814 21310 28866 21362
rect 32622 21310 32674 21362
rect 38110 21310 38162 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17054 20974 17106 21026
rect 34414 20974 34466 21026
rect 34638 20974 34690 21026
rect 35198 20974 35250 21026
rect 3838 20862 3890 20914
rect 10782 20862 10834 20914
rect 11006 20862 11058 20914
rect 11454 20862 11506 20914
rect 12910 20862 12962 20914
rect 17390 20862 17442 20914
rect 19070 20862 19122 20914
rect 19742 20862 19794 20914
rect 24894 20862 24946 20914
rect 34862 20862 34914 20914
rect 35198 20862 35250 20914
rect 37214 20862 37266 20914
rect 37774 20862 37826 20914
rect 37998 20862 38050 20914
rect 40014 20862 40066 20914
rect 1710 20750 1762 20802
rect 6190 20750 6242 20802
rect 6750 20750 6802 20802
rect 7310 20750 7362 20802
rect 13582 20750 13634 20802
rect 13918 20750 13970 20802
rect 20862 20750 20914 20802
rect 21422 20750 21474 20802
rect 27582 20750 27634 20802
rect 30942 20750 30994 20802
rect 31390 20750 31442 20802
rect 2046 20638 2098 20690
rect 2718 20638 2770 20690
rect 16270 20638 16322 20690
rect 17950 20638 18002 20690
rect 39006 20638 39058 20690
rect 5966 20526 6018 20578
rect 9662 20526 9714 20578
rect 10446 20526 10498 20578
rect 27694 20526 27746 20578
rect 33742 20526 33794 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 1822 20190 1874 20242
rect 3614 20190 3666 20242
rect 5854 20190 5906 20242
rect 16606 20190 16658 20242
rect 33742 20190 33794 20242
rect 10670 20078 10722 20130
rect 25566 20078 25618 20130
rect 30046 20078 30098 20130
rect 35870 20078 35922 20130
rect 3390 19966 3442 20018
rect 4062 19966 4114 20018
rect 8094 19966 8146 20018
rect 8766 19966 8818 20018
rect 14814 19966 14866 20018
rect 16606 19966 16658 20018
rect 17390 19966 17442 20018
rect 25678 19966 25730 20018
rect 27246 19966 27298 20018
rect 27806 19966 27858 20018
rect 32510 19966 32562 20018
rect 33518 19966 33570 20018
rect 38110 19966 38162 20018
rect 38782 19966 38834 20018
rect 39118 19966 39170 20018
rect 9774 19854 9826 19906
rect 11902 19854 11954 19906
rect 15262 19854 15314 19906
rect 20078 19854 20130 19906
rect 21758 19854 21810 19906
rect 26686 19854 26738 19906
rect 4174 19742 4226 19794
rect 5070 19742 5122 19794
rect 30830 19742 30882 19794
rect 35086 19742 35138 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 4062 19294 4114 19346
rect 7310 19294 7362 19346
rect 26126 19294 26178 19346
rect 33966 19294 34018 19346
rect 37998 19294 38050 19346
rect 11790 19182 11842 19234
rect 12462 19182 12514 19234
rect 13582 19182 13634 19234
rect 13918 19182 13970 19234
rect 20302 19182 20354 19234
rect 20862 19182 20914 19234
rect 21198 19182 21250 19234
rect 21758 19182 21810 19234
rect 32174 19182 32226 19234
rect 32622 19182 32674 19234
rect 33070 19182 33122 19234
rect 3054 19070 3106 19122
rect 6190 19070 6242 19122
rect 24110 19070 24162 19122
rect 24894 19070 24946 19122
rect 27134 19070 27186 19122
rect 34974 19070 35026 19122
rect 39006 19070 39058 19122
rect 8766 18958 8818 19010
rect 9326 18958 9378 19010
rect 12798 18958 12850 19010
rect 16382 18958 16434 19010
rect 17054 18958 17106 19010
rect 17166 18958 17218 19010
rect 17838 18958 17890 19010
rect 25790 18958 25842 19010
rect 29038 18958 29090 19010
rect 29822 18958 29874 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 3054 18622 3106 18674
rect 3838 18622 3890 18674
rect 8878 18622 8930 18674
rect 13246 18622 13298 18674
rect 10334 18510 10386 18562
rect 19518 18510 19570 18562
rect 24558 18510 24610 18562
rect 27246 18510 27298 18562
rect 2382 18398 2434 18450
rect 6078 18398 6130 18450
rect 6526 18398 6578 18450
rect 7534 18398 7586 18450
rect 8990 18398 9042 18450
rect 15598 18398 15650 18450
rect 16270 18398 16322 18450
rect 17614 18398 17666 18450
rect 18510 18398 18562 18450
rect 19070 18398 19122 18450
rect 26350 18398 26402 18450
rect 30718 18398 30770 18450
rect 33518 18398 33570 18450
rect 38670 18398 38722 18450
rect 2270 18286 2322 18338
rect 7758 18286 7810 18338
rect 11342 18286 11394 18338
rect 16606 18286 16658 18338
rect 17950 18286 18002 18338
rect 20750 18286 20802 18338
rect 23214 18286 23266 18338
rect 35310 18286 35362 18338
rect 38782 18286 38834 18338
rect 39902 18286 39954 18338
rect 12574 18174 12626 18226
rect 26238 18174 26290 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 13022 17838 13074 17890
rect 14030 17838 14082 17890
rect 3502 17726 3554 17778
rect 6302 17726 6354 17778
rect 8094 17726 8146 17778
rect 16830 17726 16882 17778
rect 20750 17726 20802 17778
rect 22878 17726 22930 17778
rect 32510 17726 32562 17778
rect 33518 17726 33570 17778
rect 34638 17726 34690 17778
rect 37998 17726 38050 17778
rect 2382 17614 2434 17666
rect 3390 17614 3442 17666
rect 4734 17614 4786 17666
rect 9550 17614 9602 17666
rect 9886 17614 9938 17666
rect 13918 17614 13970 17666
rect 20078 17614 20130 17666
rect 24110 17614 24162 17666
rect 28590 17614 28642 17666
rect 29150 17614 29202 17666
rect 35422 17614 35474 17666
rect 39790 17614 39842 17666
rect 41022 17614 41074 17666
rect 7086 17502 7138 17554
rect 39006 17502 39058 17554
rect 2158 17390 2210 17442
rect 4958 17390 5010 17442
rect 12462 17390 12514 17442
rect 13582 17390 13634 17442
rect 26910 17390 26962 17442
rect 27582 17390 27634 17442
rect 35646 17390 35698 17442
rect 39902 17390 39954 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 2158 17054 2210 17106
rect 5630 17054 5682 17106
rect 28030 17054 28082 17106
rect 36094 17054 36146 17106
rect 8878 16942 8930 16994
rect 10558 16942 10610 16994
rect 22094 16942 22146 16994
rect 28814 16942 28866 16994
rect 31054 16942 31106 16994
rect 39566 16942 39618 16994
rect 4734 16830 4786 16882
rect 5294 16830 5346 16882
rect 15486 16830 15538 16882
rect 18958 16830 19010 16882
rect 19406 16830 19458 16882
rect 19742 16830 19794 16882
rect 25342 16830 25394 16882
rect 25790 16830 25842 16882
rect 33182 16830 33234 16882
rect 33854 16830 33906 16882
rect 37214 16830 37266 16882
rect 37662 16830 37714 16882
rect 7534 16718 7586 16770
rect 15934 16718 15986 16770
rect 30046 16718 30098 16770
rect 38558 16718 38610 16770
rect 1598 16606 1650 16658
rect 22878 16606 22930 16658
rect 36878 16606 36930 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 13582 16270 13634 16322
rect 21982 16270 22034 16322
rect 30382 16270 30434 16322
rect 4062 16158 4114 16210
rect 11790 16158 11842 16210
rect 18398 16158 18450 16210
rect 29710 16158 29762 16210
rect 36430 16158 36482 16210
rect 8542 16046 8594 16098
rect 9214 16046 9266 16098
rect 13806 16046 13858 16098
rect 16158 16046 16210 16098
rect 22094 16046 22146 16098
rect 23550 16046 23602 16098
rect 23998 16046 24050 16098
rect 29934 16046 29986 16098
rect 30270 16046 30322 16098
rect 31502 16046 31554 16098
rect 31950 16046 32002 16098
rect 35534 16046 35586 16098
rect 40126 16046 40178 16098
rect 40574 16046 40626 16098
rect 3054 15934 3106 15986
rect 5518 15934 5570 15986
rect 10558 15934 10610 15986
rect 26238 15934 26290 15986
rect 37886 15934 37938 15986
rect 6078 15822 6130 15874
rect 9550 15822 9602 15874
rect 20526 15822 20578 15874
rect 27022 15822 27074 15874
rect 28590 15822 28642 15874
rect 34414 15822 34466 15874
rect 34974 15822 35026 15874
rect 35310 15822 35362 15874
rect 37102 15822 37154 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 7422 15486 7474 15538
rect 13246 15486 13298 15538
rect 35982 15486 36034 15538
rect 36542 15486 36594 15538
rect 1934 15374 1986 15426
rect 19406 15374 19458 15426
rect 21310 15374 21362 15426
rect 28702 15374 28754 15426
rect 32062 15374 32114 15426
rect 35086 15374 35138 15426
rect 39678 15374 39730 15426
rect 4734 15262 4786 15314
rect 5070 15262 5122 15314
rect 15150 15262 15202 15314
rect 15598 15262 15650 15314
rect 16718 15262 16770 15314
rect 23662 15262 23714 15314
rect 24222 15262 24274 15314
rect 29934 15262 29986 15314
rect 36766 15262 36818 15314
rect 37438 15262 37490 15314
rect 3278 15150 3330 15202
rect 8542 15150 8594 15202
rect 18398 15150 18450 15202
rect 20526 15150 20578 15202
rect 27582 15150 27634 15202
rect 30718 15150 30770 15202
rect 34078 15150 34130 15202
rect 8206 15038 8258 15090
rect 16718 15038 16770 15090
rect 40462 15038 40514 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 22318 14702 22370 14754
rect 3950 14590 4002 14642
rect 11342 14590 11394 14642
rect 20750 14590 20802 14642
rect 21422 14590 21474 14642
rect 24446 14590 24498 14642
rect 29934 14590 29986 14642
rect 34974 14590 35026 14642
rect 6414 14478 6466 14530
rect 7086 14478 7138 14530
rect 15822 14478 15874 14530
rect 16270 14478 16322 14530
rect 20302 14478 20354 14530
rect 22206 14478 22258 14530
rect 32398 14478 32450 14530
rect 32734 14478 32786 14530
rect 40014 14478 40066 14530
rect 40350 14478 40402 14530
rect 2718 14366 2770 14418
rect 10110 14366 10162 14418
rect 12350 14366 12402 14418
rect 18510 14366 18562 14418
rect 25454 14366 25506 14418
rect 30942 14366 30994 14418
rect 36318 14366 36370 14418
rect 9550 14254 9602 14306
rect 10446 14254 10498 14306
rect 19294 14254 19346 14306
rect 20190 14254 20242 14306
rect 27246 14254 27298 14306
rect 32846 14254 32898 14306
rect 36878 14254 36930 14306
rect 37662 14254 37714 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 1598 13918 1650 13970
rect 2270 13918 2322 13970
rect 5630 13918 5682 13970
rect 16382 13918 16434 13970
rect 20190 13918 20242 13970
rect 29822 13918 29874 13970
rect 36990 13918 37042 13970
rect 39790 13918 39842 13970
rect 8542 13806 8594 13858
rect 10670 13806 10722 13858
rect 23998 13806 24050 13858
rect 29038 13806 29090 13858
rect 32062 13806 32114 13858
rect 35870 13806 35922 13858
rect 37774 13806 37826 13858
rect 4622 13694 4674 13746
rect 5182 13694 5234 13746
rect 13358 13694 13410 13746
rect 13918 13694 13970 13746
rect 17502 13694 17554 13746
rect 17950 13694 18002 13746
rect 21310 13694 21362 13746
rect 21758 13694 21810 13746
rect 26126 13694 26178 13746
rect 26798 13694 26850 13746
rect 33182 13694 33234 13746
rect 33630 13694 33682 13746
rect 7534 13582 7586 13634
rect 12014 13582 12066 13634
rect 31054 13582 31106 13634
rect 38894 13582 38946 13634
rect 16942 13470 16994 13522
rect 20974 13470 21026 13522
rect 24782 13470 24834 13522
rect 36654 13470 36706 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 4174 13134 4226 13186
rect 23214 13134 23266 13186
rect 27358 13134 27410 13186
rect 16494 13022 16546 13074
rect 19518 13022 19570 13074
rect 33070 13022 33122 13074
rect 33518 13022 33570 13074
rect 33966 13022 34018 13074
rect 37102 13022 37154 13074
rect 38334 13022 38386 13074
rect 40350 13022 40402 13074
rect 3950 12910 4002 12962
rect 6974 12910 7026 12962
rect 10334 12910 10386 12962
rect 10670 12910 10722 12962
rect 12462 12910 12514 12962
rect 13582 12910 13634 12962
rect 21646 12910 21698 12962
rect 22654 12910 22706 12962
rect 23774 12910 23826 12962
rect 24334 12910 24386 12962
rect 27806 12910 27858 12962
rect 29262 12910 29314 12962
rect 29710 12910 29762 12962
rect 40126 12910 40178 12962
rect 17502 12798 17554 12850
rect 20638 12798 20690 12850
rect 21534 12798 21586 12850
rect 32734 12798 32786 12850
rect 34974 12798 35026 12850
rect 39342 12798 39394 12850
rect 6862 12686 6914 12738
rect 7198 12686 7250 12738
rect 7758 12686 7810 12738
rect 11230 12686 11282 12738
rect 12238 12686 12290 12738
rect 14142 12686 14194 12738
rect 16158 12686 16210 12738
rect 26798 12686 26850 12738
rect 27694 12686 27746 12738
rect 32174 12686 32226 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 9662 12350 9714 12402
rect 14926 12350 14978 12402
rect 17502 12350 17554 12402
rect 17950 12350 18002 12402
rect 29486 12350 29538 12402
rect 33294 12350 33346 12402
rect 37102 12350 37154 12402
rect 38110 12350 38162 12402
rect 39342 12350 39394 12402
rect 8318 12238 8370 12290
rect 19742 12238 19794 12290
rect 21198 12238 21250 12290
rect 25902 12238 25954 12290
rect 5630 12126 5682 12178
rect 6078 12126 6130 12178
rect 9886 12126 9938 12178
rect 11790 12126 11842 12178
rect 12238 12126 12290 12178
rect 12574 12126 12626 12178
rect 16718 12126 16770 12178
rect 23438 12126 23490 12178
rect 23886 12126 23938 12178
rect 28254 12126 28306 12178
rect 28590 12126 28642 12178
rect 32062 12126 32114 12178
rect 32622 12126 32674 12178
rect 33518 12126 33570 12178
rect 34078 12126 34130 12178
rect 34750 12126 34802 12178
rect 39230 12126 39282 12178
rect 18734 12014 18786 12066
rect 9102 11902 9154 11954
rect 11678 11902 11730 11954
rect 15710 11902 15762 11954
rect 16718 11902 16770 11954
rect 20414 11902 20466 11954
rect 25118 11902 25170 11954
rect 28926 11902 28978 11954
rect 37774 11902 37826 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 9326 11566 9378 11618
rect 27582 11566 27634 11618
rect 37102 11566 37154 11618
rect 7646 11454 7698 11506
rect 14926 11454 14978 11506
rect 22318 11454 22370 11506
rect 25678 11454 25730 11506
rect 33966 11454 34018 11506
rect 36542 11454 36594 11506
rect 38446 11454 38498 11506
rect 40686 11454 40738 11506
rect 12350 11342 12402 11394
rect 13022 11342 13074 11394
rect 19630 11342 19682 11394
rect 20078 11342 20130 11394
rect 27582 11342 27634 11394
rect 30046 11342 30098 11394
rect 30718 11342 30770 11394
rect 36990 11342 37042 11394
rect 8654 11230 8706 11282
rect 10110 11230 10162 11282
rect 15934 11230 15986 11282
rect 23550 11230 23602 11282
rect 27022 11230 27074 11282
rect 34974 11230 35026 11282
rect 41694 11230 41746 11282
rect 13582 11118 13634 11170
rect 14590 11118 14642 11170
rect 16606 11118 16658 11170
rect 17166 11118 17218 11170
rect 33182 11118 33234 11170
rect 33742 11118 33794 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 8318 10782 8370 10834
rect 16494 10782 16546 10834
rect 17502 10782 17554 10834
rect 21534 10782 21586 10834
rect 22654 10782 22706 10834
rect 32622 10782 32674 10834
rect 33182 10782 33234 10834
rect 34414 10782 34466 10834
rect 11566 10670 11618 10722
rect 15374 10670 15426 10722
rect 26238 10670 26290 10722
rect 30046 10670 30098 10722
rect 37886 10670 37938 10722
rect 8542 10558 8594 10610
rect 12686 10558 12738 10610
rect 13134 10558 13186 10610
rect 17726 10558 17778 10610
rect 18622 10558 18674 10610
rect 19294 10558 19346 10610
rect 22542 10558 22594 10610
rect 33070 10558 33122 10610
rect 9662 10446 9714 10498
rect 10558 10446 10610 10498
rect 27358 10446 27410 10498
rect 28030 10446 28082 10498
rect 31166 10446 31218 10498
rect 32062 10446 32114 10498
rect 36878 10446 36930 10498
rect 16158 10334 16210 10386
rect 22318 10334 22370 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 14366 9998 14418 10050
rect 28478 9998 28530 10050
rect 18958 9886 19010 9938
rect 19406 9886 19458 9938
rect 24334 9886 24386 9938
rect 30046 9886 30098 9938
rect 40238 9886 40290 9938
rect 2942 9774 2994 9826
rect 9550 9774 9602 9826
rect 9998 9774 10050 9826
rect 13806 9774 13858 9826
rect 15038 9774 15090 9826
rect 15486 9774 15538 9826
rect 27582 9774 27634 9826
rect 28590 9774 28642 9826
rect 29486 9774 29538 9826
rect 30494 9774 30546 9826
rect 2046 9662 2098 9714
rect 12238 9662 12290 9714
rect 23214 9662 23266 9714
rect 39118 9662 39170 9714
rect 13022 9550 13074 9602
rect 17726 9550 17778 9602
rect 18510 9550 18562 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 13022 9102 13074 9154
rect 16718 9102 16770 9154
rect 17726 9102 17778 9154
rect 21982 9102 22034 9154
rect 2942 8990 2994 9042
rect 10446 8990 10498 9042
rect 17838 8990 17890 9042
rect 1934 8878 1986 8930
rect 12014 8878 12066 8930
rect 13918 8878 13970 8930
rect 15374 8878 15426 8930
rect 20974 8878 21026 8930
rect 10334 8766 10386 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 11678 8318 11730 8370
rect 12126 8318 12178 8370
rect 16270 8318 16322 8370
rect 19518 8318 19570 8370
rect 2718 8206 2770 8258
rect 8206 8206 8258 8258
rect 8654 8206 8706 8258
rect 2046 8094 2098 8146
rect 10894 8094 10946 8146
rect 17278 8094 17330 8146
rect 18398 8094 18450 8146
rect 3278 7982 3330 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 14254 7534 14306 7586
rect 2942 7422 2994 7474
rect 1934 7310 1986 7362
rect 13246 7310 13298 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 2830 6638 2882 6690
rect 2046 6526 2098 6578
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 3278 6078 3330 6130
rect 2718 5854 2770 5906
rect 3502 5854 3554 5906
rect 1934 5742 1986 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 3838 5070 3890 5122
rect 4510 5070 4562 5122
rect 6974 5070 7026 5122
rect 10446 5070 10498 5122
rect 2270 4958 2322 5010
rect 2606 4958 2658 5010
rect 2942 4958 2994 5010
rect 3278 4958 3330 5010
rect 3614 4958 3666 5010
rect 4286 4958 4338 5010
rect 1710 4846 1762 4898
rect 7310 4846 7362 4898
rect 10670 4846 10722 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 2046 4510 2098 4562
rect 2942 4510 2994 4562
rect 3614 4510 3666 4562
rect 1710 4398 1762 4450
rect 2382 4398 2434 4450
rect 3278 4398 3330 4450
rect 4846 4398 4898 4450
rect 3838 4286 3890 4338
rect 4398 4174 4450 4226
rect 5294 4174 5346 4226
rect 5742 4174 5794 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 7982 3614 8034 3666
rect 11454 3614 11506 3666
rect 1710 3502 1762 3554
rect 3950 3502 4002 3554
rect 7534 3502 7586 3554
rect 11006 3502 11058 3554
rect 2046 3390 2098 3442
rect 2382 3390 2434 3442
rect 2718 3390 2770 3442
rect 3054 3390 3106 3442
rect 3390 3390 3442 3442
rect 3726 3390 3778 3442
rect 4510 3390 4562 3442
rect 4958 3390 5010 3442
rect 6078 3390 6130 3442
rect 6302 3390 6354 3442
rect 6638 3390 6690 3442
rect 10110 3390 10162 3442
rect 10334 3390 10386 3442
rect 10670 3390 10722 3442
rect 6974 3278 7026 3330
rect 9326 3278 9378 3330
rect 13134 3278 13186 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 12126 1710 12178 1762
rect 13134 1710 13186 1762
<< metal2 >>
rect 0 43200 112 44000
rect 672 43200 784 44000
rect 1344 43200 1456 44000
rect 2016 43200 2128 44000
rect 2688 43200 2800 44000
rect 3360 43200 3472 44000
rect 4032 43200 4144 44000
rect 4284 43204 4340 43214
rect 28 40180 84 43200
rect 28 40114 84 40124
rect 700 36820 756 43200
rect 1372 39060 1428 43200
rect 1932 43092 1988 43102
rect 1932 41300 1988 43036
rect 2044 41412 2100 43200
rect 2044 41356 2548 41412
rect 1932 41244 2324 41300
rect 1820 40628 1876 40638
rect 1820 40534 1876 40572
rect 1372 38994 1428 39004
rect 2044 40292 2100 40302
rect 1932 38836 1988 38846
rect 1820 38724 1876 38734
rect 1708 38722 1876 38724
rect 1708 38670 1822 38722
rect 1874 38670 1876 38722
rect 1708 38668 1876 38670
rect 1596 37716 1652 37726
rect 812 36820 868 36830
rect 700 36764 812 36820
rect 812 36754 868 36764
rect 1596 36484 1652 37660
rect 1596 36418 1652 36428
rect 1708 36482 1764 38668
rect 1820 38658 1876 38668
rect 1932 38052 1988 38780
rect 2044 38276 2100 40236
rect 2156 39060 2212 39070
rect 2156 38966 2212 39004
rect 2156 38276 2212 38286
rect 2044 38274 2212 38276
rect 2044 38222 2158 38274
rect 2210 38222 2212 38274
rect 2044 38220 2212 38222
rect 2156 38210 2212 38220
rect 1932 37996 2100 38052
rect 1932 37826 1988 37838
rect 1932 37774 1934 37826
rect 1986 37774 1988 37826
rect 1708 36430 1710 36482
rect 1762 36430 1764 36482
rect 1708 36036 1764 36430
rect 1708 35970 1764 35980
rect 1820 37154 1876 37166
rect 1820 37102 1822 37154
rect 1874 37102 1876 37154
rect 1708 35700 1764 35710
rect 1820 35700 1876 37102
rect 1932 36372 1988 37774
rect 1932 36306 1988 36316
rect 2044 36370 2100 37996
rect 2156 37492 2212 37502
rect 2268 37492 2324 41244
rect 2492 39842 2548 41356
rect 2716 40290 2772 43200
rect 3388 42644 3444 43200
rect 3388 42588 4004 42644
rect 3388 42420 3444 42430
rect 3444 42364 3556 42420
rect 3388 42354 3444 42364
rect 3388 41076 3444 41086
rect 3276 40404 3332 40414
rect 3276 40310 3332 40348
rect 2716 40238 2718 40290
rect 2770 40238 2772 40290
rect 2716 40226 2772 40238
rect 2492 39790 2494 39842
rect 2546 39790 2548 39842
rect 2492 39778 2548 39790
rect 3276 39396 3332 39406
rect 3276 39302 3332 39340
rect 2940 38948 2996 38958
rect 2940 38854 2996 38892
rect 3388 38164 3444 41020
rect 3500 38388 3556 42364
rect 3724 41748 3780 41758
rect 3724 39058 3780 41692
rect 3948 40292 4004 42588
rect 4060 40514 4116 43200
rect 4704 43200 4816 44000
rect 5376 43200 5488 44000
rect 6048 43200 6160 44000
rect 6720 43200 6832 44000
rect 7392 43200 7504 44000
rect 8064 43200 8176 44000
rect 8736 43200 8848 44000
rect 9408 43200 9520 44000
rect 10080 43200 10192 44000
rect 10752 43200 10864 44000
rect 11424 43200 11536 44000
rect 12096 43200 12208 44000
rect 12768 43200 12880 44000
rect 13440 43200 13552 44000
rect 14112 43200 14224 44000
rect 14784 43200 14896 44000
rect 15456 43200 15568 44000
rect 16128 43200 16240 44000
rect 16800 43200 16912 44000
rect 17472 43200 17584 44000
rect 18144 43200 18256 44000
rect 18816 43200 18928 44000
rect 19488 43200 19600 44000
rect 20160 43200 20272 44000
rect 20832 43200 20944 44000
rect 21504 43200 21616 44000
rect 22176 43200 22288 44000
rect 22848 43200 22960 44000
rect 23520 43200 23632 44000
rect 24192 43200 24304 44000
rect 24864 43200 24976 44000
rect 25536 43200 25648 44000
rect 26208 43200 26320 44000
rect 26880 43200 26992 44000
rect 27244 43260 27636 43316
rect 4284 41188 4340 43148
rect 4284 41122 4340 41132
rect 4732 40628 4788 43200
rect 5404 41074 5460 43200
rect 5404 41022 5406 41074
rect 5458 41022 5460 41074
rect 5404 41010 5460 41022
rect 5964 41074 6020 41086
rect 5964 41022 5966 41074
rect 6018 41022 6020 41074
rect 4732 40562 4788 40572
rect 4060 40462 4062 40514
rect 4114 40462 4116 40514
rect 4060 40450 4116 40462
rect 4956 40516 5012 40526
rect 4956 40402 5012 40460
rect 5740 40516 5796 40526
rect 4956 40350 4958 40402
rect 5010 40350 5012 40402
rect 4956 40338 5012 40350
rect 5628 40404 5684 40414
rect 3948 40236 4116 40292
rect 4060 39842 4116 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4060 39790 4062 39842
rect 4114 39790 4116 39842
rect 4060 39778 4116 39790
rect 3724 39006 3726 39058
rect 3778 39006 3780 39058
rect 3724 38994 3780 39006
rect 3948 39732 4004 39742
rect 3500 38322 3556 38332
rect 3388 38108 3892 38164
rect 3612 37940 3668 37950
rect 3500 37938 3668 37940
rect 3500 37886 3614 37938
rect 3666 37886 3668 37938
rect 3500 37884 3668 37886
rect 2716 37828 2772 37838
rect 2156 37490 2324 37492
rect 2156 37438 2158 37490
rect 2210 37438 2324 37490
rect 2156 37436 2324 37438
rect 2604 37772 2716 37828
rect 2156 37426 2212 37436
rect 2380 36820 2436 36830
rect 2436 36764 2548 36820
rect 2380 36754 2436 36764
rect 2044 36318 2046 36370
rect 2098 36318 2100 36370
rect 2044 36306 2100 36318
rect 2380 36372 2436 36382
rect 2380 36278 2436 36316
rect 2380 36036 2436 36046
rect 2044 35980 2380 36036
rect 2044 35922 2100 35980
rect 2380 35970 2436 35980
rect 2044 35870 2046 35922
rect 2098 35870 2100 35922
rect 2044 35858 2100 35870
rect 2380 35812 2436 35822
rect 2492 35812 2548 36764
rect 2380 35810 2548 35812
rect 2380 35758 2382 35810
rect 2434 35758 2548 35810
rect 2380 35756 2548 35758
rect 2380 35746 2436 35756
rect 1708 35698 1876 35700
rect 1708 35646 1710 35698
rect 1762 35646 1876 35698
rect 1708 35644 1876 35646
rect 1708 35028 1764 35644
rect 1708 34962 1764 34972
rect 2156 35252 2212 35262
rect 2044 34802 2100 34814
rect 2044 34750 2046 34802
rect 2098 34750 2100 34802
rect 2044 34356 2100 34750
rect 2044 34290 2100 34300
rect 2156 34354 2212 35196
rect 2156 34302 2158 34354
rect 2210 34302 2212 34354
rect 2156 34290 2212 34302
rect 1708 34242 1764 34254
rect 1708 34190 1710 34242
rect 1762 34190 1764 34242
rect 1708 33684 1764 34190
rect 1708 33618 1764 33628
rect 1708 33234 1764 33246
rect 1708 33182 1710 33234
rect 1762 33182 1764 33234
rect 1708 33012 1764 33182
rect 2044 33236 2100 33246
rect 2044 33142 2100 33180
rect 1708 32946 1764 32956
rect 2492 33122 2548 33134
rect 2492 33070 2494 33122
rect 2546 33070 2548 33122
rect 2492 33012 2548 33070
rect 2492 32946 2548 32956
rect 1708 32674 1764 32686
rect 1708 32622 1710 32674
rect 1762 32622 1764 32674
rect 1708 32340 1764 32622
rect 1708 32274 1764 32284
rect 2604 31948 2660 37772
rect 2716 37762 2772 37772
rect 2940 37828 2996 37838
rect 3276 37828 3332 37838
rect 2940 37826 3108 37828
rect 2940 37774 2942 37826
rect 2994 37774 3108 37826
rect 2940 37772 3108 37774
rect 2940 37762 2996 37772
rect 2940 37492 2996 37502
rect 2940 37398 2996 37436
rect 2716 37156 2772 37166
rect 2716 36370 2772 37100
rect 3052 36820 3108 37772
rect 3276 37734 3332 37772
rect 3276 37380 3332 37390
rect 2940 36764 3108 36820
rect 3164 37378 3332 37380
rect 3164 37326 3278 37378
rect 3330 37326 3332 37378
rect 3164 37324 3332 37326
rect 2716 36318 2718 36370
rect 2770 36318 2772 36370
rect 2716 36306 2772 36318
rect 2828 36708 2884 36718
rect 2716 34916 2772 34926
rect 2828 34916 2884 36652
rect 2940 35922 2996 36764
rect 2940 35870 2942 35922
rect 2994 35870 2996 35922
rect 2940 35858 2996 35870
rect 3052 36258 3108 36270
rect 3052 36206 3054 36258
rect 3106 36206 3108 36258
rect 3052 34916 3108 36206
rect 2716 34914 2884 34916
rect 2716 34862 2718 34914
rect 2770 34862 2884 34914
rect 2716 34860 2884 34862
rect 2940 34860 3108 34916
rect 3164 34916 3220 37324
rect 3276 37314 3332 37324
rect 3276 36482 3332 36494
rect 3276 36430 3278 36482
rect 3330 36430 3332 36482
rect 3276 36036 3332 36430
rect 3276 35970 3332 35980
rect 3388 36372 3444 36382
rect 3276 35812 3332 35822
rect 3276 35718 3332 35756
rect 2716 34850 2772 34860
rect 2828 34692 2884 34702
rect 2604 31892 2772 31948
rect 2716 31778 2772 31892
rect 2716 31726 2718 31778
rect 2770 31726 2772 31778
rect 2716 31714 2772 31726
rect 1932 31668 1988 31678
rect 1932 30882 1988 31612
rect 2044 31666 2100 31678
rect 2044 31614 2046 31666
rect 2098 31614 2100 31666
rect 2044 31108 2100 31614
rect 2044 31042 2100 31052
rect 1932 30830 1934 30882
rect 1986 30830 1988 30882
rect 1932 30818 1988 30830
rect 2044 30884 2100 30894
rect 1708 30098 1764 30110
rect 1708 30046 1710 30098
rect 1762 30046 1764 30098
rect 1708 29652 1764 30046
rect 2044 30098 2100 30828
rect 2716 30772 2772 30782
rect 2380 30324 2436 30334
rect 2380 30210 2436 30268
rect 2380 30158 2382 30210
rect 2434 30158 2436 30210
rect 2380 30146 2436 30158
rect 2044 30046 2046 30098
rect 2098 30046 2100 30098
rect 2044 30034 2100 30046
rect 2716 30098 2772 30716
rect 2716 30046 2718 30098
rect 2770 30046 2772 30098
rect 2716 30034 2772 30046
rect 1708 29586 1764 29596
rect 2044 29876 2100 29886
rect 2044 29650 2100 29820
rect 2044 29598 2046 29650
rect 2098 29598 2100 29650
rect 2044 29586 2100 29598
rect 1708 29426 1764 29438
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 28980 1764 29374
rect 1708 28914 1764 28924
rect 2044 29316 2100 29326
rect 1708 28642 1764 28654
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 28308 1764 28590
rect 2044 28530 2100 29260
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 28980 2548 29262
rect 2492 28914 2548 28924
rect 2044 28478 2046 28530
rect 2098 28478 2100 28530
rect 2044 28466 2100 28478
rect 2492 28642 2548 28654
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 1708 28242 1764 28252
rect 2492 28308 2548 28590
rect 2492 28242 2548 28252
rect 2044 27972 2100 27982
rect 2044 27878 2100 27916
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27636 1764 27806
rect 1708 27570 1764 27580
rect 2492 27746 2548 27758
rect 2492 27694 2494 27746
rect 2546 27694 2548 27746
rect 2492 27636 2548 27694
rect 2492 27570 2548 27580
rect 2828 27074 2884 34636
rect 2940 31948 2996 34860
rect 3164 34850 3220 34860
rect 3276 35140 3332 35150
rect 3276 34802 3332 35084
rect 3276 34750 3278 34802
rect 3330 34750 3332 34802
rect 3276 34738 3332 34750
rect 3388 34580 3444 36316
rect 3164 34524 3444 34580
rect 2940 31892 3108 31948
rect 2940 30996 2996 31006
rect 2940 30902 2996 30940
rect 2828 27022 2830 27074
rect 2882 27022 2884 27074
rect 2828 27010 2884 27022
rect 2268 26964 2324 26974
rect 2156 26850 2212 26862
rect 2156 26798 2158 26850
rect 2210 26798 2212 26850
rect 2156 26292 2212 26798
rect 2156 26226 2212 26236
rect 1820 26180 1876 26190
rect 1820 25620 1876 26124
rect 2268 26178 2324 26908
rect 2940 26516 2996 26526
rect 3052 26516 3108 31892
rect 3164 30772 3220 34524
rect 3164 30706 3220 30716
rect 3276 32564 3332 32574
rect 3164 30324 3220 30334
rect 3164 30210 3220 30268
rect 3164 30158 3166 30210
rect 3218 30158 3220 30210
rect 3164 30146 3220 30158
rect 3276 26516 3332 32508
rect 2940 26514 3108 26516
rect 2940 26462 2942 26514
rect 2994 26462 3108 26514
rect 2940 26460 3108 26462
rect 3164 26460 3332 26516
rect 3500 26516 3556 37884
rect 3612 37874 3668 37884
rect 3612 37268 3668 37278
rect 3612 37174 3668 37212
rect 3612 37044 3668 37054
rect 3612 35810 3668 36988
rect 3612 35758 3614 35810
rect 3666 35758 3668 35810
rect 3612 35138 3668 35758
rect 3612 35086 3614 35138
rect 3666 35086 3668 35138
rect 3612 35074 3668 35086
rect 3724 36258 3780 36270
rect 3724 36206 3726 36258
rect 3778 36206 3780 36258
rect 3724 32564 3780 36206
rect 3836 35364 3892 38108
rect 3948 37938 4004 39676
rect 5628 39506 5684 40348
rect 5628 39454 5630 39506
rect 5682 39454 5684 39506
rect 5628 39442 5684 39454
rect 4844 39396 4900 39406
rect 4844 39394 5572 39396
rect 4844 39342 4846 39394
rect 4898 39342 5572 39394
rect 4844 39340 5572 39342
rect 4844 39330 4900 39340
rect 5516 39058 5572 39340
rect 5516 39006 5518 39058
rect 5570 39006 5572 39058
rect 5516 38994 5572 39006
rect 5740 39060 5796 40460
rect 5964 40514 6020 41022
rect 5964 40462 5966 40514
rect 6018 40462 6020 40514
rect 5964 40450 6020 40462
rect 5964 39506 6020 39518
rect 5964 39454 5966 39506
rect 6018 39454 6020 39506
rect 5964 39060 6020 39454
rect 5740 38994 5796 39004
rect 5852 39004 6020 39060
rect 4844 38948 4900 38958
rect 4844 38854 4900 38892
rect 4396 38836 4452 38846
rect 4284 38834 4452 38836
rect 4284 38782 4398 38834
rect 4450 38782 4452 38834
rect 4284 38780 4452 38782
rect 4172 38388 4228 38398
rect 3948 37886 3950 37938
rect 4002 37886 4004 37938
rect 3948 37874 4004 37886
rect 4060 38164 4116 38174
rect 3948 37378 4004 37390
rect 3948 37326 3950 37378
rect 4002 37326 4004 37378
rect 3948 36932 4004 37326
rect 3948 36866 4004 36876
rect 4060 36596 4116 38108
rect 3948 36540 4116 36596
rect 3948 35922 4004 36540
rect 4060 36372 4116 36382
rect 4060 36278 4116 36316
rect 3948 35870 3950 35922
rect 4002 35870 4004 35922
rect 3948 35858 4004 35870
rect 3836 35308 4004 35364
rect 3836 35138 3892 35150
rect 3836 35086 3838 35138
rect 3890 35086 3892 35138
rect 3836 35026 3892 35086
rect 3948 35140 4004 35308
rect 4172 35252 4228 38332
rect 4284 38052 4340 38780
rect 4396 38770 4452 38780
rect 5068 38836 5124 38846
rect 5068 38742 5124 38780
rect 5740 38834 5796 38846
rect 5740 38782 5742 38834
rect 5794 38782 5796 38834
rect 4956 38724 5012 38734
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4284 37996 4676 38052
rect 4396 37826 4452 37838
rect 4396 37774 4398 37826
rect 4450 37774 4452 37826
rect 4396 37492 4452 37774
rect 4396 37426 4452 37436
rect 4620 37490 4676 37996
rect 4732 37940 4788 37950
rect 4732 37846 4788 37884
rect 4620 37438 4622 37490
rect 4674 37438 4676 37490
rect 4620 37426 4676 37438
rect 4844 37492 4900 37502
rect 4172 35186 4228 35196
rect 4284 37266 4340 37278
rect 4284 37214 4286 37266
rect 4338 37214 4340 37266
rect 3948 35074 4004 35084
rect 3836 34974 3838 35026
rect 3890 34974 3892 35026
rect 3836 34962 3892 34974
rect 3724 32498 3780 32508
rect 3612 29986 3668 29998
rect 3612 29934 3614 29986
rect 3666 29934 3668 29986
rect 3612 29652 3668 29934
rect 3612 29586 3668 29596
rect 3612 26516 3668 26526
rect 3500 26514 3668 26516
rect 3500 26462 3614 26514
rect 3666 26462 3668 26514
rect 3500 26460 3668 26462
rect 2940 26450 2996 26460
rect 2268 26126 2270 26178
rect 2322 26126 2324 26178
rect 2268 26114 2324 26126
rect 1820 25554 1876 25564
rect 2940 25508 2996 25518
rect 3164 25508 3220 26460
rect 3612 26450 3668 26460
rect 3276 26290 3332 26302
rect 3276 26238 3278 26290
rect 3330 26238 3332 26290
rect 3276 26180 3332 26238
rect 3276 26114 3332 26124
rect 2940 25506 3220 25508
rect 2940 25454 2942 25506
rect 2994 25454 3220 25506
rect 2940 25452 3220 25454
rect 2940 25442 2996 25452
rect 2156 25282 2212 25294
rect 2156 25230 2158 25282
rect 2210 25230 2212 25282
rect 2156 24948 2212 25230
rect 2156 24882 2212 24892
rect 2940 24724 2996 24734
rect 2940 24630 2996 24668
rect 1932 24610 1988 24622
rect 1932 24558 1934 24610
rect 1986 24558 1988 24610
rect 1932 24276 1988 24558
rect 1932 24210 1988 24220
rect 1708 23826 1764 23838
rect 1708 23774 1710 23826
rect 1762 23774 1764 23826
rect 1708 23604 1764 23774
rect 2044 23828 2100 23838
rect 2044 23734 2100 23772
rect 4284 23828 4340 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4396 36484 4452 36494
rect 4396 35922 4452 36428
rect 4732 36372 4788 36382
rect 4844 36372 4900 37436
rect 4956 37378 5012 38668
rect 5516 38276 5572 38286
rect 5292 37940 5348 37950
rect 5292 37490 5348 37884
rect 5292 37438 5294 37490
rect 5346 37438 5348 37490
rect 5292 37426 5348 37438
rect 4956 37326 4958 37378
rect 5010 37326 5012 37378
rect 4956 37314 5012 37326
rect 5516 37268 5572 38220
rect 5628 37828 5684 37838
rect 5628 37734 5684 37772
rect 5740 37492 5796 38782
rect 5740 37426 5796 37436
rect 5516 37266 5796 37268
rect 5516 37214 5518 37266
rect 5570 37214 5796 37266
rect 5516 37212 5796 37214
rect 5516 37202 5572 37212
rect 5740 36594 5796 37212
rect 5740 36542 5742 36594
rect 5794 36542 5796 36594
rect 5740 36530 5796 36542
rect 4732 36370 4900 36372
rect 4732 36318 4734 36370
rect 4786 36318 4900 36370
rect 4732 36316 4900 36318
rect 4732 36306 4788 36316
rect 4396 35870 4398 35922
rect 4450 35870 4452 35922
rect 4396 35858 4452 35870
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4956 32676 5012 32686
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4956 31218 5012 32620
rect 5740 32676 5796 32686
rect 5740 32582 5796 32620
rect 5852 31332 5908 39004
rect 6076 38668 6132 43200
rect 6636 40402 6692 40414
rect 6636 40350 6638 40402
rect 6690 40350 6692 40402
rect 6636 39732 6692 40350
rect 6188 39676 6692 39732
rect 6188 39172 6244 39676
rect 6748 39620 6804 43200
rect 6972 39620 7028 39630
rect 6748 39618 7028 39620
rect 6748 39566 6974 39618
rect 7026 39566 7028 39618
rect 6748 39564 7028 39566
rect 6636 39506 6692 39518
rect 6636 39454 6638 39506
rect 6690 39454 6692 39506
rect 6300 39396 6356 39406
rect 6300 39394 6468 39396
rect 6300 39342 6302 39394
rect 6354 39342 6468 39394
rect 6300 39340 6468 39342
rect 6300 39330 6356 39340
rect 6188 39116 6356 39172
rect 6188 38948 6244 38958
rect 6188 38854 6244 38892
rect 6076 38612 6244 38668
rect 4956 31166 4958 31218
rect 5010 31166 5012 31218
rect 4956 31154 5012 31166
rect 5516 31276 5908 31332
rect 5964 37938 6020 37950
rect 5964 37886 5966 37938
rect 6018 37886 6020 37938
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5516 29316 5572 31276
rect 5740 31108 5796 31118
rect 5740 31106 5908 31108
rect 5740 31054 5742 31106
rect 5794 31054 5908 31106
rect 5740 31052 5908 31054
rect 5740 31042 5796 31052
rect 5740 30212 5796 30222
rect 5628 29428 5684 29438
rect 5740 29428 5796 30156
rect 5628 29426 5796 29428
rect 5628 29374 5630 29426
rect 5682 29374 5796 29426
rect 5628 29372 5796 29374
rect 5628 29362 5684 29372
rect 5516 29250 5572 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5740 28644 5796 29372
rect 5852 28980 5908 31052
rect 5964 30996 6020 37886
rect 6188 37492 6244 38612
rect 6300 37938 6356 39116
rect 6300 37886 6302 37938
rect 6354 37886 6356 37938
rect 6300 37874 6356 37886
rect 6300 37492 6356 37502
rect 6188 37490 6356 37492
rect 6188 37438 6302 37490
rect 6354 37438 6356 37490
rect 6188 37436 6356 37438
rect 6300 37426 6356 37436
rect 5964 30930 6020 30940
rect 6188 31444 6244 31454
rect 6076 30884 6132 30894
rect 6076 29426 6132 30828
rect 6076 29374 6078 29426
rect 6130 29374 6132 29426
rect 6076 29362 6132 29374
rect 5852 28914 5908 28924
rect 5628 28642 5796 28644
rect 5628 28590 5742 28642
rect 5794 28590 5796 28642
rect 5628 28588 5796 28590
rect 5628 27858 5684 28588
rect 5740 28578 5796 28588
rect 6188 28642 6244 31388
rect 6412 31108 6468 39340
rect 6412 31042 6468 31052
rect 6524 38834 6580 38846
rect 6524 38782 6526 38834
rect 6578 38782 6580 38834
rect 6524 29876 6580 38782
rect 6636 38164 6692 39454
rect 6860 39396 6916 39406
rect 6860 39058 6916 39340
rect 6860 39006 6862 39058
rect 6914 39006 6916 39058
rect 6860 38994 6916 39006
rect 6972 38668 7028 39564
rect 7308 39396 7364 39406
rect 6636 38098 6692 38108
rect 6860 38612 7028 38668
rect 7084 39394 7364 39396
rect 7084 39342 7310 39394
rect 7362 39342 7364 39394
rect 7084 39340 7364 39342
rect 6636 37938 6692 37950
rect 6636 37886 6638 37938
rect 6690 37886 6692 37938
rect 6636 37156 6692 37886
rect 6860 37492 6916 38612
rect 7084 38050 7140 39340
rect 7308 39330 7364 39340
rect 7308 39172 7364 39182
rect 7084 37998 7086 38050
rect 7138 37998 7140 38050
rect 7084 37986 7140 37998
rect 7196 38834 7252 38846
rect 7196 38782 7198 38834
rect 7250 38782 7252 38834
rect 6972 37492 7028 37502
rect 6860 37490 7028 37492
rect 6860 37438 6974 37490
rect 7026 37438 7028 37490
rect 6860 37436 7028 37438
rect 6972 37426 7028 37436
rect 6636 37090 6692 37100
rect 7196 33236 7252 38782
rect 7308 38836 7364 39116
rect 7420 39060 7476 43200
rect 8092 41748 8148 43200
rect 7868 41692 8148 41748
rect 7868 40514 7924 41692
rect 8764 41412 8820 43200
rect 8764 41356 9268 41412
rect 7868 40462 7870 40514
rect 7922 40462 7924 40514
rect 7868 40450 7924 40462
rect 8764 40402 8820 40414
rect 8764 40350 8766 40402
rect 8818 40350 8820 40402
rect 8428 40180 8484 40190
rect 7868 39618 7924 39630
rect 7868 39566 7870 39618
rect 7922 39566 7924 39618
rect 7644 39394 7700 39406
rect 7644 39342 7646 39394
rect 7698 39342 7700 39394
rect 7532 39060 7588 39070
rect 7420 39058 7588 39060
rect 7420 39006 7534 39058
rect 7586 39006 7588 39058
rect 7420 39004 7588 39006
rect 7532 38994 7588 39004
rect 7308 38780 7476 38836
rect 7308 38612 7364 38622
rect 7308 37938 7364 38556
rect 7308 37886 7310 37938
rect 7362 37886 7364 37938
rect 7308 37874 7364 37886
rect 7420 37490 7476 38780
rect 7644 38724 7700 39342
rect 7868 39172 7924 39566
rect 7868 39106 7924 39116
rect 8428 39618 8484 40124
rect 8428 39566 8430 39618
rect 8482 39566 8484 39618
rect 8428 39060 8484 39566
rect 8652 39396 8708 39406
rect 8428 38994 8484 39004
rect 8540 39394 8708 39396
rect 8540 39342 8654 39394
rect 8706 39342 8708 39394
rect 8540 39340 8708 39342
rect 8316 38948 8372 38958
rect 8316 38854 8372 38892
rect 8092 38836 8148 38846
rect 8540 38836 8596 39340
rect 8652 39330 8708 39340
rect 8652 39060 8708 39070
rect 8764 39060 8820 40350
rect 9212 39732 9268 41356
rect 9324 40514 9380 40526
rect 9324 40462 9326 40514
rect 9378 40462 9380 40514
rect 9324 39956 9380 40462
rect 9436 40292 9492 43200
rect 10108 41858 10164 43200
rect 10108 41806 10110 41858
rect 10162 41806 10164 41858
rect 10108 41794 10164 41806
rect 9548 41188 9604 41198
rect 9548 40404 9604 41132
rect 9548 40402 10276 40404
rect 9548 40350 9550 40402
rect 9602 40350 10276 40402
rect 9548 40348 10276 40350
rect 9548 40338 9604 40348
rect 9436 40226 9492 40236
rect 9324 39900 9604 39956
rect 9436 39732 9492 39742
rect 9212 39730 9492 39732
rect 9212 39678 9438 39730
rect 9490 39678 9492 39730
rect 9212 39676 9492 39678
rect 9436 39666 9492 39676
rect 8652 39058 8820 39060
rect 8652 39006 8654 39058
rect 8706 39006 8820 39058
rect 8652 39004 8820 39006
rect 8988 39394 9044 39406
rect 8988 39342 8990 39394
rect 9042 39342 9044 39394
rect 8652 38994 8708 39004
rect 8876 38836 8932 38846
rect 8540 38834 8932 38836
rect 8540 38782 8878 38834
rect 8930 38782 8932 38834
rect 8540 38780 8932 38782
rect 8092 38742 8148 38780
rect 8876 38770 8932 38780
rect 8988 38668 9044 39342
rect 7644 38658 7700 38668
rect 8428 38612 9044 38668
rect 8316 38276 8372 38286
rect 7980 38052 8036 38062
rect 7644 37940 7700 37950
rect 7644 37846 7700 37884
rect 7980 37938 8036 37996
rect 8316 38050 8372 38220
rect 8316 37998 8318 38050
rect 8370 37998 8372 38050
rect 8316 37986 8372 37998
rect 7980 37886 7982 37938
rect 8034 37886 8036 37938
rect 7980 37874 8036 37886
rect 7420 37438 7422 37490
rect 7474 37438 7476 37490
rect 7420 37426 7476 37438
rect 8428 37490 8484 38612
rect 9324 38500 9380 38510
rect 9100 38388 9156 38398
rect 9100 38050 9156 38332
rect 9100 37998 9102 38050
rect 9154 37998 9156 38050
rect 9100 37986 9156 37998
rect 9324 37938 9380 38444
rect 9324 37886 9326 37938
rect 9378 37886 9380 37938
rect 9324 37874 9380 37886
rect 8652 37828 8708 37838
rect 8652 37734 8708 37772
rect 8428 37438 8430 37490
rect 8482 37438 8484 37490
rect 8428 37426 8484 37438
rect 8204 37266 8260 37278
rect 8204 37214 8206 37266
rect 8258 37214 8260 37266
rect 8204 37156 8260 37214
rect 8204 37090 8260 37100
rect 8988 37156 9044 37166
rect 8988 37062 9044 37100
rect 9548 35812 9604 39900
rect 10220 39730 10276 40348
rect 10220 39678 10222 39730
rect 10274 39678 10276 39730
rect 10220 39666 10276 39678
rect 10332 40402 10388 40414
rect 10332 40350 10334 40402
rect 10386 40350 10388 40402
rect 9996 39396 10052 39406
rect 9660 39060 9716 39070
rect 9660 38966 9716 39004
rect 9772 38164 9828 38174
rect 9772 38050 9828 38108
rect 9772 37998 9774 38050
rect 9826 37998 9828 38050
rect 9772 37986 9828 37998
rect 9996 37938 10052 39340
rect 10220 38724 10276 38734
rect 10220 38630 10276 38668
rect 9996 37886 9998 37938
rect 10050 37886 10052 37938
rect 9996 37874 10052 37886
rect 10332 37938 10388 40350
rect 10556 40292 10612 40302
rect 10556 39506 10612 40236
rect 10556 39454 10558 39506
rect 10610 39454 10612 39506
rect 10556 39442 10612 39454
rect 10780 39508 10836 43200
rect 11452 41972 11508 43200
rect 11452 41916 11956 41972
rect 11228 41858 11284 41870
rect 11228 41806 11230 41858
rect 11282 41806 11284 41858
rect 11228 40514 11284 41806
rect 11900 40626 11956 41916
rect 11900 40574 11902 40626
rect 11954 40574 11956 40626
rect 11900 40562 11956 40574
rect 12124 40628 12180 43200
rect 12796 41972 12852 43200
rect 12796 41916 13188 41972
rect 12348 40628 12404 40638
rect 12124 40626 12404 40628
rect 12124 40574 12350 40626
rect 12402 40574 12404 40626
rect 12124 40572 12404 40574
rect 12348 40562 12404 40572
rect 13132 40626 13188 41916
rect 13132 40574 13134 40626
rect 13186 40574 13188 40626
rect 13132 40562 13188 40574
rect 13468 40628 13524 43200
rect 13692 40628 13748 40638
rect 13468 40626 13748 40628
rect 13468 40574 13694 40626
rect 13746 40574 13748 40626
rect 13468 40572 13748 40574
rect 14140 40628 14196 43200
rect 14252 40628 14308 40638
rect 14140 40626 14308 40628
rect 14140 40574 14254 40626
rect 14306 40574 14308 40626
rect 14140 40572 14308 40574
rect 13692 40562 13748 40572
rect 14252 40562 14308 40572
rect 14812 40626 14868 43200
rect 15484 41298 15540 43200
rect 15484 41246 15486 41298
rect 15538 41246 15540 41298
rect 15484 41234 15540 41246
rect 16044 41298 16100 41310
rect 16044 41246 16046 41298
rect 16098 41246 16100 41298
rect 14812 40574 14814 40626
rect 14866 40574 14868 40626
rect 14812 40562 14868 40574
rect 11228 40462 11230 40514
rect 11282 40462 11284 40514
rect 11228 40450 11284 40462
rect 16044 40514 16100 41246
rect 16044 40462 16046 40514
rect 16098 40462 16100 40514
rect 16044 40450 16100 40462
rect 15148 40402 15204 40414
rect 15148 40350 15150 40402
rect 15202 40350 15204 40402
rect 11004 39508 11060 39518
rect 10780 39506 11060 39508
rect 10780 39454 11006 39506
rect 11058 39454 11060 39506
rect 10780 39452 11060 39454
rect 11004 39442 11060 39452
rect 10668 39172 10724 39182
rect 10668 38050 10724 39116
rect 15148 38500 15204 40350
rect 16156 39844 16212 43200
rect 16828 41076 16884 43200
rect 16828 41020 17332 41076
rect 17052 40514 17108 40526
rect 17052 40462 17054 40514
rect 17106 40462 17108 40514
rect 16156 39778 16212 39788
rect 16828 39844 16884 39854
rect 16828 39730 16884 39788
rect 16828 39678 16830 39730
rect 16882 39678 16884 39730
rect 16828 39666 16884 39678
rect 16380 39396 16436 39406
rect 16380 39302 16436 39340
rect 17052 39172 17108 40462
rect 17276 40404 17332 41020
rect 17500 40628 17556 43200
rect 17724 40628 17780 40638
rect 17500 40626 17780 40628
rect 17500 40574 17726 40626
rect 17778 40574 17780 40626
rect 17500 40572 17780 40574
rect 17724 40562 17780 40572
rect 18172 40628 18228 43200
rect 18172 40562 18228 40572
rect 17276 40402 17668 40404
rect 17276 40350 17278 40402
rect 17330 40350 17668 40402
rect 17276 40348 17668 40350
rect 17276 40338 17332 40348
rect 17612 39730 17668 40348
rect 17612 39678 17614 39730
rect 17666 39678 17668 39730
rect 17612 39666 17668 39678
rect 18508 40402 18564 40414
rect 18508 40350 18510 40402
rect 18562 40350 18564 40402
rect 17052 39106 17108 39116
rect 15148 38434 15204 38444
rect 10668 37998 10670 38050
rect 10722 37998 10724 38050
rect 10668 37986 10724 37998
rect 10332 37886 10334 37938
rect 10386 37886 10388 37938
rect 10332 37874 10388 37886
rect 18508 37828 18564 40350
rect 18844 39732 18900 43200
rect 19180 40628 19236 40638
rect 19516 40628 19572 43200
rect 20188 41300 20244 43200
rect 20188 41244 20468 41300
rect 20188 40962 20244 40974
rect 20188 40910 20190 40962
rect 20242 40910 20244 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19852 40628 19908 40638
rect 19516 40572 19852 40628
rect 19180 40534 19236 40572
rect 19852 40534 19908 40572
rect 20188 40626 20244 40910
rect 20188 40574 20190 40626
rect 20242 40574 20244 40626
rect 20188 40562 20244 40574
rect 18844 39730 19348 39732
rect 18844 39678 18846 39730
rect 18898 39678 19348 39730
rect 18844 39676 19348 39678
rect 18844 39666 18900 39676
rect 19292 39618 19348 39676
rect 19292 39566 19294 39618
rect 19346 39566 19348 39618
rect 19292 39554 19348 39566
rect 20412 39506 20468 41244
rect 20860 40962 20916 43200
rect 20860 40910 20862 40962
rect 20914 40910 20916 40962
rect 20860 40898 20916 40910
rect 21532 41076 21588 43200
rect 21532 41020 22036 41076
rect 20972 40628 21028 40638
rect 20412 39454 20414 39506
rect 20466 39454 20468 39506
rect 20412 39442 20468 39454
rect 20748 40514 20804 40526
rect 20748 40462 20750 40514
rect 20802 40462 20804 40514
rect 19068 39394 19124 39406
rect 19068 39342 19070 39394
rect 19122 39342 19124 39394
rect 19068 38388 19124 39342
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19068 38322 19124 38332
rect 20748 38276 20804 40462
rect 20972 40402 21028 40572
rect 20972 40350 20974 40402
rect 21026 40350 21028 40402
rect 20972 40338 21028 40350
rect 21532 39730 21588 41020
rect 21532 39678 21534 39730
rect 21586 39678 21588 39730
rect 21532 39666 21588 39678
rect 21756 40514 21812 40526
rect 21756 40462 21758 40514
rect 21810 40462 21812 40514
rect 20748 38210 20804 38220
rect 21756 38164 21812 40462
rect 21980 40402 22036 41020
rect 22204 41074 22260 43200
rect 22204 41022 22206 41074
rect 22258 41022 22260 41074
rect 22204 41010 22260 41022
rect 22876 40964 22932 43200
rect 23324 41074 23380 41086
rect 23324 41022 23326 41074
rect 23378 41022 23380 41074
rect 22876 40908 23156 40964
rect 21980 40350 21982 40402
rect 22034 40350 22036 40402
rect 21980 40338 22036 40350
rect 22428 40402 22484 40414
rect 22428 40350 22430 40402
rect 22482 40350 22484 40402
rect 21756 38098 21812 38108
rect 22428 38052 22484 40350
rect 22876 39732 22932 39742
rect 22876 39638 22932 39676
rect 23100 39506 23156 40908
rect 23324 40514 23380 41022
rect 23548 40740 23604 43200
rect 24220 41748 24276 43200
rect 24220 41692 24836 41748
rect 23548 40684 24052 40740
rect 23324 40462 23326 40514
rect 23378 40462 23380 40514
rect 23324 40450 23380 40462
rect 23996 39732 24052 40684
rect 23996 39618 24052 39676
rect 23996 39566 23998 39618
rect 24050 39566 24052 39618
rect 23996 39554 24052 39566
rect 24556 40402 24612 40414
rect 24556 40350 24558 40402
rect 24610 40350 24612 40402
rect 23100 39454 23102 39506
rect 23154 39454 23156 39506
rect 23100 39442 23156 39454
rect 22428 37986 22484 37996
rect 23772 39394 23828 39406
rect 23772 39342 23774 39394
rect 23826 39342 23828 39394
rect 23772 37940 23828 39342
rect 24556 38948 24612 40350
rect 24780 40292 24836 41692
rect 24892 40516 24948 43200
rect 24892 40460 25172 40516
rect 25004 40292 25060 40302
rect 24780 40290 25060 40292
rect 24780 40238 25006 40290
rect 25058 40238 25060 40290
rect 24780 40236 25060 40238
rect 25004 40226 25060 40236
rect 25116 40292 25172 40460
rect 25116 40226 25172 40236
rect 25564 39732 25620 43200
rect 26236 40516 26292 43200
rect 26908 43092 26964 43200
rect 27244 43092 27300 43260
rect 26908 43036 27300 43092
rect 26236 40460 26740 40516
rect 25788 40404 25844 40414
rect 26124 40404 26180 40414
rect 25788 40402 26180 40404
rect 25788 40350 25790 40402
rect 25842 40350 26126 40402
rect 26178 40350 26180 40402
rect 25788 40348 26180 40350
rect 25788 40338 25844 40348
rect 25564 39730 26068 39732
rect 25564 39678 25566 39730
rect 25618 39678 26068 39730
rect 25564 39676 26068 39678
rect 25564 39666 25620 39676
rect 26012 39618 26068 39676
rect 26012 39566 26014 39618
rect 26066 39566 26068 39618
rect 26012 39554 26068 39566
rect 24556 38882 24612 38892
rect 25788 39394 25844 39406
rect 25788 39342 25790 39394
rect 25842 39342 25844 39394
rect 23772 37874 23828 37884
rect 18508 37762 18564 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 25788 37156 25844 39342
rect 26124 38612 26180 40348
rect 26236 39058 26292 40460
rect 26572 40292 26628 40302
rect 26572 40198 26628 40236
rect 26684 39618 26740 40460
rect 27580 39730 27636 43260
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 27580 39678 27582 39730
rect 27634 39678 27636 39730
rect 27580 39666 27636 39678
rect 26684 39566 26686 39618
rect 26738 39566 26740 39618
rect 26684 39554 26740 39566
rect 26236 39006 26238 39058
rect 26290 39006 26292 39058
rect 26236 38994 26292 39006
rect 26460 39394 26516 39406
rect 26460 39342 26462 39394
rect 26514 39342 26516 39394
rect 26460 38724 26516 39342
rect 27132 39394 27188 39406
rect 27132 39342 27134 39394
rect 27186 39342 27188 39394
rect 26460 38658 26516 38668
rect 26796 38724 26852 38734
rect 27132 38724 27188 39342
rect 26796 38722 27188 38724
rect 26796 38670 26798 38722
rect 26850 38670 27188 38722
rect 26796 38668 27188 38670
rect 26124 38546 26180 38556
rect 25788 37090 25844 37100
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 9548 35746 9604 35756
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 16268 34242 16324 34254
rect 16268 34190 16270 34242
rect 16322 34190 16324 34242
rect 15036 34018 15092 34030
rect 15036 33966 15038 34018
rect 15090 33966 15092 34018
rect 7196 33170 7252 33180
rect 8764 33458 8820 33470
rect 8764 33406 8766 33458
rect 8818 33406 8820 33458
rect 6860 32450 6916 32462
rect 6860 32398 6862 32450
rect 6914 32398 6916 32450
rect 6860 30884 6916 32398
rect 8092 31892 8148 31902
rect 8652 31892 8708 31902
rect 8092 30994 8148 31836
rect 8092 30942 8094 30994
rect 8146 30942 8148 30994
rect 8092 30930 8148 30942
rect 8204 31890 8708 31892
rect 8204 31838 8654 31890
rect 8706 31838 8708 31890
rect 8204 31836 8708 31838
rect 6860 30818 6916 30828
rect 7756 30212 7812 30222
rect 7756 30118 7812 30156
rect 8204 30210 8260 31836
rect 8652 31826 8708 31836
rect 8428 31554 8484 31566
rect 8428 31502 8430 31554
rect 8482 31502 8484 31554
rect 8428 31220 8484 31502
rect 8764 31444 8820 33406
rect 14028 33460 14084 33470
rect 9772 33236 9828 33246
rect 8764 31378 8820 31388
rect 9100 33234 9828 33236
rect 9100 33182 9774 33234
rect 9826 33182 9828 33234
rect 9100 33180 9828 33182
rect 8988 31220 9044 31230
rect 8428 31164 8988 31220
rect 8652 30994 8708 31164
rect 8988 31126 9044 31164
rect 8652 30942 8654 30994
rect 8706 30942 8708 30994
rect 8204 30158 8206 30210
rect 8258 30158 8260 30210
rect 8204 30146 8260 30158
rect 8316 30884 8372 30894
rect 6524 29810 6580 29820
rect 8316 29650 8372 30828
rect 8652 30212 8708 30942
rect 8652 30146 8708 30156
rect 8316 29598 8318 29650
rect 8370 29598 8372 29650
rect 8316 29586 8372 29598
rect 8764 30100 8820 30110
rect 6188 28590 6190 28642
rect 6242 28590 6244 28642
rect 6188 28578 6244 28590
rect 6972 28980 7028 28990
rect 5628 27806 5630 27858
rect 5682 27806 5684 27858
rect 5628 27794 5684 27806
rect 6076 27858 6132 27870
rect 6076 27806 6078 27858
rect 6130 27806 6132 27858
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 6076 27188 6132 27806
rect 6076 27122 6132 27132
rect 6860 27188 6916 27198
rect 6860 27094 6916 27132
rect 6188 27076 6244 27086
rect 5404 26964 5460 26974
rect 5404 26514 5460 26908
rect 5404 26462 5406 26514
rect 5458 26462 5460 26514
rect 5404 26450 5460 26462
rect 6188 26514 6244 27020
rect 6188 26462 6190 26514
rect 6242 26462 6244 26514
rect 6188 26450 6244 26462
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 6972 25618 7028 28924
rect 8652 28420 8708 28430
rect 8764 28420 8820 30044
rect 9100 29650 9156 33180
rect 9772 33170 9828 33180
rect 9884 32674 9940 32686
rect 9884 32622 9886 32674
rect 9938 32622 9940 32674
rect 9772 31666 9828 31678
rect 9772 31614 9774 31666
rect 9826 31614 9828 31666
rect 9660 31220 9716 31230
rect 9436 30772 9492 30782
rect 9100 29598 9102 29650
rect 9154 29598 9156 29650
rect 9100 29586 9156 29598
rect 9212 30770 9492 30772
rect 9212 30718 9438 30770
rect 9490 30718 9492 30770
rect 9212 30716 9492 30718
rect 8652 28418 8820 28420
rect 8652 28366 8654 28418
rect 8706 28366 8820 28418
rect 8652 28364 8820 28366
rect 9100 29428 9156 29438
rect 8652 28354 8708 28364
rect 9100 28082 9156 29372
rect 9212 28866 9268 30716
rect 9436 30706 9492 30716
rect 9212 28814 9214 28866
rect 9266 28814 9268 28866
rect 9212 28802 9268 28814
rect 9660 29652 9716 31164
rect 9772 30770 9828 31614
rect 9772 30718 9774 30770
rect 9826 30718 9828 30770
rect 9772 30706 9828 30718
rect 9100 28030 9102 28082
rect 9154 28030 9156 28082
rect 9100 28018 9156 28030
rect 9548 28644 9604 28654
rect 9660 28644 9716 29596
rect 9548 28642 9716 28644
rect 9548 28590 9550 28642
rect 9602 28590 9716 28642
rect 9548 28588 9716 28590
rect 9772 30548 9828 30558
rect 9772 28644 9828 30492
rect 9884 29428 9940 32622
rect 10892 32450 10948 32462
rect 10892 32398 10894 32450
rect 10946 32398 10948 32450
rect 10332 30994 10388 31006
rect 10332 30942 10334 30994
rect 10386 30942 10388 30994
rect 10108 30884 10164 30894
rect 10108 30790 10164 30828
rect 9884 29362 9940 29372
rect 10332 30212 10388 30942
rect 10780 30884 10836 30894
rect 10332 29426 10388 30156
rect 10668 30882 10836 30884
rect 10668 30830 10782 30882
rect 10834 30830 10836 30882
rect 10668 30828 10836 30830
rect 10668 29986 10724 30828
rect 10780 30818 10836 30828
rect 10892 30548 10948 32398
rect 11676 31892 11732 31902
rect 11676 31890 12180 31892
rect 11676 31838 11678 31890
rect 11730 31838 12180 31890
rect 11676 31836 12180 31838
rect 11676 31826 11732 31836
rect 11228 31554 11284 31566
rect 11228 31502 11230 31554
rect 11282 31502 11284 31554
rect 11228 31220 11284 31502
rect 11228 31154 11284 31164
rect 11676 31220 11732 31230
rect 10892 30482 10948 30492
rect 11004 30994 11060 31006
rect 11004 30942 11006 30994
rect 11058 30942 11060 30994
rect 11004 30212 11060 30942
rect 11676 30994 11732 31164
rect 11676 30942 11678 30994
rect 11730 30942 11732 30994
rect 11676 30930 11732 30942
rect 12124 30994 12180 31836
rect 12796 31668 12852 31678
rect 12796 31666 13076 31668
rect 12796 31614 12798 31666
rect 12850 31614 13076 31666
rect 12796 31612 13076 31614
rect 12796 31602 12852 31612
rect 12124 30942 12126 30994
rect 12178 30942 12180 30994
rect 12124 30930 12180 30942
rect 11004 30146 11060 30156
rect 11676 30212 11732 30222
rect 11676 30118 11732 30156
rect 12572 30212 12628 30222
rect 11452 30100 11508 30110
rect 11452 30006 11508 30044
rect 12348 30098 12404 30110
rect 12348 30046 12350 30098
rect 12402 30046 12404 30098
rect 10668 29934 10670 29986
rect 10722 29934 10724 29986
rect 10668 29922 10724 29934
rect 11228 29986 11284 29998
rect 11228 29934 11230 29986
rect 11282 29934 11284 29986
rect 10332 29374 10334 29426
rect 10386 29374 10388 29426
rect 10108 29316 10164 29326
rect 9996 29314 10164 29316
rect 9996 29262 10110 29314
rect 10162 29262 10164 29314
rect 9996 29260 10164 29262
rect 9884 28644 9940 28654
rect 9772 28642 9940 28644
rect 9772 28590 9886 28642
rect 9938 28590 9940 28642
rect 9772 28588 9940 28590
rect 8316 27970 8372 27982
rect 8316 27918 8318 27970
rect 8370 27918 8372 27970
rect 7868 26964 7924 27002
rect 7868 26898 7924 26908
rect 6972 25566 6974 25618
rect 7026 25566 7028 25618
rect 6972 25554 7028 25566
rect 7308 26852 7364 26862
rect 7308 25618 7364 26796
rect 8316 26516 8372 27918
rect 8652 27076 8708 27086
rect 8652 26962 8708 27020
rect 8652 26910 8654 26962
rect 8706 26910 8708 26962
rect 8652 26898 8708 26910
rect 8876 27074 8932 27086
rect 8876 27022 8878 27074
rect 8930 27022 8932 27074
rect 8876 26964 8932 27022
rect 9548 26908 9604 28588
rect 9884 28578 9940 28588
rect 9884 28420 9940 28430
rect 9884 27970 9940 28364
rect 9884 27918 9886 27970
rect 9938 27918 9940 27970
rect 9884 27906 9940 27918
rect 8876 26898 8932 26908
rect 9212 26852 9268 26862
rect 9212 26758 9268 26796
rect 9324 26852 9604 26908
rect 9996 26962 10052 29260
rect 10108 29250 10164 29260
rect 9996 26910 9998 26962
rect 10050 26910 10052 26962
rect 9996 26898 10052 26910
rect 10108 26964 10164 26974
rect 10332 26964 10388 29374
rect 10668 29652 10724 29662
rect 10668 29426 10724 29596
rect 10668 29374 10670 29426
rect 10722 29374 10724 29426
rect 10668 29362 10724 29374
rect 11228 28644 11284 29934
rect 12236 29652 12292 29662
rect 11228 28578 11284 28588
rect 11340 29426 11396 29438
rect 11340 29374 11342 29426
rect 11394 29374 11396 29426
rect 11228 27746 11284 27758
rect 11228 27694 11230 27746
rect 11282 27694 11284 27746
rect 11228 27076 11284 27694
rect 11228 27010 11284 27020
rect 10164 26908 10388 26964
rect 11340 26908 11396 29374
rect 12236 28082 12292 29596
rect 12348 28418 12404 30046
rect 12572 28756 12628 30156
rect 13020 28866 13076 31612
rect 13468 30212 13524 30222
rect 13020 28814 13022 28866
rect 13074 28814 13076 28866
rect 13020 28802 13076 28814
rect 13132 30100 13188 30110
rect 12572 28690 12628 28700
rect 12348 28366 12350 28418
rect 12402 28366 12404 28418
rect 12348 28354 12404 28366
rect 12236 28030 12238 28082
rect 12290 28030 12292 28082
rect 12236 28018 12292 28030
rect 12684 27858 12740 27870
rect 12684 27806 12686 27858
rect 12738 27806 12740 27858
rect 12236 27076 12292 27086
rect 12236 26982 12292 27020
rect 12684 27074 12740 27806
rect 13132 27858 13188 30044
rect 13468 28756 13524 30156
rect 14028 30210 14084 33404
rect 14924 32450 14980 32462
rect 14924 32398 14926 32450
rect 14978 32398 14980 32450
rect 14588 31554 14644 31566
rect 14588 31502 14590 31554
rect 14642 31502 14644 31554
rect 14588 31220 14644 31502
rect 14588 31154 14644 31164
rect 14700 31220 14756 31230
rect 14700 31218 14868 31220
rect 14700 31166 14702 31218
rect 14754 31166 14868 31218
rect 14700 31164 14868 31166
rect 14700 31154 14756 31164
rect 14028 30158 14030 30210
rect 14082 30158 14084 30210
rect 14028 30146 14084 30158
rect 14364 30548 14420 30558
rect 13692 29650 13748 29662
rect 13692 29598 13694 29650
rect 13746 29598 13748 29650
rect 13132 27806 13134 27858
rect 13186 27806 13188 27858
rect 13132 27794 13188 27806
rect 13356 28700 13524 28756
rect 13580 28756 13636 28766
rect 12684 27022 12686 27074
rect 12738 27022 12740 27074
rect 12684 26908 12740 27022
rect 8316 26450 8372 26460
rect 8540 26740 8596 26750
rect 8540 26290 8596 26684
rect 9324 26628 9380 26852
rect 8540 26238 8542 26290
rect 8594 26238 8596 26290
rect 8540 26226 8596 26238
rect 9100 26572 9604 26628
rect 9100 26290 9156 26572
rect 9100 26238 9102 26290
rect 9154 26238 9156 26290
rect 9100 26226 9156 26238
rect 9324 25730 9380 25742
rect 9324 25678 9326 25730
rect 9378 25678 9380 25730
rect 7308 25566 7310 25618
rect 7362 25566 7364 25618
rect 7308 25554 7364 25566
rect 9100 25620 9156 25630
rect 9324 25620 9380 25678
rect 9100 25618 9380 25620
rect 9100 25566 9102 25618
rect 9154 25566 9380 25618
rect 9100 25564 9380 25566
rect 9548 25618 9604 26572
rect 9772 26404 9828 26414
rect 9772 26310 9828 26348
rect 10108 26402 10164 26908
rect 10108 26350 10110 26402
rect 10162 26350 10164 26402
rect 10108 26338 10164 26350
rect 10556 26852 10612 26862
rect 11340 26852 11844 26908
rect 12684 26852 13076 26908
rect 10556 26402 10612 26796
rect 10556 26350 10558 26402
rect 10610 26350 10612 26402
rect 10556 26338 10612 26350
rect 11788 26178 11844 26852
rect 13020 26292 13076 26852
rect 13356 26292 13412 28700
rect 13580 28642 13636 28700
rect 13692 28754 13748 29598
rect 14364 29650 14420 30492
rect 14812 29876 14868 31164
rect 14924 30100 14980 32398
rect 15036 31892 15092 33966
rect 15148 33460 15204 33470
rect 15148 33366 15204 33404
rect 16156 33236 16212 33246
rect 15036 31826 15092 31836
rect 15260 33234 16212 33236
rect 15260 33182 16158 33234
rect 16210 33182 16212 33234
rect 15260 33180 16212 33182
rect 15260 31218 15316 33180
rect 16156 33170 16212 33180
rect 15932 32674 15988 32686
rect 15932 32622 15934 32674
rect 15986 32622 15988 32674
rect 15708 31778 15764 31790
rect 15708 31726 15710 31778
rect 15762 31726 15764 31778
rect 15260 31166 15262 31218
rect 15314 31166 15316 31218
rect 15260 31154 15316 31166
rect 15596 31220 15652 31230
rect 15596 31126 15652 31164
rect 15708 30212 15764 31726
rect 15932 30548 15988 32622
rect 16268 31948 16324 34190
rect 19740 34242 19796 34254
rect 19740 34190 19742 34242
rect 19794 34190 19796 34242
rect 18732 34018 18788 34030
rect 18732 33966 18734 34018
rect 18786 33966 18788 34018
rect 18396 33460 18452 33470
rect 18396 33458 18564 33460
rect 18396 33406 18398 33458
rect 18450 33406 18564 33458
rect 18396 33404 18564 33406
rect 18396 33394 18452 33404
rect 15932 30482 15988 30492
rect 16044 31892 16324 31948
rect 17052 33234 17108 33246
rect 17052 33182 17054 33234
rect 17106 33182 17108 33234
rect 15708 30146 15764 30156
rect 14924 30034 14980 30044
rect 14812 29820 15092 29876
rect 14364 29598 14366 29650
rect 14418 29598 14420 29650
rect 14364 29586 14420 29598
rect 15036 29650 15092 29820
rect 15036 29598 15038 29650
rect 15090 29598 15092 29650
rect 15036 29586 15092 29598
rect 14924 29314 14980 29326
rect 14924 29262 14926 29314
rect 14978 29262 14980 29314
rect 13692 28702 13694 28754
rect 13746 28702 13748 28754
rect 13692 28690 13748 28702
rect 14140 28756 14196 28766
rect 13580 28590 13582 28642
rect 13634 28590 13636 28642
rect 13580 28578 13636 28590
rect 13020 26290 13412 26292
rect 13020 26238 13022 26290
rect 13074 26238 13358 26290
rect 13410 26238 13412 26290
rect 13020 26236 13412 26238
rect 13020 26226 13076 26236
rect 13356 26226 13412 26236
rect 13916 28084 13972 28094
rect 13916 26290 13972 28028
rect 14140 27186 14196 28700
rect 14924 28756 14980 29262
rect 14924 28690 14980 28700
rect 15820 29202 15876 29214
rect 15820 29150 15822 29202
rect 15874 29150 15876 29202
rect 14476 28530 14532 28542
rect 14476 28478 14478 28530
rect 14530 28478 14532 28530
rect 14476 27972 14532 28478
rect 15036 28420 15092 28430
rect 14476 27906 14532 27916
rect 14924 28418 15092 28420
rect 14924 28366 15038 28418
rect 15090 28366 15092 28418
rect 14924 28364 15092 28366
rect 14140 27134 14142 27186
rect 14194 27134 14196 27186
rect 14140 27122 14196 27134
rect 14924 27076 14980 28364
rect 15036 28354 15092 28364
rect 14924 26982 14980 27020
rect 15596 28082 15652 28094
rect 15596 28030 15598 28082
rect 15650 28030 15652 28082
rect 15596 26628 15652 28030
rect 15596 26562 15652 26572
rect 13916 26238 13918 26290
rect 13970 26238 13972 26290
rect 13916 26226 13972 26238
rect 11788 26126 11790 26178
rect 11842 26126 11844 26178
rect 11788 26114 11844 26126
rect 9548 25566 9550 25618
rect 9602 25566 9604 25618
rect 9100 25554 9156 25564
rect 8092 25394 8148 25406
rect 8092 25342 8094 25394
rect 8146 25342 8148 25394
rect 7532 24834 7588 24846
rect 7532 24782 7534 24834
rect 7586 24782 7588 24834
rect 6188 24610 6244 24622
rect 6188 24558 6190 24610
rect 6242 24558 6244 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23762 4340 23772
rect 4732 23828 4788 23838
rect 1708 23538 1764 23548
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 2044 23492 2100 23502
rect 1596 22930 1652 22942
rect 1596 22878 1598 22930
rect 1650 22878 1652 22930
rect 1596 20692 1652 22878
rect 1708 22932 1764 22942
rect 1708 22484 1764 22876
rect 1708 22370 1764 22428
rect 1708 22318 1710 22370
rect 1762 22318 1764 22370
rect 1708 22306 1764 22318
rect 2044 22258 2100 23436
rect 2044 22206 2046 22258
rect 2098 22206 2100 22258
rect 2044 22194 2100 22206
rect 2380 23266 2436 23278
rect 2380 23214 2382 23266
rect 2434 23214 2436 23266
rect 2380 21700 2436 23214
rect 4732 23154 4788 23772
rect 6188 23828 6244 24558
rect 6188 23762 6244 23772
rect 7420 23716 7476 23726
rect 6972 23714 7476 23716
rect 6972 23662 7422 23714
rect 7474 23662 7476 23714
rect 6972 23660 7476 23662
rect 6972 23266 7028 23660
rect 7420 23650 7476 23660
rect 6972 23214 6974 23266
rect 7026 23214 7028 23266
rect 6972 23202 7028 23214
rect 4732 23102 4734 23154
rect 4786 23102 4788 23154
rect 4732 23090 4788 23102
rect 5292 23154 5348 23166
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 5292 23044 5348 23102
rect 5628 23044 5684 23054
rect 5292 23042 5684 23044
rect 5292 22990 5630 23042
rect 5682 22990 5684 23042
rect 5292 22988 5684 22990
rect 5292 22820 5348 22830
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2492 22484 2548 22494
rect 2492 22390 2548 22428
rect 4844 22260 4900 22270
rect 2380 21634 2436 21644
rect 3500 21700 3556 21710
rect 4508 21700 4564 21710
rect 1820 21588 1876 21598
rect 2156 21588 2212 21598
rect 1820 21494 1876 21532
rect 2044 21586 2212 21588
rect 2044 21534 2158 21586
rect 2210 21534 2212 21586
rect 2044 21532 2212 21534
rect 1708 20916 1764 20926
rect 1708 20804 1764 20860
rect 1708 20802 1876 20804
rect 1708 20750 1710 20802
rect 1762 20750 1876 20802
rect 1708 20748 1876 20750
rect 1708 20738 1764 20748
rect 1596 20626 1652 20636
rect 1820 20242 1876 20748
rect 2044 20690 2100 21532
rect 2156 21522 2212 21532
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 2044 20626 2100 20638
rect 2716 20692 2772 20702
rect 2716 20598 2772 20636
rect 1820 20190 1822 20242
rect 1874 20190 1876 20242
rect 1820 20178 1876 20190
rect 3388 20356 3444 20366
rect 3388 20018 3444 20300
rect 3388 19966 3390 20018
rect 3442 19966 3444 20018
rect 3052 19122 3108 19134
rect 3052 19070 3054 19122
rect 3106 19070 3108 19122
rect 3052 18674 3108 19070
rect 3052 18622 3054 18674
rect 3106 18622 3108 18674
rect 3052 18610 3108 18622
rect 2380 18450 2436 18462
rect 2380 18398 2382 18450
rect 2434 18398 2436 18450
rect 2268 18338 2324 18350
rect 2268 18286 2270 18338
rect 2322 18286 2324 18338
rect 2156 17442 2212 17454
rect 2156 17390 2158 17442
rect 2210 17390 2212 17442
rect 2156 17106 2212 17390
rect 2156 17054 2158 17106
rect 2210 17054 2212 17106
rect 2156 17042 2212 17054
rect 1596 16660 1652 16670
rect 1596 16658 1988 16660
rect 1596 16606 1598 16658
rect 1650 16606 1988 16658
rect 1596 16604 1988 16606
rect 1596 16594 1652 16604
rect 1932 15426 1988 16604
rect 1932 15374 1934 15426
rect 1986 15374 1988 15426
rect 1932 15362 1988 15374
rect 1596 14420 1652 14430
rect 1596 13970 1652 14364
rect 1596 13918 1598 13970
rect 1650 13918 1652 13970
rect 1596 13906 1652 13918
rect 2268 13970 2324 18286
rect 2380 17668 2436 18398
rect 2380 17574 2436 17612
rect 3388 17668 3444 19966
rect 3500 17778 3556 21644
rect 3612 21698 4564 21700
rect 3612 21646 4510 21698
rect 4562 21646 4564 21698
rect 3612 21644 4564 21646
rect 3612 20242 3668 21644
rect 4508 21634 4564 21644
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3612 20190 3614 20242
rect 3666 20190 3668 20242
rect 3612 20178 3668 20190
rect 3836 20914 3892 20926
rect 3836 20862 3838 20914
rect 3890 20862 3892 20914
rect 3836 18900 3892 20862
rect 4844 20804 4900 22204
rect 5292 21810 5348 22764
rect 5292 21758 5294 21810
rect 5346 21758 5348 21810
rect 5292 21746 5348 21758
rect 5628 21588 5684 22988
rect 7532 22820 7588 24782
rect 8092 23716 8148 25342
rect 9548 24836 9604 25566
rect 8092 23650 8148 23660
rect 8204 23714 8260 23726
rect 8204 23662 8206 23714
rect 8258 23662 8260 23714
rect 7532 22754 7588 22764
rect 7980 23042 8036 23054
rect 7980 22990 7982 23042
rect 8034 22990 8036 23042
rect 7084 22260 7140 22270
rect 7084 22166 7140 22204
rect 6972 22036 7028 22046
rect 6972 21698 7028 21980
rect 6972 21646 6974 21698
rect 7026 21646 7028 21698
rect 6972 21634 7028 21646
rect 7980 21700 8036 22990
rect 8092 22484 8148 22494
rect 8092 22390 8148 22428
rect 8204 22148 8260 23662
rect 8204 22082 8260 22092
rect 9436 23716 9492 23726
rect 9436 21810 9492 23660
rect 9548 22370 9604 24780
rect 9548 22318 9550 22370
rect 9602 22318 9604 22370
rect 9548 21924 9604 22318
rect 9660 25730 9716 25742
rect 9660 25678 9662 25730
rect 9714 25678 9716 25730
rect 9660 22372 9716 25678
rect 11452 25620 11508 25630
rect 10556 25618 11508 25620
rect 10556 25566 11454 25618
rect 11506 25566 11508 25618
rect 10556 25564 11508 25566
rect 10444 24836 10500 24846
rect 10444 24742 10500 24780
rect 10556 23938 10612 25564
rect 11452 25554 11508 25564
rect 15484 25620 15540 25630
rect 12796 25394 12852 25406
rect 12796 25342 12798 25394
rect 12850 25342 12852 25394
rect 10556 23886 10558 23938
rect 10610 23886 10612 23938
rect 10556 23874 10612 23886
rect 10892 24836 10948 24846
rect 10892 23940 10948 24780
rect 10892 23938 11284 23940
rect 10892 23886 10894 23938
rect 10946 23886 11284 23938
rect 10892 23884 11284 23886
rect 10892 23874 10948 23884
rect 11228 23604 11284 23884
rect 11564 23828 11620 23838
rect 11900 23828 11956 23838
rect 11228 23378 11284 23548
rect 11228 23326 11230 23378
rect 11282 23326 11284 23378
rect 11228 23314 11284 23326
rect 11340 23826 11620 23828
rect 11340 23774 11566 23826
rect 11618 23774 11620 23826
rect 11340 23772 11620 23774
rect 11340 22708 11396 23772
rect 11564 23762 11620 23772
rect 11676 23772 11900 23828
rect 11676 23268 11732 23772
rect 11900 23734 11956 23772
rect 12348 23828 12404 23838
rect 12348 23734 12404 23772
rect 12796 23716 12852 25342
rect 15484 24722 15540 25564
rect 15820 24836 15876 29150
rect 15932 28868 15988 28878
rect 16044 28868 16100 31892
rect 16156 31780 16212 31790
rect 16156 31686 16212 31724
rect 17052 30210 17108 33182
rect 17276 33124 17332 33134
rect 17276 31218 17332 33068
rect 18396 31556 18452 31566
rect 18396 31462 18452 31500
rect 17276 31166 17278 31218
rect 17330 31166 17332 31218
rect 17276 31154 17332 31166
rect 17836 31108 17892 31118
rect 17052 30158 17054 30210
rect 17106 30158 17108 30210
rect 17052 30146 17108 30158
rect 17388 30212 17444 30222
rect 17444 30156 17556 30212
rect 17388 30118 17444 30156
rect 16492 29986 16548 29998
rect 16492 29934 16494 29986
rect 16546 29934 16548 29986
rect 15932 28866 16100 28868
rect 15932 28814 15934 28866
rect 15986 28814 16100 28866
rect 15932 28812 16100 28814
rect 16156 29540 16212 29550
rect 15932 28802 15988 28812
rect 16156 28082 16212 29484
rect 16156 28030 16158 28082
rect 16210 28030 16212 28082
rect 16156 28018 16212 28030
rect 16492 27970 16548 29934
rect 16716 29988 16772 29998
rect 16492 27918 16494 27970
rect 16546 27918 16548 27970
rect 16492 27906 16548 27918
rect 16604 29426 16660 29438
rect 16604 29374 16606 29426
rect 16658 29374 16660 29426
rect 16156 27860 16212 27870
rect 16156 27076 16212 27804
rect 16604 27860 16660 29374
rect 16716 28530 16772 29932
rect 16716 28478 16718 28530
rect 16770 28478 16772 28530
rect 16716 28466 16772 28478
rect 17500 29316 17556 30156
rect 17836 30210 17892 31052
rect 17836 30158 17838 30210
rect 17890 30158 17892 30210
rect 17836 30146 17892 30158
rect 18060 31106 18116 31118
rect 18060 31054 18062 31106
rect 18114 31054 18116 31106
rect 16828 28420 16884 28430
rect 16828 27970 16884 28364
rect 16828 27918 16830 27970
rect 16882 27918 16884 27970
rect 16828 27906 16884 27918
rect 17500 28082 17556 29260
rect 17948 29316 18004 29326
rect 17948 29222 18004 29260
rect 18060 28756 18116 31054
rect 18060 28690 18116 28700
rect 18396 29314 18452 29326
rect 18396 29262 18398 29314
rect 18450 29262 18452 29314
rect 17500 28030 17502 28082
rect 17554 28030 17556 28082
rect 16604 27794 16660 27804
rect 16156 26982 16212 27020
rect 17164 26964 17220 26974
rect 17052 26908 17164 26964
rect 16380 26514 16436 26526
rect 16380 26462 16382 26514
rect 16434 26462 16436 26514
rect 16268 25620 16324 25630
rect 16268 25506 16324 25564
rect 16268 25454 16270 25506
rect 16322 25454 16324 25506
rect 16268 25442 16324 25454
rect 16380 24948 16436 26462
rect 16940 26404 16996 26414
rect 16940 26310 16996 26348
rect 16380 24882 16436 24892
rect 16604 25620 16660 25630
rect 16604 24946 16660 25564
rect 16604 24894 16606 24946
rect 16658 24894 16660 24946
rect 16604 24882 16660 24894
rect 15876 24780 15988 24836
rect 15820 24742 15876 24780
rect 15484 24670 15486 24722
rect 15538 24670 15540 24722
rect 15484 24658 15540 24670
rect 15260 24050 15316 24062
rect 15260 23998 15262 24050
rect 15314 23998 15316 24050
rect 12796 23650 12852 23660
rect 14252 23826 14308 23838
rect 14252 23774 14254 23826
rect 14306 23774 14308 23826
rect 13356 23604 13412 23614
rect 10220 22652 11396 22708
rect 11452 23212 11732 23268
rect 12572 23268 12628 23278
rect 9884 22372 9940 22382
rect 9660 22370 9940 22372
rect 9660 22318 9886 22370
rect 9938 22318 9940 22370
rect 9660 22316 9940 22318
rect 9884 22306 9940 22316
rect 9548 21858 9604 21868
rect 9436 21758 9438 21810
rect 9490 21758 9492 21810
rect 9436 21746 9492 21758
rect 10220 21810 10276 22652
rect 10668 22148 10724 22158
rect 10724 22092 10836 22148
rect 10668 22082 10724 22092
rect 10220 21758 10222 21810
rect 10274 21758 10276 21810
rect 10220 21746 10276 21758
rect 10668 21924 10724 21934
rect 7980 21634 8036 21644
rect 5628 21494 5684 21532
rect 6748 21588 6804 21598
rect 4844 20738 4900 20748
rect 6188 20802 6244 20814
rect 6188 20750 6190 20802
rect 6242 20750 6244 20802
rect 5964 20578 6020 20590
rect 5964 20526 5966 20578
rect 6018 20526 6020 20578
rect 4060 20356 4116 20366
rect 4060 20018 4116 20300
rect 5852 20244 5908 20254
rect 5964 20244 6020 20526
rect 6188 20356 6244 20750
rect 6748 20802 6804 21532
rect 7980 21476 8036 21486
rect 7980 21382 8036 21420
rect 6748 20750 6750 20802
rect 6802 20750 6804 20802
rect 6748 20738 6804 20750
rect 7308 20802 7364 20814
rect 7308 20750 7310 20802
rect 7362 20750 7364 20802
rect 6188 20290 6244 20300
rect 5852 20242 6020 20244
rect 5852 20190 5854 20242
rect 5906 20190 6020 20242
rect 5852 20188 6020 20190
rect 5852 20178 5908 20188
rect 4060 19966 4062 20018
rect 4114 19966 4116 20018
rect 4060 19954 4116 19966
rect 4172 19796 4228 19806
rect 3836 18834 3892 18844
rect 3948 19794 4228 19796
rect 3948 19742 4174 19794
rect 4226 19742 4228 19794
rect 3948 19740 4228 19742
rect 3836 18676 3892 18686
rect 3948 18676 4004 19740
rect 4172 19730 4228 19740
rect 5068 19794 5124 19806
rect 5068 19742 5070 19794
rect 5122 19742 5124 19794
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4060 19348 4116 19358
rect 4060 19254 4116 19292
rect 5068 19124 5124 19742
rect 7308 19346 7364 20750
rect 9660 20578 9716 20590
rect 9660 20526 9662 20578
rect 9714 20526 9716 20578
rect 7308 19294 7310 19346
rect 7362 19294 7364 19346
rect 7308 19282 7364 19294
rect 7756 20132 7812 20142
rect 6188 19124 6244 19134
rect 5068 19122 6244 19124
rect 5068 19070 6190 19122
rect 6242 19070 6244 19122
rect 5068 19068 6244 19070
rect 6188 19058 6244 19068
rect 7084 19012 7140 19022
rect 3836 18674 4004 18676
rect 3836 18622 3838 18674
rect 3890 18622 4004 18674
rect 3836 18620 4004 18622
rect 6076 18900 6132 18910
rect 3836 18610 3892 18620
rect 6076 18450 6132 18844
rect 6524 18452 6580 18462
rect 6076 18398 6078 18450
rect 6130 18398 6132 18450
rect 6076 18386 6132 18398
rect 6300 18450 6580 18452
rect 6300 18398 6526 18450
rect 6578 18398 6580 18450
rect 6300 18396 6580 18398
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 3500 17726 3502 17778
rect 3554 17726 3556 17778
rect 3500 17714 3556 17726
rect 6300 17778 6356 18396
rect 6524 18386 6580 18396
rect 6300 17726 6302 17778
rect 6354 17726 6356 17778
rect 3388 17556 3444 17612
rect 4732 17668 4788 17678
rect 4732 17574 4788 17612
rect 3388 17500 3556 17556
rect 3052 15988 3108 15998
rect 3052 15894 3108 15932
rect 3276 15204 3332 15214
rect 3276 15202 3444 15204
rect 3276 15150 3278 15202
rect 3330 15150 3444 15202
rect 3276 15148 3444 15150
rect 3276 15138 3332 15148
rect 2716 14420 2772 14430
rect 2716 14326 2772 14364
rect 2268 13918 2270 13970
rect 2322 13918 2324 13970
rect 2268 13906 2324 13918
rect 3388 13748 3444 15148
rect 3500 14420 3556 17500
rect 4956 17442 5012 17454
rect 4956 17390 4958 17442
rect 5010 17390 5012 17442
rect 4732 16882 4788 16894
rect 4732 16830 4734 16882
rect 4786 16830 4788 16882
rect 4732 16772 4788 16830
rect 4732 16706 4788 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4956 16436 5012 17390
rect 5628 17108 5684 17118
rect 5292 17052 5628 17108
rect 5292 16884 5348 17052
rect 5628 17014 5684 17052
rect 6300 17108 6356 17726
rect 7084 17554 7140 18956
rect 7532 18452 7588 18462
rect 7532 17668 7588 18396
rect 7756 18338 7812 20076
rect 9660 20132 9716 20526
rect 9660 20066 9716 20076
rect 10444 20578 10500 20590
rect 10444 20526 10446 20578
rect 10498 20526 10500 20578
rect 8092 20018 8148 20030
rect 8092 19966 8094 20018
rect 8146 19966 8148 20018
rect 8092 19348 8148 19966
rect 8764 20018 8820 20030
rect 8764 19966 8766 20018
rect 8818 19966 8820 20018
rect 8764 19908 8820 19966
rect 9772 19908 9828 19918
rect 8764 19906 9828 19908
rect 8764 19854 9774 19906
rect 9826 19854 9828 19906
rect 8764 19852 9828 19854
rect 8092 19282 8148 19292
rect 8764 19012 8820 19022
rect 9324 19012 9380 19022
rect 8764 18918 8820 18956
rect 8876 19010 9380 19012
rect 8876 18958 9326 19010
rect 9378 18958 9380 19010
rect 8876 18956 9380 18958
rect 8876 18674 8932 18956
rect 9324 18946 9380 18956
rect 8876 18622 8878 18674
rect 8930 18622 8932 18674
rect 8876 18610 8932 18622
rect 7756 18286 7758 18338
rect 7810 18286 7812 18338
rect 7756 18274 7812 18286
rect 8988 18450 9044 18462
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 18340 9044 18398
rect 8988 18274 9044 18284
rect 8876 18228 8932 18238
rect 8092 17780 8148 17790
rect 8092 17686 8148 17724
rect 7532 17602 7588 17612
rect 7084 17502 7086 17554
rect 7138 17502 7140 17554
rect 7084 17490 7140 17502
rect 6356 17052 6468 17108
rect 6300 17042 6356 17052
rect 4956 16370 5012 16380
rect 5180 16882 5348 16884
rect 5180 16830 5294 16882
rect 5346 16830 5348 16882
rect 5180 16828 5348 16830
rect 4060 16210 4116 16222
rect 4060 16158 4062 16210
rect 4114 16158 4116 16210
rect 3948 16100 4004 16110
rect 3948 14642 4004 16044
rect 4060 15316 4116 16158
rect 5180 15540 5236 16828
rect 5292 16818 5348 16828
rect 5516 15988 5572 15998
rect 5516 15894 5572 15932
rect 4060 15250 4116 15260
rect 4732 15484 5236 15540
rect 4732 15314 4788 15484
rect 4732 15262 4734 15314
rect 4786 15262 4788 15314
rect 4732 15250 4788 15262
rect 5068 15316 5124 15326
rect 5068 15222 5124 15260
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 3948 14590 3950 14642
rect 4002 14590 4004 14642
rect 3948 14578 4004 14590
rect 3500 14364 4004 14420
rect 3388 13682 3444 13692
rect 3948 12962 4004 14364
rect 5180 13972 5236 15484
rect 6076 15874 6132 15886
rect 6076 15822 6078 15874
rect 6130 15822 6132 15874
rect 5628 13972 5684 13982
rect 5180 13970 5684 13972
rect 5180 13918 5630 13970
rect 5682 13918 5684 13970
rect 5180 13916 5684 13918
rect 4620 13748 4676 13758
rect 4620 13654 4676 13692
rect 5180 13746 5236 13916
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 5180 13682 5236 13694
rect 4172 13524 4228 13534
rect 4172 13186 4228 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4172 13134 4174 13186
rect 4226 13134 4228 13186
rect 4172 13122 4228 13134
rect 3948 12910 3950 12962
rect 4002 12910 4004 12962
rect 3948 12898 4004 12910
rect 5628 12178 5684 13916
rect 6076 13524 6132 15822
rect 6412 14644 6468 17052
rect 8876 16994 8932 18172
rect 8876 16942 8878 16994
rect 8930 16942 8932 16994
rect 8876 16930 8932 16942
rect 9548 17668 9604 17678
rect 9772 17668 9828 19852
rect 10332 18562 10388 18574
rect 10332 18510 10334 18562
rect 10386 18510 10388 18562
rect 10332 17892 10388 18510
rect 10332 17826 10388 17836
rect 9548 17666 9828 17668
rect 9548 17614 9550 17666
rect 9602 17614 9828 17666
rect 9548 17612 9828 17614
rect 9884 17668 9940 17678
rect 9548 16996 9604 17612
rect 9884 17574 9940 17612
rect 7532 16772 7588 16782
rect 7532 16678 7588 16716
rect 7420 16436 7476 16446
rect 7420 15538 7476 16380
rect 8540 16100 8596 16110
rect 8540 16006 8596 16044
rect 9212 16098 9268 16110
rect 9212 16046 9214 16098
rect 9266 16046 9268 16098
rect 9212 15876 9268 16046
rect 9548 15876 9604 16940
rect 10444 15988 10500 20526
rect 10668 20130 10724 21868
rect 10780 20914 10836 22092
rect 10780 20862 10782 20914
rect 10834 20862 10836 20914
rect 10780 20850 10836 20862
rect 11004 20916 11060 20926
rect 11452 20916 11508 23212
rect 12572 23174 12628 23212
rect 11788 22930 11844 22942
rect 11788 22878 11790 22930
rect 11842 22878 11844 22930
rect 11788 22260 11844 22878
rect 13356 22484 13412 23548
rect 13580 22484 13636 22494
rect 13132 22482 13636 22484
rect 13132 22430 13582 22482
rect 13634 22430 13636 22482
rect 13132 22428 13636 22430
rect 11788 22194 11844 22204
rect 12460 22260 12516 22270
rect 12460 22146 12516 22204
rect 12460 22094 12462 22146
rect 12514 22094 12516 22146
rect 12460 22082 12516 22094
rect 13020 22148 13076 22158
rect 13020 22054 13076 22092
rect 12460 21588 12516 21598
rect 13132 21588 13188 22428
rect 13580 22418 13636 22428
rect 13804 22484 13860 22494
rect 13804 22036 13860 22428
rect 14252 22484 14308 23774
rect 14252 22418 14308 22428
rect 14588 23268 14644 23278
rect 14588 22482 14644 23212
rect 14924 23156 14980 23166
rect 14924 23154 15092 23156
rect 14924 23102 14926 23154
rect 14978 23102 15092 23154
rect 14924 23100 15092 23102
rect 14924 23090 14980 23100
rect 14588 22430 14590 22482
rect 14642 22430 14644 22482
rect 14588 22418 14644 22430
rect 14924 22932 14980 22942
rect 14924 22482 14980 22876
rect 14924 22430 14926 22482
rect 14978 22430 14980 22482
rect 13916 22260 13972 22270
rect 13916 22166 13972 22204
rect 14252 22260 14308 22270
rect 14252 22166 14308 22204
rect 14924 22260 14980 22430
rect 14924 22194 14980 22204
rect 13804 21980 13972 22036
rect 12460 21494 12516 21532
rect 12908 21586 13188 21588
rect 12908 21534 13134 21586
rect 13186 21534 13188 21586
rect 12908 21532 13188 21534
rect 11004 20914 11508 20916
rect 11004 20862 11006 20914
rect 11058 20862 11454 20914
rect 11506 20862 11508 20914
rect 11004 20860 11508 20862
rect 11004 20850 11060 20860
rect 11452 20850 11508 20860
rect 12908 20914 12964 21532
rect 13132 21522 13188 21532
rect 13468 21588 13524 21598
rect 13804 21588 13860 21598
rect 13468 21586 13636 21588
rect 13468 21534 13470 21586
rect 13522 21534 13636 21586
rect 13468 21532 13636 21534
rect 13468 21522 13524 21532
rect 12908 20862 12910 20914
rect 12962 20862 12964 20914
rect 12908 20850 12964 20862
rect 10668 20078 10670 20130
rect 10722 20078 10724 20130
rect 10668 20066 10724 20078
rect 13580 20802 13636 21532
rect 13580 20750 13582 20802
rect 13634 20750 13636 20802
rect 13580 20244 13636 20750
rect 11900 19906 11956 19918
rect 11900 19854 11902 19906
rect 11954 19854 11956 19906
rect 11788 19234 11844 19246
rect 11788 19182 11790 19234
rect 11842 19182 11844 19234
rect 11340 18452 11396 18462
rect 11340 18338 11396 18396
rect 11340 18286 11342 18338
rect 11394 18286 11396 18338
rect 11340 18274 11396 18286
rect 10556 16996 10612 17006
rect 10556 16902 10612 16940
rect 11788 16210 11844 19182
rect 11900 18340 11956 19854
rect 12460 19234 12516 19246
rect 12460 19182 12462 19234
rect 12514 19182 12516 19234
rect 12460 19012 12516 19182
rect 13580 19234 13636 20188
rect 13580 19182 13582 19234
rect 13634 19182 13636 19234
rect 13580 19170 13636 19182
rect 13692 21586 13860 21588
rect 13692 21534 13806 21586
rect 13858 21534 13860 21586
rect 13692 21532 13860 21534
rect 12796 19012 12852 19022
rect 12460 19010 12852 19012
rect 12460 18958 12798 19010
rect 12850 18958 12852 19010
rect 12460 18956 12852 18958
rect 11900 18274 11956 18284
rect 12572 18228 12628 18238
rect 12572 18134 12628 18172
rect 12460 17442 12516 17454
rect 12460 17390 12462 17442
rect 12514 17390 12516 17442
rect 12460 16324 12516 17390
rect 12796 16996 12852 18956
rect 13244 18674 13300 18686
rect 13244 18622 13246 18674
rect 13298 18622 13300 18674
rect 13020 17892 13076 17902
rect 13020 17798 13076 17836
rect 13244 17892 13300 18622
rect 13244 17826 13300 17836
rect 12796 16930 12852 16940
rect 13580 17442 13636 17454
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13580 16996 13636 17390
rect 13580 16930 13636 16940
rect 12460 16258 12516 16268
rect 13580 16324 13636 16334
rect 13580 16230 13636 16268
rect 11788 16158 11790 16210
rect 11842 16158 11844 16210
rect 11788 16146 11844 16158
rect 10556 15988 10612 15998
rect 10444 15986 10612 15988
rect 10444 15934 10558 15986
rect 10610 15934 10612 15986
rect 10444 15932 10612 15934
rect 10556 15922 10612 15932
rect 9212 15874 9604 15876
rect 9212 15822 9550 15874
rect 9602 15822 9604 15874
rect 9212 15820 9604 15822
rect 7420 15486 7422 15538
rect 7474 15486 7476 15538
rect 7420 15474 7476 15486
rect 8540 15202 8596 15214
rect 8540 15150 8542 15202
rect 8594 15150 8596 15202
rect 8204 15092 8260 15102
rect 8204 15090 8484 15092
rect 8204 15038 8206 15090
rect 8258 15038 8484 15090
rect 8204 15036 8484 15038
rect 8204 15026 8260 15036
rect 6412 14530 6468 14588
rect 6412 14478 6414 14530
rect 6466 14478 6468 14530
rect 6412 14466 6468 14478
rect 7084 14530 7140 14542
rect 7084 14478 7086 14530
rect 7138 14478 7140 14530
rect 7084 13636 7140 14478
rect 8428 13860 8484 15036
rect 8540 14644 8596 15150
rect 8540 14578 8596 14588
rect 9548 14644 9604 15820
rect 13244 15540 13300 15550
rect 9548 14578 9604 14588
rect 10332 14812 10612 14868
rect 10108 14420 10164 14430
rect 10108 14326 10164 14364
rect 9548 14306 9604 14318
rect 9548 14254 9550 14306
rect 9602 14254 9604 14306
rect 8540 13860 8596 13870
rect 8428 13858 8596 13860
rect 8428 13806 8542 13858
rect 8594 13806 8596 13858
rect 8428 13804 8596 13806
rect 8540 13794 8596 13804
rect 7532 13636 7588 13646
rect 7084 13634 7588 13636
rect 7084 13582 7534 13634
rect 7586 13582 7588 13634
rect 7084 13580 7588 13582
rect 7532 13570 7588 13580
rect 6076 13458 6132 13468
rect 9324 13188 9380 13198
rect 6972 12964 7028 12974
rect 6972 12870 7028 12908
rect 8540 12964 8596 12974
rect 6860 12740 6916 12750
rect 6860 12646 6916 12684
rect 7196 12738 7252 12750
rect 7196 12686 7198 12738
rect 7250 12686 7252 12738
rect 5628 12126 5630 12178
rect 5682 12126 5684 12178
rect 5628 12114 5684 12126
rect 6076 12178 6132 12190
rect 6076 12126 6078 12178
rect 6130 12126 6132 12178
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 6076 11508 6132 12126
rect 6076 11442 6132 11452
rect 7196 11284 7252 12686
rect 7756 12740 7812 12750
rect 7756 12646 7812 12684
rect 8316 12290 8372 12302
rect 8316 12238 8318 12290
rect 8370 12238 8372 12290
rect 7644 11508 7700 11518
rect 7644 11414 7700 11452
rect 7196 11218 7252 11228
rect 8316 10834 8372 12238
rect 8316 10782 8318 10834
rect 8370 10782 8372 10834
rect 8316 10770 8372 10782
rect 8540 10610 8596 12908
rect 9100 11954 9156 11966
rect 9100 11902 9102 11954
rect 9154 11902 9156 11954
rect 8652 11284 8708 11294
rect 8652 11190 8708 11228
rect 9100 10724 9156 11902
rect 9324 11618 9380 13132
rect 9548 12404 9604 14254
rect 9884 12964 9940 12974
rect 9772 12740 9828 12750
rect 9660 12404 9716 12414
rect 9548 12402 9716 12404
rect 9548 12350 9662 12402
rect 9714 12350 9716 12402
rect 9548 12348 9716 12350
rect 9660 12338 9716 12348
rect 9324 11566 9326 11618
rect 9378 11566 9380 11618
rect 9324 11554 9380 11566
rect 9100 10658 9156 10668
rect 8540 10558 8542 10610
rect 8594 10558 8596 10610
rect 8540 10546 8596 10558
rect 9660 10500 9716 10510
rect 9772 10500 9828 12684
rect 9884 12180 9940 12908
rect 10332 12962 10388 14812
rect 10332 12910 10334 12962
rect 10386 12910 10388 12962
rect 10332 12898 10388 12910
rect 10444 14644 10500 14654
rect 10556 14644 10612 14812
rect 11340 14644 11396 14654
rect 10556 14642 11396 14644
rect 10556 14590 11342 14642
rect 11394 14590 11396 14642
rect 10556 14588 11396 14590
rect 10444 14306 10500 14588
rect 11340 14578 11396 14588
rect 12348 14420 12404 14430
rect 12348 14326 12404 14364
rect 10444 14254 10446 14306
rect 10498 14254 10500 14306
rect 10444 12964 10500 14254
rect 13244 13972 13300 15484
rect 13692 14980 13748 21532
rect 13804 21522 13860 21532
rect 13804 21364 13860 21374
rect 13804 19236 13860 21308
rect 13916 20802 13972 21980
rect 15036 21476 15092 23100
rect 15260 22372 15316 23998
rect 15372 23716 15428 23726
rect 15372 22932 15428 23660
rect 15708 23714 15764 23726
rect 15708 23662 15710 23714
rect 15762 23662 15764 23714
rect 15708 23492 15764 23662
rect 15484 23436 15708 23492
rect 15484 23154 15540 23436
rect 15708 23426 15764 23436
rect 15484 23102 15486 23154
rect 15538 23102 15540 23154
rect 15484 23090 15540 23102
rect 15932 23266 15988 24780
rect 16156 24612 16212 24622
rect 16156 24610 16436 24612
rect 16156 24558 16158 24610
rect 16210 24558 16436 24610
rect 16156 24556 16436 24558
rect 16156 24546 16212 24556
rect 16268 23268 16324 23278
rect 15932 23214 15934 23266
rect 15986 23214 15988 23266
rect 15932 22932 15988 23214
rect 15372 22876 15764 22932
rect 15708 22594 15764 22876
rect 15932 22866 15988 22876
rect 16156 23212 16268 23268
rect 15708 22542 15710 22594
rect 15762 22542 15764 22594
rect 15708 22530 15764 22542
rect 15260 22306 15316 22316
rect 16156 21810 16212 23212
rect 16268 23202 16324 23212
rect 16156 21758 16158 21810
rect 16210 21758 16212 21810
rect 16156 21746 16212 21758
rect 16268 23042 16324 23054
rect 16268 22990 16270 23042
rect 16322 22990 16324 23042
rect 15036 21410 15092 21420
rect 13916 20750 13918 20802
rect 13970 20750 13972 20802
rect 13916 20738 13972 20750
rect 16268 20690 16324 22990
rect 16268 20638 16270 20690
rect 16322 20638 16324 20690
rect 16268 20626 16324 20638
rect 14812 20018 14868 20030
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19908 14868 19966
rect 15260 19908 15316 19918
rect 14812 19852 15260 19908
rect 13916 19236 13972 19246
rect 13804 19234 13972 19236
rect 13804 19182 13918 19234
rect 13970 19182 13972 19234
rect 13804 19180 13972 19182
rect 13916 19170 13972 19180
rect 14028 17892 14084 17902
rect 14028 17798 14084 17836
rect 13916 17666 13972 17678
rect 13916 17614 13918 17666
rect 13970 17614 13972 17666
rect 13804 16100 13860 16110
rect 13916 16100 13972 17614
rect 13804 16098 13972 16100
rect 13804 16046 13806 16098
rect 13858 16046 13972 16098
rect 13804 16044 13972 16046
rect 13804 15540 13860 16044
rect 13804 15474 13860 15484
rect 15148 15316 15204 15326
rect 15260 15316 15316 19852
rect 16380 19010 16436 24556
rect 16492 23938 16548 23950
rect 16492 23886 16494 23938
rect 16546 23886 16548 23938
rect 16492 23492 16548 23886
rect 16492 23426 16548 23436
rect 17052 23828 17108 26908
rect 17164 26898 17220 26908
rect 17500 26514 17556 28030
rect 18396 28084 18452 29262
rect 18508 28644 18564 33404
rect 18732 31108 18788 33966
rect 19740 33124 19796 34190
rect 26236 34018 26292 34030
rect 26236 33966 26238 34018
rect 26290 33966 26292 34018
rect 24780 33572 24836 33582
rect 19740 33058 19796 33068
rect 24556 33458 24612 33470
rect 24556 33406 24558 33458
rect 24610 33406 24612 33458
rect 23996 33012 24052 33022
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19180 32676 19236 32686
rect 19180 31890 19236 32620
rect 20076 32676 20132 32686
rect 20076 32582 20132 32620
rect 19404 32450 19460 32462
rect 19404 32398 19406 32450
rect 19458 32398 19460 32450
rect 19404 31948 19460 32398
rect 21196 32450 21252 32462
rect 21196 32398 21198 32450
rect 21250 32398 21252 32450
rect 21196 31948 21252 32398
rect 19404 31892 19572 31948
rect 19180 31838 19182 31890
rect 19234 31838 19236 31890
rect 19180 31826 19236 31838
rect 18732 31042 18788 31052
rect 19404 31666 19460 31678
rect 19404 31614 19406 31666
rect 19458 31614 19460 31666
rect 19404 29988 19460 31614
rect 19404 29922 19460 29932
rect 19404 29540 19460 29550
rect 19404 29446 19460 29484
rect 19516 29316 19572 31892
rect 20524 31892 21252 31948
rect 20300 31780 20356 31790
rect 20188 31778 20356 31780
rect 20188 31726 20302 31778
rect 20354 31726 20356 31778
rect 20188 31724 20356 31726
rect 19740 31668 19796 31678
rect 20188 31668 20244 31724
rect 20300 31714 20356 31724
rect 19740 31666 20244 31668
rect 19740 31614 19742 31666
rect 19794 31614 20244 31666
rect 19740 31612 20244 31614
rect 19740 31602 19796 31612
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 29988 20244 31612
rect 20300 31556 20356 31566
rect 20300 31462 20356 31500
rect 20412 30996 20468 31006
rect 20524 30996 20580 31892
rect 23324 31778 23380 31790
rect 23324 31726 23326 31778
rect 23378 31726 23380 31778
rect 21420 31554 21476 31566
rect 21420 31502 21422 31554
rect 21474 31502 21476 31554
rect 20412 30994 20580 30996
rect 20412 30942 20414 30994
rect 20466 30942 20580 30994
rect 20412 30940 20580 30942
rect 20748 30996 20804 31006
rect 21084 30996 21140 31006
rect 21420 30996 21476 31502
rect 20748 30994 21476 30996
rect 20748 30942 20750 30994
rect 20802 30942 21086 30994
rect 21138 30942 21476 30994
rect 20748 30940 21476 30942
rect 21756 30994 21812 31006
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 20412 30930 20468 30940
rect 20188 29922 20244 29932
rect 20300 30100 20356 30110
rect 20300 29986 20356 30044
rect 20300 29934 20302 29986
rect 20354 29934 20356 29986
rect 20300 29922 20356 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18956 28644 19012 28654
rect 18508 28642 19012 28644
rect 18508 28590 18958 28642
rect 19010 28590 19012 28642
rect 18508 28588 19012 28590
rect 18956 28578 19012 28588
rect 19516 28644 19572 29260
rect 20524 29428 20580 29438
rect 20748 29428 20804 30940
rect 21084 30930 21140 30940
rect 21756 30884 21812 30942
rect 21756 30818 21812 30828
rect 21756 30210 21812 30222
rect 21756 30158 21758 30210
rect 21810 30158 21812 30210
rect 21532 30100 21588 30110
rect 21532 30006 21588 30044
rect 21756 30100 21812 30158
rect 21756 30034 21812 30044
rect 22204 30212 22260 30222
rect 20524 29426 20804 29428
rect 20524 29374 20526 29426
rect 20578 29374 20804 29426
rect 20524 29372 20804 29374
rect 20860 29986 20916 29998
rect 20860 29934 20862 29986
rect 20914 29934 20916 29986
rect 19852 28756 19908 28766
rect 19852 28662 19908 28700
rect 20524 28756 20580 29372
rect 20524 28690 20580 28700
rect 19516 28550 19572 28588
rect 20636 28644 20692 28654
rect 20636 28550 20692 28588
rect 20188 28532 20244 28542
rect 20188 28438 20244 28476
rect 20860 28532 20916 29934
rect 21196 29988 21252 29998
rect 21084 29426 21140 29438
rect 21084 29374 21086 29426
rect 21138 29374 21140 29426
rect 21084 29092 21140 29374
rect 21084 29026 21140 29036
rect 20860 28466 20916 28476
rect 21196 28420 21252 29932
rect 22204 28756 22260 30156
rect 22764 30210 22820 30222
rect 22764 30158 22766 30210
rect 22818 30158 22820 30210
rect 22764 29764 22820 30158
rect 23324 30212 23380 31726
rect 23996 31778 24052 32956
rect 24332 32450 24388 32462
rect 24332 32398 24334 32450
rect 24386 32398 24388 32450
rect 24332 31948 24388 32398
rect 23996 31726 23998 31778
rect 24050 31726 24052 31778
rect 23996 31714 24052 31726
rect 24220 31892 24388 31948
rect 24220 31218 24276 31892
rect 24556 31780 24612 33406
rect 24556 31714 24612 31724
rect 24668 32452 24724 32462
rect 24220 31166 24222 31218
rect 24274 31166 24276 31218
rect 24220 31154 24276 31166
rect 23324 30146 23380 30156
rect 22764 29698 22820 29708
rect 24668 30100 24724 32396
rect 24780 31218 24836 33516
rect 24780 31166 24782 31218
rect 24834 31166 24836 31218
rect 24780 31154 24836 31166
rect 25676 33234 25732 33246
rect 25676 33182 25678 33234
rect 25730 33182 25732 33234
rect 25676 31220 25732 33182
rect 26236 33012 26292 33966
rect 26236 32946 26292 32956
rect 26348 33460 26404 33470
rect 26012 32452 26068 32462
rect 26012 32358 26068 32396
rect 26236 32450 26292 32462
rect 26236 32398 26238 32450
rect 26290 32398 26292 32450
rect 26236 31666 26292 32398
rect 26236 31614 26238 31666
rect 26290 31614 26292 31666
rect 26236 31602 26292 31614
rect 25676 31154 25732 31164
rect 25676 30994 25732 31006
rect 25676 30942 25678 30994
rect 25730 30942 25732 30994
rect 25340 30884 25396 30894
rect 25676 30884 25732 30942
rect 26348 30994 26404 33404
rect 26796 31948 26852 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 40684 36596 40740 36606
rect 40572 36594 40740 36596
rect 40572 36542 40686 36594
rect 40738 36542 40740 36594
rect 40572 36540 40740 36542
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 40348 35026 40404 35038
rect 40348 34974 40350 35026
rect 40402 34974 40404 35026
rect 39116 34804 39172 34814
rect 38556 34802 39172 34804
rect 38556 34750 39118 34802
rect 39170 34750 39172 34802
rect 38556 34748 39172 34750
rect 27244 34242 27300 34254
rect 27244 34190 27246 34242
rect 27298 34190 27300 34242
rect 27244 33572 27300 34190
rect 35644 34242 35700 34254
rect 35644 34190 35646 34242
rect 35698 34190 35700 34242
rect 27244 33506 27300 33516
rect 34412 34018 34468 34030
rect 34412 33966 34414 34018
rect 34466 33966 34468 34018
rect 27132 33460 27188 33470
rect 27132 33366 27188 33404
rect 29596 33460 29652 33470
rect 28140 33236 28196 33246
rect 27020 33234 28196 33236
rect 27020 33182 28142 33234
rect 28194 33182 28196 33234
rect 27020 33180 28196 33182
rect 26348 30942 26350 30994
rect 26402 30942 26404 30994
rect 26348 30930 26404 30942
rect 26572 31892 26852 31948
rect 26908 32562 26964 32574
rect 26908 32510 26910 32562
rect 26962 32510 26964 32562
rect 25340 30882 25732 30884
rect 25340 30830 25342 30882
rect 25394 30830 25732 30882
rect 25340 30828 25732 30830
rect 23548 29650 23604 29662
rect 23548 29598 23550 29650
rect 23602 29598 23604 29650
rect 23548 29540 23604 29598
rect 23548 29474 23604 29484
rect 24332 29540 24388 29550
rect 24332 29446 24388 29484
rect 24108 29428 24164 29438
rect 24108 29334 24164 29372
rect 24668 29314 24724 30044
rect 24668 29262 24670 29314
rect 24722 29262 24724 29314
rect 22204 28690 22260 28700
rect 22316 29092 22372 29102
rect 22316 28754 22372 29036
rect 22316 28702 22318 28754
rect 22370 28702 22372 28754
rect 22316 28690 22372 28702
rect 24668 28756 24724 29262
rect 24668 28690 24724 28700
rect 24780 30324 24836 30334
rect 24332 28644 24388 28654
rect 24332 28550 24388 28588
rect 24780 28642 24836 30268
rect 24780 28590 24782 28642
rect 24834 28590 24836 28642
rect 24780 28578 24836 28590
rect 25116 29986 25172 29998
rect 25116 29934 25118 29986
rect 25170 29934 25172 29986
rect 23548 28532 23604 28542
rect 23548 28438 23604 28476
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18396 28018 18452 28028
rect 19740 27972 19796 27982
rect 19740 27878 19796 27916
rect 20188 27860 20244 27870
rect 20188 27766 20244 27804
rect 18396 27746 18452 27758
rect 18396 27694 18398 27746
rect 18450 27694 18452 27746
rect 18284 27186 18340 27198
rect 18284 27134 18286 27186
rect 18338 27134 18340 27186
rect 18284 26964 18340 27134
rect 18284 26898 18340 26908
rect 18396 26740 18452 27694
rect 21196 27746 21252 28364
rect 21196 27694 21198 27746
rect 21250 27694 21252 27746
rect 21196 27682 21252 27694
rect 25004 27972 25060 27982
rect 25116 27972 25172 29934
rect 25340 29316 25396 30828
rect 25788 30100 25844 30110
rect 25788 30006 25844 30044
rect 25340 28644 25396 29260
rect 26124 29986 26180 29998
rect 26124 29934 26126 29986
rect 26178 29934 26180 29986
rect 26124 29316 26180 29934
rect 26124 29250 26180 29260
rect 26236 29764 26292 29774
rect 26236 29314 26292 29708
rect 26236 29262 26238 29314
rect 26290 29262 26292 29314
rect 26236 29250 26292 29262
rect 25228 27972 25284 27982
rect 25116 27970 25284 27972
rect 25116 27918 25230 27970
rect 25282 27918 25284 27970
rect 25116 27916 25284 27918
rect 25004 27298 25060 27916
rect 25228 27906 25284 27916
rect 25004 27246 25006 27298
rect 25058 27246 25060 27298
rect 25004 27234 25060 27246
rect 21868 27074 21924 27086
rect 21868 27022 21870 27074
rect 21922 27022 21924 27074
rect 18396 26674 18452 26684
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 17500 26462 17502 26514
rect 17554 26462 17556 26514
rect 17276 26066 17332 26078
rect 17276 26014 17278 26066
rect 17330 26014 17332 26066
rect 17164 23940 17220 23950
rect 17276 23940 17332 26014
rect 17500 25618 17556 26462
rect 19404 26404 19460 26414
rect 19404 26310 19460 26348
rect 20188 26404 20244 26414
rect 20188 26310 20244 26348
rect 20412 26290 20468 26302
rect 20412 26238 20414 26290
rect 20466 26238 20468 26290
rect 18396 26180 18452 26190
rect 17612 26178 18452 26180
rect 17612 26126 18398 26178
rect 18450 26126 18452 26178
rect 17612 26124 18452 26126
rect 17612 26066 17668 26124
rect 18396 26114 18452 26124
rect 19628 26180 19684 26190
rect 17612 26014 17614 26066
rect 17666 26014 17668 26066
rect 17612 26002 17668 26014
rect 17500 25566 17502 25618
rect 17554 25566 17556 25618
rect 17388 24948 17444 24958
rect 17388 24834 17444 24892
rect 17388 24782 17390 24834
rect 17442 24782 17444 24834
rect 17388 24770 17444 24782
rect 17164 23938 17332 23940
rect 17164 23886 17166 23938
rect 17218 23886 17332 23938
rect 17164 23884 17332 23886
rect 17164 23874 17220 23884
rect 17052 23268 17108 23772
rect 17500 23492 17556 25566
rect 17612 24836 17668 24846
rect 17612 24722 17668 24780
rect 17612 24670 17614 24722
rect 17666 24670 17668 24722
rect 17612 24658 17668 24670
rect 18284 24836 18340 24846
rect 18284 24722 18340 24780
rect 18844 24836 18900 24846
rect 18844 24742 18900 24780
rect 18284 24670 18286 24722
rect 18338 24670 18340 24722
rect 18284 24658 18340 24670
rect 19628 24722 19684 26124
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24670 19630 24722
rect 19682 24670 19684 24722
rect 19628 24658 19684 24670
rect 20076 24724 20132 24734
rect 20076 24630 20132 24668
rect 18060 24610 18116 24622
rect 18060 24558 18062 24610
rect 18114 24558 18116 24610
rect 17500 23378 17556 23436
rect 17500 23326 17502 23378
rect 17554 23326 17556 23378
rect 17052 23212 17220 23268
rect 16716 22932 16772 22942
rect 16492 22148 16548 22158
rect 16492 22146 16660 22148
rect 16492 22094 16494 22146
rect 16546 22094 16660 22146
rect 16492 22092 16660 22094
rect 16492 22082 16548 22092
rect 16604 20242 16660 22092
rect 16604 20190 16606 20242
rect 16658 20190 16660 20242
rect 16604 20178 16660 20190
rect 16604 20020 16660 20030
rect 16716 20020 16772 22876
rect 16828 22484 16884 22494
rect 16828 21028 16884 22428
rect 16940 21364 16996 21374
rect 16940 21270 16996 21308
rect 17052 21028 17108 21038
rect 16828 21026 17108 21028
rect 16828 20974 17054 21026
rect 17106 20974 17108 21026
rect 16828 20972 17108 20974
rect 17052 20962 17108 20972
rect 16604 20018 16772 20020
rect 16604 19966 16606 20018
rect 16658 19966 16772 20018
rect 16604 19964 16772 19966
rect 17164 20020 17220 23212
rect 17500 21812 17556 23326
rect 17836 23492 17892 23502
rect 17836 23154 17892 23436
rect 18060 23268 18116 24558
rect 19180 24612 19236 24622
rect 20412 24612 20468 26238
rect 21084 26290 21140 26302
rect 21084 26238 21086 26290
rect 21138 26238 21140 26290
rect 21084 26180 21140 26238
rect 21084 26114 21140 26124
rect 21532 26290 21588 26302
rect 21532 26238 21534 26290
rect 21586 26238 21588 26290
rect 20524 25620 20580 25630
rect 20524 25526 20580 25564
rect 19180 24610 19460 24612
rect 19180 24558 19182 24610
rect 19234 24558 19460 24610
rect 19180 24556 19460 24558
rect 19180 24546 19236 24556
rect 19404 23826 19460 24556
rect 20412 24050 20468 24556
rect 20412 23998 20414 24050
rect 20466 23998 20468 24050
rect 20412 23986 20468 23998
rect 21532 24052 21588 26238
rect 21868 25508 21924 27022
rect 21980 26852 22036 26862
rect 21980 26850 22372 26852
rect 21980 26798 21982 26850
rect 22034 26798 22372 26850
rect 21980 26796 22372 26798
rect 21980 26786 22036 26796
rect 22204 25508 22260 25518
rect 21868 25506 22260 25508
rect 21868 25454 22206 25506
rect 22258 25454 22260 25506
rect 21868 25452 22260 25454
rect 21532 23986 21588 23996
rect 22204 25284 22260 25452
rect 19404 23774 19406 23826
rect 19458 23774 19460 23826
rect 19404 23762 19460 23774
rect 20748 23826 20804 23838
rect 20748 23774 20750 23826
rect 20802 23774 20804 23826
rect 18060 23202 18116 23212
rect 19180 23716 19236 23726
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17836 23090 17892 23102
rect 18284 23154 18340 23166
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 17388 21810 17556 21812
rect 17388 21758 17502 21810
rect 17554 21758 17556 21810
rect 17388 21756 17556 21758
rect 17388 20914 17444 21756
rect 17500 21746 17556 21756
rect 17388 20862 17390 20914
rect 17442 20862 17444 20914
rect 17388 20244 17444 20862
rect 17948 21364 18004 21374
rect 17948 20690 18004 21308
rect 18284 20916 18340 23102
rect 18732 22372 18788 22382
rect 18732 22278 18788 22316
rect 19180 22372 19236 23660
rect 20188 23716 20244 23726
rect 20188 23714 20356 23716
rect 20188 23662 20190 23714
rect 20242 23662 20356 23714
rect 20188 23660 20356 23662
rect 20188 23650 20244 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19180 22370 19684 22372
rect 19180 22318 19182 22370
rect 19234 22318 19684 22370
rect 19180 22316 19684 22318
rect 19180 22306 19236 22316
rect 18732 21476 18788 21486
rect 18732 21382 18788 21420
rect 18284 20850 18340 20860
rect 19068 20916 19124 20926
rect 19628 20916 19684 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20300 21924 20356 23660
rect 20748 23378 20804 23774
rect 21420 23716 21476 23726
rect 21420 23622 21476 23660
rect 20748 23326 20750 23378
rect 20802 23326 20804 23378
rect 20748 23314 20804 23326
rect 21420 23380 21476 23390
rect 21420 23286 21476 23324
rect 20972 23268 21028 23278
rect 19836 21914 20100 21924
rect 20188 21868 20356 21924
rect 20412 22372 20468 22382
rect 20188 21812 20244 21868
rect 20076 21756 20244 21812
rect 20076 21698 20132 21756
rect 20076 21646 20078 21698
rect 20130 21646 20132 21698
rect 20076 21634 20132 21646
rect 19740 20916 19796 20926
rect 19628 20914 19796 20916
rect 19628 20862 19742 20914
rect 19794 20862 19796 20914
rect 19628 20860 19796 20862
rect 19068 20822 19124 20860
rect 19740 20850 19796 20860
rect 17948 20638 17950 20690
rect 18002 20638 18004 20690
rect 17948 20626 18004 20638
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 17388 20132 17668 20188
rect 17388 20020 17444 20030
rect 17164 20018 17444 20020
rect 17164 19966 17390 20018
rect 17442 19966 17444 20018
rect 17164 19964 17444 19966
rect 16604 19954 16660 19964
rect 17164 19908 17220 19964
rect 17388 19954 17444 19964
rect 17164 19842 17220 19852
rect 16380 18958 16382 19010
rect 16434 18958 16436 19010
rect 16380 18946 16436 18958
rect 17052 19010 17108 19022
rect 17052 18958 17054 19010
rect 17106 18958 17108 19010
rect 15596 18452 15652 18462
rect 15596 18358 15652 18396
rect 16268 18450 16324 18462
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 16268 18340 16324 18398
rect 16604 18340 16660 18350
rect 16268 18338 16660 18340
rect 16268 18286 16606 18338
rect 16658 18286 16660 18338
rect 16268 18284 16660 18286
rect 15484 16882 15540 16894
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16772 15540 16830
rect 16604 16884 16660 18284
rect 16604 16818 16660 16828
rect 16828 17778 16884 17790
rect 16828 17726 16830 17778
rect 16882 17726 16884 17778
rect 15932 16772 15988 16782
rect 15484 16770 15988 16772
rect 15484 16718 15934 16770
rect 15986 16718 15988 16770
rect 15484 16716 15988 16718
rect 15932 16100 15988 16716
rect 16156 16100 16212 16110
rect 15932 16098 16212 16100
rect 15932 16046 16158 16098
rect 16210 16046 16212 16098
rect 15932 16044 16212 16046
rect 16156 15876 16212 16044
rect 16156 15810 16212 15820
rect 15596 15316 15652 15326
rect 15148 15314 15652 15316
rect 15148 15262 15150 15314
rect 15202 15262 15598 15314
rect 15650 15262 15652 15314
rect 15148 15260 15652 15262
rect 15148 15250 15204 15260
rect 15596 15250 15652 15260
rect 16716 15316 16772 15326
rect 16828 15316 16884 17726
rect 17052 17220 17108 18958
rect 17164 19012 17220 19022
rect 17164 18918 17220 18956
rect 17612 18450 17668 20132
rect 20076 19906 20132 19918
rect 20076 19854 20078 19906
rect 20130 19854 20132 19906
rect 19068 19796 19124 19806
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 17836 19010 17892 19022
rect 17836 18958 17838 19010
rect 17890 18958 17892 19010
rect 17836 18452 17892 18958
rect 17836 18386 17892 18396
rect 18508 18452 18564 18462
rect 18508 18358 18564 18396
rect 19068 18450 19124 19740
rect 20076 19796 20132 19854
rect 20076 19730 20132 19740
rect 20412 19796 20468 22316
rect 20636 22146 20692 22158
rect 20636 22094 20638 22146
rect 20690 22094 20692 22146
rect 20636 21140 20692 22094
rect 20972 21810 21028 23212
rect 21644 22372 21700 22382
rect 21644 22278 21700 22316
rect 22204 22372 22260 25228
rect 22316 24946 22372 26796
rect 22428 26404 22484 26414
rect 22428 25730 22484 26348
rect 23772 26404 23828 26414
rect 23772 26310 23828 26348
rect 22428 25678 22430 25730
rect 22482 25678 22484 25730
rect 22428 25666 22484 25678
rect 23436 26180 23492 26190
rect 22316 24894 22318 24946
rect 22370 24894 22372 24946
rect 22316 24882 22372 24894
rect 22988 25508 23044 25518
rect 22316 24052 22372 24062
rect 22316 23958 22372 23996
rect 22316 23268 22372 23278
rect 22316 23174 22372 23212
rect 22204 22306 22260 22316
rect 22876 22372 22932 22382
rect 22988 22372 23044 25452
rect 23324 25506 23380 25518
rect 23324 25454 23326 25506
rect 23378 25454 23380 25506
rect 23100 24498 23156 24510
rect 23100 24446 23102 24498
rect 23154 24446 23156 24498
rect 23100 23828 23156 24446
rect 23324 24052 23380 25454
rect 23436 25508 23492 26124
rect 25340 26180 25396 28588
rect 25564 28644 25620 28654
rect 25564 27970 25620 28588
rect 25564 27918 25566 27970
rect 25618 27918 25620 27970
rect 25564 27906 25620 27918
rect 26348 27858 26404 27870
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26124 27748 26180 27758
rect 26348 27748 26404 27806
rect 26124 27746 26404 27748
rect 26124 27694 26126 27746
rect 26178 27694 26404 27746
rect 26124 27692 26404 27694
rect 26124 26964 26180 27692
rect 26572 27636 26628 31892
rect 26908 31556 26964 32510
rect 27020 32002 27076 33180
rect 28140 33170 28196 33180
rect 29372 33124 29428 33134
rect 29372 33122 29540 33124
rect 29372 33070 29374 33122
rect 29426 33070 29540 33122
rect 29372 33068 29540 33070
rect 29372 33058 29428 33068
rect 27468 33012 27524 33022
rect 27468 32562 27524 32956
rect 27468 32510 27470 32562
rect 27522 32510 27524 32562
rect 27468 32498 27524 32510
rect 29372 32900 29428 32910
rect 27020 31950 27022 32002
rect 27074 31950 27076 32002
rect 27020 31938 27076 31950
rect 29036 32004 29092 32014
rect 28588 31780 28644 31790
rect 28588 31686 28644 31724
rect 29036 31778 29092 31948
rect 29036 31726 29038 31778
rect 29090 31726 29092 31778
rect 27356 31556 27412 31566
rect 26908 31500 27356 31556
rect 27020 30324 27076 30334
rect 27020 30230 27076 30268
rect 27244 29538 27300 29550
rect 27244 29486 27246 29538
rect 27298 29486 27300 29538
rect 27244 29428 27300 29486
rect 27244 29362 27300 29372
rect 27356 29316 27412 31500
rect 28476 31554 28532 31566
rect 28476 31502 28478 31554
rect 28530 31502 28532 31554
rect 28476 31220 28532 31502
rect 29036 31556 29092 31726
rect 29036 31490 29092 31500
rect 28588 31220 28644 31230
rect 28476 31218 28644 31220
rect 28476 31166 28590 31218
rect 28642 31166 28644 31218
rect 28476 31164 28644 31166
rect 28588 31154 28644 31164
rect 29372 31218 29428 32844
rect 29372 31166 29374 31218
rect 29426 31166 29428 31218
rect 29372 31154 29428 31166
rect 29484 32564 29540 33068
rect 29484 31780 29540 32508
rect 29484 30884 29540 31724
rect 29596 31778 29652 33404
rect 30156 33458 30212 33470
rect 30156 33406 30158 33458
rect 30210 33406 30212 33458
rect 29820 33122 29876 33134
rect 29820 33070 29822 33122
rect 29874 33070 29876 33122
rect 29820 32788 29876 33070
rect 30156 33012 30212 33406
rect 32956 33460 33012 33470
rect 32956 33366 33012 33404
rect 30156 32946 30212 32956
rect 30492 33236 30548 33246
rect 30156 32788 30212 32798
rect 29820 32732 30156 32788
rect 29708 32674 29764 32686
rect 29708 32622 29710 32674
rect 29762 32622 29764 32674
rect 29708 31948 29764 32622
rect 30156 32004 30212 32732
rect 30492 32786 30548 33180
rect 31164 33234 31220 33246
rect 31164 33182 31166 33234
rect 31218 33182 31220 33234
rect 31164 32900 31220 33182
rect 33964 33236 34020 33246
rect 33964 33142 34020 33180
rect 31164 32834 31220 32844
rect 32732 33122 32788 33134
rect 32732 33070 32734 33122
rect 32786 33070 32788 33122
rect 30492 32734 30494 32786
rect 30546 32734 30548 32786
rect 30492 32722 30548 32734
rect 32396 32788 32452 32798
rect 32396 32694 32452 32732
rect 31164 32564 31220 32574
rect 31164 32470 31220 32508
rect 31948 32564 32004 32574
rect 31948 32470 32004 32508
rect 32732 32564 32788 33070
rect 32732 32498 32788 32508
rect 32956 33124 33012 33134
rect 29708 31892 29876 31948
rect 29596 31726 29598 31778
rect 29650 31726 29652 31778
rect 29596 31714 29652 31726
rect 29708 30884 29764 30894
rect 29484 30882 29764 30884
rect 29484 30830 29710 30882
rect 29762 30830 29764 30882
rect 29484 30828 29764 30830
rect 29596 30210 29652 30828
rect 29708 30818 29764 30828
rect 29820 30434 29876 31892
rect 30156 31218 30212 31948
rect 31388 32338 31444 32350
rect 31388 32286 31390 32338
rect 31442 32286 31444 32338
rect 31388 31556 31444 32286
rect 31388 31490 31444 31500
rect 31836 32340 31892 32350
rect 30156 31166 30158 31218
rect 30210 31166 30212 31218
rect 30156 31154 30212 31166
rect 30268 31220 30324 31230
rect 29820 30382 29822 30434
rect 29874 30382 29876 30434
rect 29820 30370 29876 30382
rect 29596 30158 29598 30210
rect 29650 30158 29652 30210
rect 28028 30100 28084 30110
rect 28028 30006 28084 30044
rect 29596 29652 29652 30158
rect 30268 30210 30324 31164
rect 31836 31106 31892 32284
rect 31948 31556 32004 31566
rect 31948 31462 32004 31500
rect 32732 31554 32788 31566
rect 32732 31502 32734 31554
rect 32786 31502 32788 31554
rect 31836 31054 31838 31106
rect 31890 31054 31892 31106
rect 31836 31042 31892 31054
rect 30604 30884 30660 30894
rect 30604 30790 30660 30828
rect 30268 30158 30270 30210
rect 30322 30158 30324 30210
rect 30268 30146 30324 30158
rect 31724 30100 31780 30110
rect 31052 29988 31108 29998
rect 31052 29894 31108 29932
rect 27356 29250 27412 29260
rect 28140 29316 28196 29326
rect 28140 29222 28196 29260
rect 29036 29314 29092 29326
rect 29036 29262 29038 29314
rect 29090 29262 29092 29314
rect 28252 28756 28308 28766
rect 28028 28644 28084 28654
rect 28028 28550 28084 28588
rect 27244 28418 27300 28430
rect 27244 28366 27246 28418
rect 27298 28366 27300 28418
rect 27244 28196 27300 28366
rect 27804 28420 27860 28430
rect 27804 28326 27860 28364
rect 28140 28418 28196 28430
rect 28140 28366 28142 28418
rect 28194 28366 28196 28418
rect 28140 28196 28196 28366
rect 27244 28140 28196 28196
rect 26124 26898 26180 26908
rect 26348 27580 26628 27636
rect 25788 26850 25844 26862
rect 25788 26798 25790 26850
rect 25842 26798 25844 26850
rect 25788 26516 25844 26798
rect 25900 26516 25956 26526
rect 25788 26514 25956 26516
rect 25788 26462 25902 26514
rect 25954 26462 25956 26514
rect 25788 26460 25956 26462
rect 25900 26450 25956 26460
rect 25788 26292 25844 26302
rect 25340 26086 25396 26124
rect 25676 26290 25844 26292
rect 25676 26238 25790 26290
rect 25842 26238 25844 26290
rect 25676 26236 25844 26238
rect 23436 24946 23492 25452
rect 23436 24894 23438 24946
rect 23490 24894 23492 24946
rect 23436 24882 23492 24894
rect 24556 26066 24612 26078
rect 24556 26014 24558 26066
rect 24610 26014 24612 26066
rect 23436 24052 23492 24062
rect 23324 23996 23436 24052
rect 23436 23986 23492 23996
rect 23324 23828 23380 23838
rect 23100 23826 23380 23828
rect 23100 23774 23326 23826
rect 23378 23774 23380 23826
rect 23100 23772 23380 23774
rect 23324 23762 23380 23772
rect 24556 23828 24612 26014
rect 24556 23762 24612 23772
rect 24892 25620 24948 25630
rect 23436 23044 23492 23054
rect 22876 22370 23044 22372
rect 22876 22318 22878 22370
rect 22930 22318 23044 22370
rect 22876 22316 23044 22318
rect 23324 23042 23492 23044
rect 23324 22990 23438 23042
rect 23490 22990 23492 23042
rect 23324 22988 23492 22990
rect 23324 22370 23380 22988
rect 23436 22978 23492 22988
rect 23324 22318 23326 22370
rect 23378 22318 23380 22370
rect 22876 22306 22932 22316
rect 23324 22306 23380 22318
rect 20972 21758 20974 21810
rect 21026 21758 21028 21810
rect 20972 21746 21028 21758
rect 21756 22146 21812 22158
rect 21756 22094 21758 22146
rect 21810 22094 21812 22146
rect 21756 21810 21812 22094
rect 21756 21758 21758 21810
rect 21810 21758 21812 21810
rect 21756 21746 21812 21758
rect 20636 21074 20692 21084
rect 23996 21586 24052 21598
rect 23996 21534 23998 21586
rect 24050 21534 24052 21586
rect 23884 20916 23940 20926
rect 20860 20804 20916 20814
rect 21420 20804 21476 20814
rect 20916 20802 21476 20804
rect 20916 20750 21422 20802
rect 21474 20750 21476 20802
rect 20916 20748 21476 20750
rect 20860 20710 20916 20748
rect 21420 20738 21476 20748
rect 20412 19730 20468 19740
rect 21196 20580 21252 20590
rect 20300 19234 20356 19246
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 19516 19012 19572 19022
rect 19516 18562 19572 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18498 19572 18510
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18386 19124 18398
rect 17052 17154 17108 17164
rect 17948 18338 18004 18350
rect 17948 18286 17950 18338
rect 18002 18286 18004 18338
rect 17948 16884 18004 18286
rect 20300 18340 20356 19182
rect 20300 18274 20356 18284
rect 20748 19236 20804 19246
rect 20748 18338 20804 19180
rect 20748 18286 20750 18338
rect 20802 18286 20804 18338
rect 20748 18274 20804 18286
rect 20860 19234 20916 19246
rect 20860 19182 20862 19234
rect 20914 19182 20916 19234
rect 20748 18116 20804 18126
rect 20076 17780 20132 17790
rect 20076 17666 20132 17724
rect 20748 17780 20804 18060
rect 20748 17686 20804 17724
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 17602 20132 17614
rect 19836 17276 20100 17286
rect 19180 17220 19236 17230
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19236 17164 19348 17220
rect 19836 17210 20100 17220
rect 19180 17154 19236 17164
rect 17948 16818 18004 16828
rect 18396 16884 18452 16894
rect 18396 16212 18452 16828
rect 18956 16884 19012 16894
rect 18956 16790 19012 16828
rect 16716 15314 16884 15316
rect 16716 15262 16718 15314
rect 16770 15262 16884 15314
rect 16716 15260 16884 15262
rect 16716 15250 16772 15260
rect 16716 15092 16772 15102
rect 16716 14998 16772 15036
rect 13692 14914 13748 14924
rect 15820 14644 15876 14654
rect 15820 14530 15876 14588
rect 15820 14478 15822 14530
rect 15874 14478 15876 14530
rect 15820 14466 15876 14478
rect 16268 14530 16324 14542
rect 16828 14532 16884 15260
rect 18284 16210 18452 16212
rect 18284 16158 18398 16210
rect 18450 16158 18452 16210
rect 18284 16156 18452 16158
rect 16268 14478 16270 14530
rect 16322 14478 16324 14530
rect 13244 13916 13524 13972
rect 10668 13858 10724 13870
rect 10668 13806 10670 13858
rect 10722 13806 10724 13858
rect 10668 13188 10724 13806
rect 13356 13746 13412 13758
rect 13356 13694 13358 13746
rect 13410 13694 13412 13746
rect 12012 13634 12068 13646
rect 12012 13582 12014 13634
rect 12066 13582 12068 13634
rect 12012 13188 12068 13582
rect 12012 13132 12404 13188
rect 10668 13122 10724 13132
rect 10668 12964 10724 12974
rect 10444 12962 10724 12964
rect 10444 12910 10670 12962
rect 10722 12910 10724 12962
rect 10444 12908 10724 12910
rect 10668 12740 10724 12908
rect 11788 12964 11844 12974
rect 10668 12674 10724 12684
rect 11228 12740 11284 12750
rect 11228 12646 11284 12684
rect 9884 12086 9940 12124
rect 10108 12404 10164 12414
rect 10108 11282 10164 12348
rect 10108 11230 10110 11282
rect 10162 11230 10164 11282
rect 10108 11218 10164 11230
rect 10444 12180 10500 12190
rect 9660 10498 9828 10500
rect 9660 10446 9662 10498
rect 9714 10446 9828 10498
rect 9660 10444 9828 10446
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2940 9828 2996 9838
rect 8204 9828 8260 9838
rect 2940 9826 3332 9828
rect 2940 9774 2942 9826
rect 2994 9774 3332 9826
rect 2940 9772 3332 9774
rect 2940 9762 2996 9772
rect 2044 9716 2100 9726
rect 2044 9622 2100 9660
rect 2940 9042 2996 9054
rect 2940 8990 2942 9042
rect 2994 8990 2996 9042
rect 1932 8932 1988 8942
rect 1932 8838 1988 8876
rect 2940 8428 2996 8990
rect 3276 8428 3332 9772
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2940 8372 3220 8428
rect 3276 8372 3668 8428
rect 2716 8258 2772 8270
rect 2716 8206 2718 8258
rect 2770 8206 2772 8258
rect 2044 8148 2100 8158
rect 2044 8054 2100 8092
rect 1932 7362 1988 7374
rect 1932 7310 1934 7362
rect 1986 7310 1988 7362
rect 1932 6804 1988 7310
rect 1932 6738 1988 6748
rect 2044 6578 2100 6590
rect 2044 6526 2046 6578
rect 2098 6526 2100 6578
rect 2044 6132 2100 6526
rect 2716 6580 2772 8206
rect 2940 7474 2996 7486
rect 2940 7422 2942 7474
rect 2994 7422 2996 7474
rect 2716 6514 2772 6524
rect 2828 6690 2884 6702
rect 2828 6638 2830 6690
rect 2882 6638 2884 6690
rect 2044 6066 2100 6076
rect 2716 5908 2772 5918
rect 2604 5906 2772 5908
rect 2604 5854 2718 5906
rect 2770 5854 2772 5906
rect 2604 5852 2772 5854
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5460 1988 5742
rect 1932 5394 1988 5404
rect 2044 5124 2100 5134
rect 1708 4900 1764 4910
rect 1708 4898 1876 4900
rect 1708 4846 1710 4898
rect 1762 4846 1876 4898
rect 1708 4844 1876 4846
rect 1708 4834 1764 4844
rect 1708 4452 1764 4490
rect 1708 4386 1764 4396
rect 1708 4228 1764 4238
rect 1708 3556 1764 4172
rect 1708 3462 1764 3500
rect 1820 1764 1876 4844
rect 2044 4562 2100 5068
rect 2268 5012 2324 5022
rect 2044 4510 2046 4562
rect 2098 4510 2100 4562
rect 2044 4498 2100 4510
rect 2156 5010 2324 5012
rect 2156 4958 2270 5010
rect 2322 4958 2324 5010
rect 2156 4956 2324 4958
rect 2044 3444 2100 3454
rect 2156 3444 2212 4956
rect 2268 4946 2324 4956
rect 2604 5010 2660 5852
rect 2716 5842 2772 5852
rect 2604 4958 2606 5010
rect 2658 4958 2660 5010
rect 2604 4946 2660 4958
rect 2716 5236 2772 5246
rect 2380 4450 2436 4462
rect 2380 4398 2382 4450
rect 2434 4398 2436 4450
rect 2380 4116 2436 4398
rect 2380 4050 2436 4060
rect 2044 3442 2212 3444
rect 2044 3390 2046 3442
rect 2098 3390 2212 3442
rect 2044 3388 2212 3390
rect 2380 3556 2436 3566
rect 2380 3442 2436 3500
rect 2380 3390 2382 3442
rect 2434 3390 2436 3442
rect 2044 3378 2100 3388
rect 1820 1698 1876 1708
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2380 756 2436 3390
rect 2716 3442 2772 5180
rect 2828 4564 2884 6638
rect 2940 5010 2996 7422
rect 3164 6132 3220 8372
rect 3276 8034 3332 8046
rect 3276 7982 3278 8034
rect 3330 7982 3332 8034
rect 3276 7476 3332 7982
rect 3276 7410 3332 7420
rect 3276 6132 3332 6142
rect 3164 6130 3332 6132
rect 3164 6078 3278 6130
rect 3330 6078 3332 6130
rect 3164 6076 3332 6078
rect 3276 6066 3332 6076
rect 3500 5908 3556 5918
rect 3388 5906 3556 5908
rect 3388 5854 3502 5906
rect 3554 5854 3556 5906
rect 3388 5852 3556 5854
rect 2940 4958 2942 5010
rect 2994 4958 2996 5010
rect 2940 4946 2996 4958
rect 3276 5012 3332 5022
rect 3276 4918 3332 4956
rect 2940 4564 2996 4574
rect 2828 4562 2996 4564
rect 2828 4510 2942 4562
rect 2994 4510 2996 4562
rect 2828 4508 2996 4510
rect 2940 4498 2996 4508
rect 3276 4564 3332 4574
rect 3276 4450 3332 4508
rect 3276 4398 3278 4450
rect 3330 4398 3332 4450
rect 3276 4386 3332 4398
rect 3052 3444 3108 3454
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3378 2772 3390
rect 2940 3388 3052 3444
rect 2380 690 2436 700
rect 2688 0 2800 800
rect 2940 84 2996 3388
rect 3052 3350 3108 3388
rect 3388 3442 3444 5852
rect 3500 5842 3556 5852
rect 3612 5010 3668 8372
rect 8204 8258 8260 9772
rect 9548 9828 9604 9838
rect 9660 9828 9716 10444
rect 9604 9772 9716 9828
rect 9996 9826 10052 9838
rect 9996 9774 9998 9826
rect 10050 9774 10052 9826
rect 8204 8206 8206 8258
rect 8258 8206 8260 8258
rect 8204 8194 8260 8206
rect 8652 9492 8708 9502
rect 8652 8258 8708 9436
rect 9548 8932 9604 9772
rect 9996 9380 10052 9774
rect 9996 9314 10052 9324
rect 10444 9042 10500 12124
rect 11788 12180 11844 12908
rect 12236 12738 12292 12750
rect 12236 12686 12238 12738
rect 12290 12686 12292 12738
rect 12236 12404 12292 12686
rect 12236 12338 12292 12348
rect 11788 12086 11844 12124
rect 12236 12178 12292 12190
rect 12236 12126 12238 12178
rect 12290 12126 12292 12178
rect 12236 12068 12292 12126
rect 12348 12180 12404 13132
rect 12460 12964 12516 12974
rect 12460 12870 12516 12908
rect 12572 12180 12628 12190
rect 12348 12178 12628 12180
rect 12348 12126 12574 12178
rect 12626 12126 12628 12178
rect 12348 12124 12628 12126
rect 12572 12114 12628 12124
rect 12236 12012 12516 12068
rect 11676 11954 11732 11966
rect 11676 11902 11678 11954
rect 11730 11902 11732 11954
rect 11676 10836 11732 11902
rect 12348 11394 12404 11406
rect 12348 11342 12350 11394
rect 12402 11342 12404 11394
rect 11676 10780 12292 10836
rect 11564 10724 11620 10734
rect 11564 10630 11620 10668
rect 10556 10498 10612 10510
rect 10556 10446 10558 10498
rect 10610 10446 10612 10498
rect 10556 9492 10612 10446
rect 12236 9714 12292 10780
rect 12348 10052 12404 11342
rect 12460 11396 12516 12012
rect 13020 11396 13076 11406
rect 13356 11396 13412 13694
rect 13468 12964 13524 13916
rect 13916 13746 13972 13758
rect 13916 13694 13918 13746
rect 13970 13694 13972 13746
rect 13580 12964 13636 12974
rect 13524 12962 13860 12964
rect 13524 12910 13582 12962
rect 13634 12910 13860 12962
rect 13524 12908 13860 12910
rect 13468 12870 13524 12908
rect 13580 12898 13636 12908
rect 12460 11394 13412 11396
rect 12460 11342 13022 11394
rect 13074 11342 13412 11394
rect 12460 11340 13412 11342
rect 12684 10610 12740 11340
rect 13020 11330 13076 11340
rect 13356 11172 13412 11340
rect 13580 11172 13636 11182
rect 13356 11116 13580 11172
rect 13580 11078 13636 11116
rect 12684 10558 12686 10610
rect 12738 10558 12740 10610
rect 12684 10546 12740 10558
rect 13132 10612 13188 10622
rect 13132 10610 13300 10612
rect 13132 10558 13134 10610
rect 13186 10558 13300 10610
rect 13132 10556 13300 10558
rect 13132 10546 13188 10556
rect 12460 10052 12516 10062
rect 12348 9996 12460 10052
rect 12460 9986 12516 9996
rect 12236 9662 12238 9714
rect 12290 9662 12292 9714
rect 12236 9650 12292 9662
rect 13020 9604 13076 9614
rect 13020 9602 13188 9604
rect 13020 9550 13022 9602
rect 13074 9550 13188 9602
rect 13020 9548 13188 9550
rect 13020 9538 13076 9548
rect 10556 9426 10612 9436
rect 12012 9380 12068 9390
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 8978 10500 8990
rect 11676 9156 11732 9166
rect 9548 8866 9604 8876
rect 10332 8818 10388 8830
rect 10332 8766 10334 8818
rect 10386 8766 10388 8818
rect 10332 8428 10388 8766
rect 10332 8372 10948 8428
rect 8652 8206 8654 8258
rect 8706 8206 8708 8258
rect 8652 8194 8708 8206
rect 10892 8146 10948 8372
rect 11676 8370 11732 9100
rect 12012 8930 12068 9324
rect 13020 9156 13076 9166
rect 13020 9062 13076 9100
rect 12012 8878 12014 8930
rect 12066 8878 12068 8930
rect 12012 8866 12068 8878
rect 12124 8932 12180 8942
rect 11676 8318 11678 8370
rect 11730 8318 11732 8370
rect 11676 8306 11732 8318
rect 12124 8370 12180 8876
rect 12124 8318 12126 8370
rect 12178 8318 12180 8370
rect 12124 8306 12180 8318
rect 10892 8094 10894 8146
rect 10946 8094 10948 8146
rect 10892 8082 10948 8094
rect 13132 7588 13188 9548
rect 13132 7522 13188 7532
rect 13244 7362 13300 10556
rect 13804 9826 13860 12908
rect 13916 11508 13972 13694
rect 16268 13076 16324 14478
rect 16716 14476 16828 14532
rect 16380 13972 16436 13982
rect 16380 13970 16660 13972
rect 16380 13918 16382 13970
rect 16434 13918 16660 13970
rect 16380 13916 16660 13918
rect 16380 13906 16436 13916
rect 16492 13076 16548 13086
rect 16268 13074 16548 13076
rect 16268 13022 16494 13074
rect 16546 13022 16548 13074
rect 16268 13020 16548 13022
rect 16492 13010 16548 13020
rect 14140 12740 14196 12750
rect 14140 12738 14980 12740
rect 14140 12686 14142 12738
rect 14194 12686 14980 12738
rect 14140 12684 14980 12686
rect 14140 12674 14196 12684
rect 14924 12402 14980 12684
rect 14924 12350 14926 12402
rect 14978 12350 14980 12402
rect 14924 12338 14980 12350
rect 16156 12738 16212 12750
rect 16156 12686 16158 12738
rect 16210 12686 16212 12738
rect 15708 11956 15764 11966
rect 15708 11954 15988 11956
rect 15708 11902 15710 11954
rect 15762 11902 15988 11954
rect 15708 11900 15988 11902
rect 15708 11890 15764 11900
rect 14924 11508 14980 11518
rect 13916 11506 14980 11508
rect 13916 11454 14926 11506
rect 14978 11454 14980 11506
rect 13916 11452 14980 11454
rect 14924 11442 14980 11452
rect 15932 11282 15988 11900
rect 16156 11396 16212 12686
rect 16604 12180 16660 13916
rect 16604 12114 16660 12124
rect 16716 12178 16772 14476
rect 16828 14466 16884 14476
rect 17500 14644 17556 14654
rect 17500 13748 17556 14588
rect 18284 14644 18340 16156
rect 18396 16146 18452 16156
rect 19292 15428 19348 17164
rect 19404 16884 19460 16894
rect 19740 16884 19796 16894
rect 19404 16790 19460 16828
rect 19516 16882 19796 16884
rect 19516 16830 19742 16882
rect 19794 16830 19796 16882
rect 19516 16828 19796 16830
rect 19404 15428 19460 15438
rect 19292 15426 19460 15428
rect 19292 15374 19406 15426
rect 19458 15374 19460 15426
rect 19292 15372 19460 15374
rect 19404 15362 19460 15372
rect 18396 15202 18452 15214
rect 18396 15150 18398 15202
rect 18450 15150 18452 15202
rect 18396 14980 18452 15150
rect 18396 14914 18452 14924
rect 18508 15092 18564 15102
rect 18284 14578 18340 14588
rect 18508 14418 18564 15036
rect 18508 14366 18510 14418
rect 18562 14366 18564 14418
rect 18508 14354 18564 14366
rect 19292 14308 19348 14318
rect 19292 14306 19460 14308
rect 19292 14254 19294 14306
rect 19346 14254 19460 14306
rect 19292 14252 19460 14254
rect 19292 14242 19348 14252
rect 17500 13746 17668 13748
rect 17500 13694 17502 13746
rect 17554 13694 17668 13746
rect 17500 13692 17668 13694
rect 17500 13682 17556 13692
rect 16940 13524 16996 13534
rect 16940 13522 17556 13524
rect 16940 13470 16942 13522
rect 16994 13470 17556 13522
rect 16940 13468 17556 13470
rect 16940 13458 16996 13468
rect 17500 12850 17556 13468
rect 17500 12798 17502 12850
rect 17554 12798 17556 12850
rect 17500 12786 17556 12798
rect 17500 12404 17556 12414
rect 17612 12404 17668 13692
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 12964 18004 13694
rect 17948 12898 18004 12908
rect 18732 12964 18788 12974
rect 17948 12404 18004 12414
rect 17500 12402 18004 12404
rect 17500 12350 17502 12402
rect 17554 12350 17950 12402
rect 18002 12350 18004 12402
rect 17500 12348 18004 12350
rect 17500 12338 17556 12348
rect 16716 12126 16718 12178
rect 16770 12126 16772 12178
rect 16716 12114 16772 12126
rect 17500 12180 17556 12190
rect 16716 11954 16772 11966
rect 16716 11902 16718 11954
rect 16770 11902 16772 11954
rect 16716 11620 16772 11902
rect 16716 11564 17220 11620
rect 16492 11396 16548 11406
rect 16156 11340 16492 11396
rect 15932 11230 15934 11282
rect 15986 11230 15988 11282
rect 15932 11218 15988 11230
rect 14588 11172 14644 11182
rect 14588 10836 14644 11116
rect 15036 10836 15092 10846
rect 14588 10780 15036 10836
rect 14364 10724 14420 10734
rect 14364 10050 14420 10668
rect 14364 9998 14366 10050
rect 14418 9998 14420 10050
rect 14364 9986 14420 9998
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13804 9762 13860 9774
rect 15036 9826 15092 10780
rect 16492 10836 16548 11340
rect 16604 11172 16660 11182
rect 16604 11078 16660 11116
rect 17164 11170 17220 11564
rect 17164 11118 17166 11170
rect 17218 11118 17220 11170
rect 17164 11106 17220 11118
rect 16492 10742 16548 10780
rect 17500 10834 17556 12124
rect 17948 11396 18004 12348
rect 18732 12066 18788 12908
rect 19404 12516 19460 14252
rect 19516 13074 19572 16828
rect 19740 16818 19796 16828
rect 20860 16884 20916 19182
rect 21196 19234 21252 20524
rect 23884 20188 23940 20860
rect 23772 20132 23940 20188
rect 21756 19908 21812 19918
rect 21196 19182 21198 19234
rect 21250 19182 21252 19234
rect 21196 19170 21252 19182
rect 21644 19906 21812 19908
rect 21644 19854 21758 19906
rect 21810 19854 21812 19906
rect 21644 19852 21812 19854
rect 21644 18228 21700 19852
rect 21756 19842 21812 19852
rect 21756 19236 21812 19246
rect 21756 19142 21812 19180
rect 23772 19012 23828 20132
rect 23996 19348 24052 21534
rect 24444 21588 24500 21598
rect 23996 19282 24052 19292
rect 24108 21140 24164 21150
rect 24108 19122 24164 21084
rect 24444 20580 24500 21532
rect 24892 20916 24948 25564
rect 25676 25284 25732 26236
rect 25788 26226 25844 26236
rect 25676 24722 25732 25228
rect 25900 25282 25956 25294
rect 25900 25230 25902 25282
rect 25954 25230 25956 25282
rect 25900 24946 25956 25230
rect 25900 24894 25902 24946
rect 25954 24894 25956 24946
rect 25900 24882 25956 24894
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 25676 24658 25732 24670
rect 25116 24052 25172 24062
rect 25116 23958 25172 23996
rect 26124 23828 26180 23838
rect 26124 23734 26180 23772
rect 26348 23380 26404 27580
rect 26460 27412 26516 27422
rect 26460 25730 26516 27356
rect 28140 27076 28196 27086
rect 28252 27076 28308 28700
rect 29036 28756 29092 29262
rect 29036 28690 29092 28700
rect 29036 28532 29092 28542
rect 29036 27298 29092 28476
rect 29036 27246 29038 27298
rect 29090 27246 29092 27298
rect 29036 27234 29092 27246
rect 29260 28418 29316 28430
rect 29260 28366 29262 28418
rect 29314 28366 29316 28418
rect 28140 27074 28308 27076
rect 28140 27022 28142 27074
rect 28194 27022 28308 27074
rect 28140 27020 28308 27022
rect 28700 27074 28756 27086
rect 28700 27022 28702 27074
rect 28754 27022 28756 27074
rect 28140 27010 28196 27020
rect 26908 26964 26964 26974
rect 26460 25678 26462 25730
rect 26514 25678 26516 25730
rect 26460 25666 26516 25678
rect 26796 26180 26852 26190
rect 26796 25620 26852 26124
rect 26572 25618 26852 25620
rect 26572 25566 26798 25618
rect 26850 25566 26852 25618
rect 26572 25564 26852 25566
rect 26348 23314 26404 23324
rect 26460 23380 26516 23390
rect 26572 23380 26628 25564
rect 26796 25554 26852 25564
rect 26460 23378 26628 23380
rect 26460 23326 26462 23378
rect 26514 23326 26628 23378
rect 26460 23324 26628 23326
rect 26908 23378 26964 26908
rect 27244 26292 27300 26302
rect 27244 25620 27300 26236
rect 28364 26292 28420 26302
rect 28364 26198 28420 26236
rect 27244 25526 27300 25564
rect 28700 25508 28756 27022
rect 28924 26180 28980 26190
rect 28924 26086 28980 26124
rect 29260 25508 29316 28366
rect 29596 28082 29652 29596
rect 31388 29652 31444 29662
rect 31724 29652 31780 30044
rect 31444 29596 31780 29652
rect 31388 29558 31444 29596
rect 29596 28030 29598 28082
rect 29650 28030 29652 28082
rect 29596 28018 29652 28030
rect 30268 29538 30324 29550
rect 30268 29486 30270 29538
rect 30322 29486 30324 29538
rect 30268 27412 30324 29486
rect 31724 29426 31780 29596
rect 31836 29988 31892 29998
rect 31836 29650 31892 29932
rect 31836 29598 31838 29650
rect 31890 29598 31892 29650
rect 31836 29586 31892 29598
rect 32732 29540 32788 31502
rect 32956 31218 33012 33068
rect 33292 33012 33348 33022
rect 32956 31166 32958 31218
rect 33010 31166 33012 31218
rect 32956 31154 33012 31166
rect 33068 31778 33124 31790
rect 33068 31726 33070 31778
rect 33122 31726 33124 31778
rect 32732 29474 32788 29484
rect 31724 29374 31726 29426
rect 31778 29374 31780 29426
rect 31724 29362 31780 29374
rect 33068 29316 33124 31726
rect 33292 31780 33348 32956
rect 34412 33012 34468 33966
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35644 33124 35700 34190
rect 37324 34242 37380 34254
rect 37324 34190 37326 34242
rect 37378 34190 37380 34242
rect 35644 33058 35700 33068
rect 36540 33124 36596 33134
rect 34412 32946 34468 32956
rect 35084 32786 35140 32798
rect 35084 32734 35086 32786
rect 35138 32734 35140 32786
rect 33516 32564 33572 32574
rect 33516 32470 33572 32508
rect 33404 32450 33460 32462
rect 33404 32398 33406 32450
rect 33458 32398 33460 32450
rect 33404 31948 33460 32398
rect 34412 32340 34468 32350
rect 34412 32246 34468 32284
rect 33404 31892 33684 31948
rect 33404 31780 33460 31790
rect 33292 31778 33460 31780
rect 33292 31726 33406 31778
rect 33458 31726 33460 31778
rect 33292 31724 33460 31726
rect 33404 31714 33460 31724
rect 33628 31218 33684 31892
rect 35084 31892 35140 32734
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35084 31826 35140 31836
rect 36540 31890 36596 33068
rect 37212 33122 37268 33134
rect 37212 33070 37214 33122
rect 37266 33070 37268 33122
rect 37212 32452 37268 33070
rect 37324 33124 37380 34190
rect 37324 33058 37380 33068
rect 37548 34020 37604 34030
rect 37548 32562 37604 33964
rect 38444 34020 38500 34030
rect 38444 33926 38500 33964
rect 38444 33460 38500 33470
rect 37772 33458 38500 33460
rect 37772 33406 38446 33458
rect 38498 33406 38500 33458
rect 37772 33404 38500 33406
rect 37548 32510 37550 32562
rect 37602 32510 37604 32562
rect 37548 32498 37604 32510
rect 37660 33122 37716 33134
rect 37660 33070 37662 33122
rect 37714 33070 37716 33122
rect 37212 31948 37268 32396
rect 37436 32004 37492 32014
rect 37660 32004 37716 33070
rect 37492 31948 37716 32004
rect 36540 31838 36542 31890
rect 36594 31838 36596 31890
rect 36540 31826 36596 31838
rect 37100 31892 37156 31902
rect 37212 31892 37380 31948
rect 37100 31798 37156 31836
rect 37324 31778 37380 31892
rect 37324 31726 37326 31778
rect 37378 31726 37380 31778
rect 33628 31166 33630 31218
rect 33682 31166 33684 31218
rect 33628 31154 33684 31166
rect 35756 31554 35812 31566
rect 35756 31502 35758 31554
rect 35810 31502 35812 31554
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35756 30322 35812 31502
rect 36092 30994 36148 31006
rect 36092 30942 36094 30994
rect 36146 30942 36148 30994
rect 36092 30884 36148 30942
rect 36652 30994 36708 31006
rect 36652 30942 36654 30994
rect 36706 30942 36708 30994
rect 36652 30884 36708 30942
rect 36988 30884 37044 30894
rect 36652 30882 37044 30884
rect 36652 30830 36990 30882
rect 37042 30830 37044 30882
rect 36652 30828 37044 30830
rect 36092 30818 36148 30828
rect 36988 30770 37044 30828
rect 36988 30718 36990 30770
rect 37042 30718 37044 30770
rect 36876 30436 36932 30446
rect 35756 30270 35758 30322
rect 35810 30270 35812 30322
rect 35756 30258 35812 30270
rect 36764 30324 36820 30334
rect 33404 30210 33460 30222
rect 33404 30158 33406 30210
rect 33458 30158 33460 30210
rect 33404 29764 33460 30158
rect 33404 29698 33460 29708
rect 33964 30210 34020 30222
rect 33964 30158 33966 30210
rect 34018 30158 34020 30210
rect 33852 29652 33908 29662
rect 33852 29558 33908 29596
rect 33404 29316 33460 29326
rect 33516 29316 33572 29326
rect 33068 29314 33516 29316
rect 33068 29262 33406 29314
rect 33458 29262 33516 29314
rect 33068 29260 33516 29262
rect 33404 29250 33460 29260
rect 30268 27346 30324 27356
rect 30492 28754 30548 28766
rect 33292 28756 33348 28766
rect 30492 28702 30494 28754
rect 30546 28702 30548 28754
rect 28700 25506 29316 25508
rect 28700 25454 29262 25506
rect 29314 25454 29316 25506
rect 28700 25452 29316 25454
rect 28812 24612 28868 24622
rect 28812 24518 28868 24556
rect 26908 23326 26910 23378
rect 26962 23326 26964 23378
rect 26460 23314 26516 23324
rect 26908 23156 26964 23326
rect 27244 23156 27300 23166
rect 26908 23154 27300 23156
rect 26908 23102 27246 23154
rect 27298 23102 27300 23154
rect 26908 23100 27300 23102
rect 26908 22484 26964 23100
rect 27244 23090 27300 23100
rect 26796 22428 26964 22484
rect 26348 22260 26404 22270
rect 26348 22166 26404 22204
rect 25564 22146 25620 22158
rect 25564 22094 25566 22146
rect 25618 22094 25620 22146
rect 25116 21588 25172 21598
rect 25116 21494 25172 21532
rect 24892 20822 24948 20860
rect 24444 20514 24500 20524
rect 25564 20130 25620 22094
rect 25788 21588 25844 21598
rect 25788 21494 25844 21532
rect 25564 20078 25566 20130
rect 25618 20078 25620 20130
rect 25564 20066 25620 20078
rect 25676 20018 25732 20030
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25676 19796 25732 19966
rect 25676 19730 25732 19740
rect 26684 19906 26740 19918
rect 26684 19854 26686 19906
rect 26738 19854 26740 19906
rect 26124 19348 26180 19358
rect 26124 19254 26180 19292
rect 24108 19070 24110 19122
rect 24162 19070 24164 19122
rect 24108 19058 24164 19070
rect 24892 19124 24948 19134
rect 24892 19030 24948 19068
rect 23212 18340 23268 18350
rect 23212 18246 23268 18284
rect 21756 18228 21812 18238
rect 21644 18172 21756 18228
rect 21756 18162 21812 18172
rect 22876 18228 22932 18238
rect 22876 17778 22932 18172
rect 22876 17726 22878 17778
rect 22930 17726 22932 17778
rect 22876 17714 22932 17726
rect 22092 16996 22148 17006
rect 20860 16818 20916 16828
rect 21980 16994 22148 16996
rect 21980 16942 22094 16994
rect 22146 16942 22148 16994
rect 21980 16940 22148 16942
rect 21980 16322 22036 16940
rect 22092 16930 22148 16940
rect 23548 16772 23604 16782
rect 22876 16660 22932 16670
rect 22876 16566 22932 16604
rect 21980 16270 21982 16322
rect 22034 16270 22036 16322
rect 21980 16258 22036 16270
rect 22092 16098 22148 16110
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 20524 15876 20580 15886
rect 20524 15782 20580 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 21308 15426 21364 15438
rect 21308 15374 21310 15426
rect 21362 15374 21364 15426
rect 20524 15204 20580 15214
rect 20524 15110 20580 15148
rect 21308 14868 21364 15374
rect 21308 14802 21364 14812
rect 20748 14644 20804 14654
rect 21420 14644 21476 14654
rect 20748 14550 20804 14588
rect 21308 14588 21420 14644
rect 20300 14532 20356 14542
rect 20300 14438 20356 14476
rect 20188 14306 20244 14318
rect 20188 14254 20190 14306
rect 20242 14254 20244 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13970 20244 14254
rect 20188 13918 20190 13970
rect 20242 13918 20244 13970
rect 20188 13906 20244 13918
rect 21308 13746 21364 14588
rect 21420 14550 21476 14588
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 21308 13682 21364 13694
rect 21644 14532 21700 14542
rect 22092 14532 22148 16046
rect 23548 16098 23604 16716
rect 23548 16046 23550 16098
rect 23602 16046 23604 16098
rect 23548 16034 23604 16046
rect 23772 15876 23828 18956
rect 25788 19012 25844 19022
rect 24556 18564 24612 18574
rect 24556 18470 24612 18508
rect 25788 18452 25844 18956
rect 25788 18386 25844 18396
rect 26348 18452 26404 18462
rect 26684 18452 26740 19854
rect 26348 18450 26740 18452
rect 26348 18398 26350 18450
rect 26402 18398 26740 18450
rect 26348 18396 26740 18398
rect 24108 18228 24164 18238
rect 24108 17666 24164 18172
rect 24108 17614 24110 17666
rect 24162 17614 24164 17666
rect 24108 17602 24164 17614
rect 26236 18226 26292 18238
rect 26236 18174 26238 18226
rect 26290 18174 26292 18226
rect 25340 16884 25396 16894
rect 25340 16790 25396 16828
rect 25788 16882 25844 16894
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 24220 16772 24276 16782
rect 23772 15810 23828 15820
rect 23996 16098 24052 16110
rect 23996 16046 23998 16098
rect 24050 16046 24052 16098
rect 23996 15652 24052 16046
rect 23996 15586 24052 15596
rect 23660 15314 23716 15326
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 23548 15204 23604 15214
rect 22316 14868 22372 14878
rect 22316 14754 22372 14812
rect 22316 14702 22318 14754
rect 22370 14702 22372 14754
rect 22316 14690 22372 14702
rect 22204 14532 22260 14542
rect 22092 14476 22204 14532
rect 20972 13524 21028 13534
rect 19516 13022 19518 13074
rect 19570 13022 19572 13074
rect 19516 13010 19572 13022
rect 20636 13522 21028 13524
rect 20636 13470 20974 13522
rect 21026 13470 21028 13522
rect 20636 13468 21028 13470
rect 20636 12850 20692 13468
rect 20972 13458 21028 13468
rect 21644 12964 21700 14476
rect 22204 14438 22260 14476
rect 23212 13860 23268 13870
rect 21644 12870 21700 12908
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 20636 12798 20638 12850
rect 20690 12798 20692 12850
rect 20636 12786 20692 12798
rect 21532 12850 21588 12862
rect 21532 12798 21534 12850
rect 21586 12798 21588 12850
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19404 12460 19684 12516
rect 19836 12506 20100 12516
rect 19628 12292 19684 12460
rect 19740 12292 19796 12302
rect 19628 12290 19796 12292
rect 19628 12238 19742 12290
rect 19794 12238 19796 12290
rect 19628 12236 19796 12238
rect 19740 12226 19796 12236
rect 21196 12290 21252 12302
rect 21196 12238 21198 12290
rect 21250 12238 21252 12290
rect 18732 12014 18734 12066
rect 18786 12014 18788 12066
rect 18732 12002 18788 12014
rect 20412 11954 20468 11966
rect 20412 11902 20414 11954
rect 20466 11902 20468 11954
rect 17948 11330 18004 11340
rect 18620 11396 18676 11406
rect 17500 10782 17502 10834
rect 17554 10782 17556 10834
rect 17500 10770 17556 10782
rect 15372 10724 15428 10734
rect 15372 10630 15428 10668
rect 17724 10612 17780 10622
rect 18620 10612 18676 11340
rect 19628 11394 19684 11406
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19292 10612 19348 10622
rect 17780 10556 17892 10612
rect 17724 10518 17780 10556
rect 16156 10386 16212 10398
rect 16156 10334 16158 10386
rect 16210 10334 16212 10386
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 15036 9762 15092 9774
rect 15372 10052 15428 10062
rect 13916 8932 13972 8942
rect 13916 8838 13972 8876
rect 15372 8930 15428 9996
rect 15372 8878 15374 8930
rect 15426 8878 15428 8930
rect 15372 8866 15428 8878
rect 15484 9826 15540 9838
rect 15484 9774 15486 9826
rect 15538 9774 15540 9826
rect 15484 8428 15540 9774
rect 16156 9380 16212 10334
rect 17724 9602 17780 9614
rect 17724 9550 17726 9602
rect 17778 9550 17780 9602
rect 16156 9314 16212 9324
rect 17276 9380 17332 9390
rect 16716 9156 16772 9166
rect 16716 9062 16772 9100
rect 15484 8372 16324 8428
rect 16268 8370 16324 8372
rect 16268 8318 16270 8370
rect 16322 8318 16324 8370
rect 16268 8306 16324 8318
rect 17276 8146 17332 9324
rect 17724 9154 17780 9550
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17724 9090 17780 9102
rect 17836 9042 17892 10556
rect 18620 10610 19012 10612
rect 18620 10558 18622 10610
rect 18674 10558 19012 10610
rect 18620 10556 19012 10558
rect 18620 10546 18676 10556
rect 18956 9940 19012 10556
rect 19292 10610 19572 10612
rect 19292 10558 19294 10610
rect 19346 10558 19572 10610
rect 19292 10556 19572 10558
rect 19292 10546 19348 10556
rect 19516 10052 19572 10556
rect 19516 9986 19572 9996
rect 19404 9940 19460 9950
rect 18956 9938 19460 9940
rect 18956 9886 18958 9938
rect 19010 9886 19406 9938
rect 19458 9886 19460 9938
rect 18956 9884 19460 9886
rect 18956 9874 19012 9884
rect 19404 9874 19460 9884
rect 17836 8990 17838 9042
rect 17890 8990 17892 9042
rect 17836 8978 17892 8990
rect 18508 9602 18564 9614
rect 18508 9550 18510 9602
rect 18562 9550 18564 9602
rect 18508 8428 18564 9550
rect 19628 8428 19684 11342
rect 20076 11396 20132 11406
rect 20076 11302 20132 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20412 9156 20468 11902
rect 21196 10836 21252 12238
rect 21196 10770 21252 10780
rect 21532 10834 21588 12798
rect 21756 12628 21812 13694
rect 23212 13186 23268 13804
rect 23212 13134 23214 13186
rect 23266 13134 23268 13186
rect 23212 13122 23268 13134
rect 22540 12964 22596 12974
rect 22652 12964 22708 12974
rect 22596 12962 22708 12964
rect 22596 12910 22654 12962
rect 22706 12910 22708 12962
rect 22596 12908 22708 12910
rect 21756 12572 21924 12628
rect 21868 11508 21924 12572
rect 22316 11508 22372 11518
rect 21868 11506 22372 11508
rect 21868 11454 22318 11506
rect 22370 11454 22372 11506
rect 21868 11452 22372 11454
rect 22316 11442 22372 11452
rect 21532 10782 21534 10834
rect 21586 10782 21588 10834
rect 21532 10770 21588 10782
rect 21980 11172 22036 11182
rect 20412 9090 20468 9100
rect 20972 10052 21028 10062
rect 20972 8930 21028 9996
rect 21980 9154 22036 11116
rect 22540 10612 22596 12908
rect 22652 12898 22708 12908
rect 23436 12178 23492 12190
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 23436 11060 23492 12126
rect 23548 11282 23604 15148
rect 23660 14644 23716 15262
rect 24220 15314 24276 16716
rect 24220 15262 24222 15314
rect 24274 15262 24276 15314
rect 24220 15250 24276 15262
rect 25452 16660 25508 16670
rect 24444 14644 24500 14654
rect 23660 14642 24500 14644
rect 23660 14590 24446 14642
rect 24498 14590 24500 14642
rect 23660 14588 24500 14590
rect 24444 14578 24500 14588
rect 25452 14418 25508 16604
rect 25788 15204 25844 16830
rect 25788 15138 25844 15148
rect 26124 16884 26180 16894
rect 25452 14366 25454 14418
rect 25506 14366 25508 14418
rect 25452 14354 25508 14366
rect 23996 13860 24052 13870
rect 23996 13766 24052 13804
rect 23772 13748 23828 13758
rect 23772 12964 23828 13692
rect 26124 13748 26180 16828
rect 26236 15986 26292 18174
rect 26348 17444 26404 18396
rect 26796 18228 26852 22428
rect 27020 22372 27076 22382
rect 27692 22372 27748 22382
rect 26908 22370 27748 22372
rect 26908 22318 27022 22370
rect 27074 22318 27694 22370
rect 27746 22318 27748 22370
rect 26908 22316 27748 22318
rect 26908 20356 26964 22316
rect 27020 22306 27076 22316
rect 27692 22306 27748 22316
rect 29260 22372 29316 25452
rect 29708 27076 29764 27086
rect 29708 25506 29764 27020
rect 30492 27076 30548 28702
rect 32172 28754 33348 28756
rect 32172 28702 33294 28754
rect 33346 28702 33348 28754
rect 32172 28700 33348 28702
rect 31500 28532 31556 28542
rect 31500 28438 31556 28476
rect 30492 27010 30548 27020
rect 32172 27074 32228 28700
rect 33292 28690 33348 28700
rect 33404 28756 33460 28766
rect 32844 27300 32900 27310
rect 32172 27022 32174 27074
rect 32226 27022 32228 27074
rect 32172 27010 32228 27022
rect 32732 27298 32900 27300
rect 32732 27246 32846 27298
rect 32898 27246 32900 27298
rect 32732 27244 32900 27246
rect 32732 27074 32788 27244
rect 32844 27234 32900 27244
rect 32732 27022 32734 27074
rect 32786 27022 32788 27074
rect 32732 27010 32788 27022
rect 29820 26962 29876 26974
rect 29820 26910 29822 26962
rect 29874 26910 29876 26962
rect 29820 26852 29876 26910
rect 33180 26962 33236 26974
rect 33180 26910 33182 26962
rect 33234 26910 33236 26962
rect 29820 26786 29876 26796
rect 30716 26852 30772 26862
rect 29708 25454 29710 25506
rect 29762 25454 29764 25506
rect 29708 25442 29764 25454
rect 30156 25284 30212 25294
rect 30156 24834 30212 25228
rect 30716 24946 30772 26796
rect 33180 26292 33236 26910
rect 33180 26198 33236 26236
rect 33404 26068 33460 28700
rect 33516 27298 33572 29260
rect 33964 29316 34020 30158
rect 34748 30210 34804 30222
rect 34748 30158 34750 30210
rect 34802 30158 34804 30210
rect 34524 29986 34580 29998
rect 34524 29934 34526 29986
rect 34578 29934 34580 29986
rect 33964 29250 34020 29260
rect 34188 29764 34244 29774
rect 34188 29314 34244 29708
rect 34188 29262 34190 29314
rect 34242 29262 34244 29314
rect 34188 29250 34244 29262
rect 34300 28532 34356 28542
rect 34300 28438 34356 28476
rect 33516 27246 33518 27298
rect 33570 27246 33572 27298
rect 33516 26964 33572 27246
rect 33964 27858 34020 27870
rect 33964 27806 33966 27858
rect 34018 27806 34020 27858
rect 33964 26964 34020 27806
rect 33516 26962 34020 26964
rect 33516 26910 33518 26962
rect 33570 26910 34020 26962
rect 33516 26908 34020 26910
rect 34412 26964 34468 26974
rect 33516 26898 33572 26908
rect 33404 26012 33572 26068
rect 30716 24894 30718 24946
rect 30770 24894 30772 24946
rect 30716 24882 30772 24894
rect 32172 25282 32228 25294
rect 32172 25230 32174 25282
rect 32226 25230 32228 25282
rect 30156 24782 30158 24834
rect 30210 24782 30212 24834
rect 30156 24770 30212 24782
rect 32172 24834 32228 25230
rect 32172 24782 32174 24834
rect 32226 24782 32228 24834
rect 32172 24770 32228 24782
rect 32732 25282 32788 25294
rect 32732 25230 32734 25282
rect 32786 25230 32788 25282
rect 32732 24836 32788 25230
rect 32844 25284 32900 25294
rect 32844 25190 32900 25228
rect 33180 24948 33236 24958
rect 33180 24854 33236 24892
rect 32732 24770 32788 24780
rect 30604 24724 30660 24734
rect 30268 23716 30324 23726
rect 30604 23716 30660 24668
rect 31724 24724 31780 24734
rect 31724 24630 31780 24668
rect 31276 24276 31332 24286
rect 30828 23940 30884 23950
rect 30828 23938 30996 23940
rect 30828 23886 30830 23938
rect 30882 23886 30996 23938
rect 30828 23884 30996 23886
rect 30828 23874 30884 23884
rect 30156 23714 30660 23716
rect 30156 23662 30270 23714
rect 30322 23662 30660 23714
rect 30156 23660 30660 23662
rect 30156 23042 30212 23660
rect 30268 23650 30324 23660
rect 30156 22990 30158 23042
rect 30210 22990 30212 23042
rect 30156 22978 30212 22990
rect 27244 22148 27300 22158
rect 28252 22148 28308 22158
rect 27244 22146 28084 22148
rect 27244 22094 27246 22146
rect 27298 22094 28084 22146
rect 27244 22092 28084 22094
rect 27244 22082 27300 22092
rect 28028 21810 28084 22092
rect 28252 22054 28308 22092
rect 29036 22146 29092 22158
rect 29036 22094 29038 22146
rect 29090 22094 29092 22146
rect 29036 22036 29092 22094
rect 29036 21970 29092 21980
rect 28028 21758 28030 21810
rect 28082 21758 28084 21810
rect 28028 21746 28084 21758
rect 29148 21588 29204 21598
rect 29260 21588 29316 22316
rect 30940 22372 30996 23884
rect 31276 23938 31332 24220
rect 31276 23886 31278 23938
rect 31330 23886 31332 23938
rect 31276 23874 31332 23886
rect 33516 23826 33572 26012
rect 33628 25396 33684 25406
rect 33628 25302 33684 25340
rect 33740 25172 33796 26908
rect 33516 23774 33518 23826
rect 33570 23774 33572 23826
rect 33516 23762 33572 23774
rect 33628 24612 33684 24622
rect 33740 24612 33796 25116
rect 33628 24610 33796 24612
rect 33628 24558 33630 24610
rect 33682 24558 33796 24610
rect 33628 24556 33796 24558
rect 34076 24610 34132 24622
rect 34076 24558 34078 24610
rect 34130 24558 34132 24610
rect 33516 23604 33572 23614
rect 33180 23042 33236 23054
rect 33180 22990 33182 23042
rect 33234 22990 33236 23042
rect 33180 22930 33236 22990
rect 33180 22878 33182 22930
rect 33234 22878 33236 22930
rect 30940 22306 30996 22316
rect 32172 22370 32228 22382
rect 32172 22318 32174 22370
rect 32226 22318 32228 22370
rect 29596 22148 29652 22158
rect 29596 22054 29652 22092
rect 32060 21812 32116 21822
rect 32060 21718 32116 21756
rect 29148 21586 29316 21588
rect 29148 21534 29150 21586
rect 29202 21534 29316 21586
rect 29148 21532 29316 21534
rect 29596 21588 29652 21598
rect 29148 21522 29204 21532
rect 29596 21494 29652 21532
rect 28812 21362 28868 21374
rect 28812 21310 28814 21362
rect 28866 21310 28868 21362
rect 27580 20802 27636 20814
rect 27580 20750 27582 20802
rect 27634 20750 27636 20802
rect 27020 20580 27076 20590
rect 27076 20524 27188 20580
rect 27020 20514 27076 20524
rect 26908 20300 27076 20356
rect 27020 19796 27076 20300
rect 27132 20188 27188 20524
rect 27132 20132 27300 20188
rect 27020 19730 27076 19740
rect 27244 20018 27300 20132
rect 27244 19966 27246 20018
rect 27298 19966 27300 20018
rect 27132 19124 27188 19134
rect 27132 19030 27188 19068
rect 26796 18162 26852 18172
rect 27244 18562 27300 19966
rect 27244 18510 27246 18562
rect 27298 18510 27300 18562
rect 26348 17378 26404 17388
rect 26908 17444 26964 17454
rect 26908 17350 26964 17388
rect 27244 16884 27300 18510
rect 27580 17444 27636 20750
rect 27692 20578 27748 20590
rect 27692 20526 27694 20578
rect 27746 20526 27748 20578
rect 27692 20188 27748 20526
rect 27692 20132 28084 20188
rect 27804 20018 27860 20030
rect 27804 19966 27806 20018
rect 27858 19966 27860 20018
rect 27636 17388 27748 17444
rect 27580 17350 27636 17388
rect 27244 16818 27300 16828
rect 26236 15934 26238 15986
rect 26290 15934 26292 15986
rect 26236 15922 26292 15934
rect 27020 15876 27076 15886
rect 27020 15782 27076 15820
rect 27244 15316 27300 15326
rect 27244 14306 27300 15260
rect 27692 15316 27748 17388
rect 27804 17108 27860 19966
rect 27804 17042 27860 17052
rect 28028 17106 28084 20132
rect 28812 19124 28868 21310
rect 32172 21252 32228 22318
rect 32284 22372 32340 22382
rect 32508 22372 32564 22382
rect 32844 22372 32900 22382
rect 33180 22372 33236 22878
rect 32340 22370 33236 22372
rect 32340 22318 32510 22370
rect 32562 22318 32846 22370
rect 32898 22318 33236 22370
rect 32340 22316 33236 22318
rect 33516 22370 33572 23548
rect 33628 22930 33684 24556
rect 34076 24276 34132 24558
rect 34076 24210 34132 24220
rect 34300 24164 34356 24174
rect 34300 24070 34356 24108
rect 33628 22878 33630 22930
rect 33682 22878 33684 22930
rect 33628 22866 33684 22878
rect 33740 23042 33796 23054
rect 33740 22990 33742 23042
rect 33794 22990 33796 23042
rect 33516 22318 33518 22370
rect 33570 22318 33572 22370
rect 32284 22306 32340 22316
rect 32508 22306 32564 22316
rect 32844 22306 32900 22316
rect 33516 22306 33572 22318
rect 33180 21812 33236 21822
rect 33180 21718 33236 21756
rect 33404 21588 33460 21598
rect 33740 21588 33796 22990
rect 34076 23042 34132 23054
rect 34076 22990 34078 23042
rect 34130 22990 34132 23042
rect 34076 21700 34132 22990
rect 34076 21634 34132 21644
rect 33404 21586 33796 21588
rect 33404 21534 33406 21586
rect 33458 21534 33796 21586
rect 33404 21532 33796 21534
rect 32620 21364 32676 21374
rect 32620 21270 32676 21308
rect 32172 21186 32228 21196
rect 30940 20802 30996 20814
rect 30940 20750 30942 20802
rect 30994 20750 30996 20802
rect 30044 20132 30100 20142
rect 28812 19058 28868 19068
rect 29708 20130 30100 20132
rect 29708 20078 30046 20130
rect 30098 20078 30100 20130
rect 29708 20076 30100 20078
rect 29036 19010 29092 19022
rect 29036 18958 29038 19010
rect 29090 18958 29092 19010
rect 29036 18564 29092 18958
rect 29036 18498 29092 18508
rect 28588 18228 28644 18238
rect 28588 17668 28644 18172
rect 29148 17668 29204 17678
rect 28588 17666 29204 17668
rect 28588 17614 28590 17666
rect 28642 17614 29150 17666
rect 29202 17614 29204 17666
rect 28588 17612 29204 17614
rect 28588 17602 28644 17612
rect 29148 17602 29204 17612
rect 28028 17054 28030 17106
rect 28082 17054 28084 17106
rect 28028 17042 28084 17054
rect 28812 16996 28868 17006
rect 28812 16902 28868 16940
rect 29708 16210 29764 20076
rect 30044 20066 30100 20076
rect 30940 20132 30996 20750
rect 31388 20804 31444 20814
rect 31388 20710 31444 20748
rect 33404 20188 33460 21532
rect 33964 21252 34020 21262
rect 33740 20578 33796 20590
rect 33740 20526 33742 20578
rect 33794 20526 33796 20578
rect 33740 20242 33796 20526
rect 33740 20190 33742 20242
rect 33794 20190 33796 20242
rect 30940 20066 30996 20076
rect 32620 20132 32676 20142
rect 33404 20132 33572 20188
rect 33740 20178 33796 20190
rect 32508 20020 32564 20030
rect 30828 19796 30884 19806
rect 30828 19702 30884 19740
rect 32172 19348 32228 19358
rect 32172 19234 32228 19292
rect 32172 19182 32174 19234
rect 32226 19182 32228 19234
rect 32172 19170 32228 19182
rect 29820 19010 29876 19022
rect 29820 18958 29822 19010
rect 29874 18958 29876 19010
rect 29820 17332 29876 18958
rect 30716 18452 30772 18462
rect 30716 18358 30772 18396
rect 32508 17780 32564 19964
rect 32508 17686 32564 17724
rect 32620 19236 32676 20076
rect 33516 20020 33572 20132
rect 33516 19926 33572 19964
rect 33964 19346 34020 21196
rect 34412 21026 34468 26908
rect 34524 25396 34580 29934
rect 34748 29652 34804 30158
rect 35868 30210 35924 30222
rect 35868 30158 35870 30210
rect 35922 30158 35924 30210
rect 35868 30100 35924 30158
rect 35924 30044 36148 30100
rect 35868 30034 35924 30044
rect 34804 29596 35140 29652
rect 34748 29586 34804 29596
rect 35084 28644 35140 29596
rect 36092 29650 36148 30044
rect 36092 29598 36094 29650
rect 36146 29598 36148 29650
rect 36092 29586 36148 29598
rect 36764 29650 36820 30268
rect 36764 29598 36766 29650
rect 36818 29598 36820 29650
rect 36764 29586 36820 29598
rect 35308 29540 35364 29550
rect 35308 29446 35364 29484
rect 36540 29316 36596 29326
rect 36540 29222 36596 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 36876 28866 36932 30380
rect 36988 30210 37044 30718
rect 36988 30158 36990 30210
rect 37042 30158 37044 30210
rect 36988 29316 37044 30158
rect 37324 30100 37380 31726
rect 37436 30996 37492 31948
rect 37436 30994 37604 30996
rect 37436 30942 37438 30994
rect 37490 30942 37604 30994
rect 37436 30940 37604 30942
rect 37436 30930 37492 30940
rect 37548 30770 37604 30940
rect 37548 30718 37550 30770
rect 37602 30718 37604 30770
rect 37548 30706 37604 30718
rect 37660 30212 37716 30222
rect 37772 30212 37828 33404
rect 38444 33394 38500 33404
rect 38108 32564 38164 32574
rect 38108 32004 38164 32508
rect 38556 31948 38612 34748
rect 39116 34738 39172 34748
rect 39452 33236 39508 33246
rect 39228 33234 39508 33236
rect 39228 33182 39454 33234
rect 39506 33182 39508 33234
rect 39228 33180 39508 33182
rect 39116 32562 39172 32574
rect 39116 32510 39118 32562
rect 39170 32510 39172 32562
rect 39116 32452 39172 32510
rect 39116 32386 39172 32396
rect 39228 31948 39284 33180
rect 39452 33170 39508 33180
rect 40348 32788 40404 34974
rect 40236 32732 40404 32788
rect 39900 32564 39956 32574
rect 39900 32470 39956 32508
rect 38108 31892 38276 31948
rect 38220 31778 38276 31892
rect 38220 31726 38222 31778
rect 38274 31726 38276 31778
rect 38220 31714 38276 31726
rect 38332 31892 38612 31948
rect 39116 31892 39284 31948
rect 39340 32338 39396 32350
rect 39340 32286 39342 32338
rect 39394 32286 39396 32338
rect 39340 31948 39396 32286
rect 40236 31948 40292 32732
rect 40348 32564 40404 32574
rect 40348 32562 40516 32564
rect 40348 32510 40350 32562
rect 40402 32510 40516 32562
rect 40348 32508 40516 32510
rect 40348 32498 40404 32508
rect 40460 32452 40516 32508
rect 40460 32386 40516 32396
rect 39340 31892 39844 31948
rect 37884 30884 37940 30894
rect 37884 30790 37940 30828
rect 37660 30210 37828 30212
rect 37660 30158 37662 30210
rect 37714 30158 37828 30210
rect 37660 30156 37828 30158
rect 37660 30146 37716 30156
rect 37324 30034 37380 30044
rect 37548 29988 37604 29998
rect 37548 29650 37604 29932
rect 37548 29598 37550 29650
rect 37602 29598 37604 29650
rect 37548 29586 37604 29598
rect 36988 29250 37044 29260
rect 36876 28814 36878 28866
rect 36930 28814 36932 28866
rect 36876 28802 36932 28814
rect 35308 28756 35364 28766
rect 35308 28662 35364 28700
rect 34636 27858 34692 27870
rect 34636 27806 34638 27858
rect 34690 27806 34692 27858
rect 34636 27188 34692 27806
rect 34636 27122 34692 27132
rect 34972 27186 35028 27198
rect 34972 27134 34974 27186
rect 35026 27134 35028 27186
rect 34524 25330 34580 25340
rect 34972 23604 35028 27134
rect 35084 24948 35140 28588
rect 36316 28644 36372 28654
rect 36316 28550 36372 28588
rect 37660 28420 37716 28430
rect 37660 28326 37716 28364
rect 38332 28308 38388 31892
rect 38892 31106 38948 31118
rect 38892 31054 38894 31106
rect 38946 31054 38948 31106
rect 38892 30324 38948 31054
rect 39116 30436 39172 31892
rect 39116 30370 39172 30380
rect 39228 31666 39284 31678
rect 39228 31614 39230 31666
rect 39282 31614 39284 31666
rect 38892 30258 38948 30268
rect 37772 28252 38388 28308
rect 37660 28084 37716 28094
rect 37772 28084 37828 28252
rect 37660 28082 37828 28084
rect 37660 28030 37662 28082
rect 37714 28030 37828 28082
rect 37660 28028 37828 28030
rect 37660 28018 37716 28028
rect 36876 27970 36932 27982
rect 36876 27918 36878 27970
rect 36930 27918 36932 27970
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35980 26964 36036 26974
rect 35980 26870 36036 26908
rect 36876 26516 36932 27918
rect 38892 27970 38948 27982
rect 38892 27918 38894 27970
rect 38946 27918 38948 27970
rect 37884 27748 37940 27758
rect 36876 26450 36932 26460
rect 37772 27746 37940 27748
rect 37772 27694 37886 27746
rect 37938 27694 37940 27746
rect 37772 27692 37940 27694
rect 35644 26178 35700 26190
rect 35644 26126 35646 26178
rect 35698 26126 35700 26178
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35644 25172 35700 26126
rect 36988 25844 37044 25854
rect 35644 25106 35700 25116
rect 35980 25506 36036 25518
rect 35980 25454 35982 25506
rect 36034 25454 36036 25506
rect 35084 24052 35140 24892
rect 35308 24836 35364 24846
rect 35308 24742 35364 24780
rect 35980 24498 36036 25454
rect 36316 25508 36372 25518
rect 35980 24446 35982 24498
rect 36034 24446 36036 24498
rect 35980 24434 36036 24446
rect 36092 25172 36148 25182
rect 36316 25172 36372 25452
rect 36148 25116 36596 25172
rect 36092 24946 36148 25116
rect 36092 24894 36094 24946
rect 36146 24894 36148 24946
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 23938 35140 23996
rect 35756 24052 35812 24062
rect 35756 23958 35812 23996
rect 36092 24052 36148 24894
rect 36540 24946 36596 25116
rect 36540 24894 36542 24946
rect 36594 24894 36596 24946
rect 36540 24882 36596 24894
rect 36876 24612 36932 24622
rect 36652 24610 36932 24612
rect 36652 24558 36878 24610
rect 36930 24558 36932 24610
rect 36652 24556 36932 24558
rect 36652 24498 36708 24556
rect 36876 24546 36932 24556
rect 36652 24446 36654 24498
rect 36706 24446 36708 24498
rect 36652 24434 36708 24446
rect 36988 24162 37044 25788
rect 37100 25508 37156 25518
rect 37100 25414 37156 25452
rect 37772 25506 37828 27692
rect 37884 27682 37940 27692
rect 37996 27188 38052 27198
rect 37996 27094 38052 27132
rect 38780 26516 38836 26526
rect 38780 26422 38836 26460
rect 37772 25454 37774 25506
rect 37826 25454 37828 25506
rect 37772 25442 37828 25454
rect 38668 26290 38724 26302
rect 38668 26238 38670 26290
rect 38722 26238 38724 26290
rect 38668 24948 38724 26238
rect 38892 25844 38948 27918
rect 38892 25778 38948 25788
rect 38724 24892 39172 24948
rect 38668 24882 38724 24892
rect 36988 24110 36990 24162
rect 37042 24110 37044 24162
rect 36988 24098 37044 24110
rect 37884 24834 37940 24846
rect 37884 24782 37886 24834
rect 37938 24782 37940 24834
rect 37884 24164 37940 24782
rect 39116 24724 39172 24892
rect 39228 24724 39284 31614
rect 39788 30100 39844 31892
rect 40012 31892 40292 31948
rect 39900 30100 39956 30110
rect 39788 30098 39956 30100
rect 39788 30046 39902 30098
rect 39954 30046 39956 30098
rect 39788 30044 39956 30046
rect 39900 30034 39956 30044
rect 39900 29428 39956 29438
rect 39900 29334 39956 29372
rect 39788 29316 39844 29326
rect 39788 28082 39844 29260
rect 40012 28642 40068 31892
rect 40348 31890 40404 31902
rect 40348 31838 40350 31890
rect 40402 31838 40404 31890
rect 40012 28590 40014 28642
rect 40066 28590 40068 28642
rect 40012 28578 40068 28590
rect 40236 29652 40292 29662
rect 39788 28030 39790 28082
rect 39842 28030 39844 28082
rect 39788 28018 39844 28030
rect 39900 28420 39956 28430
rect 39900 27298 39956 28364
rect 39900 27246 39902 27298
rect 39954 27246 39956 27298
rect 39900 27234 39956 27246
rect 40236 28082 40292 29596
rect 40236 28030 40238 28082
rect 40290 28030 40292 28082
rect 40124 27076 40180 27086
rect 40236 27076 40292 28030
rect 40124 27074 40292 27076
rect 40124 27022 40126 27074
rect 40178 27022 40292 27074
rect 40124 27020 40292 27022
rect 40124 27010 40180 27020
rect 39340 26962 39396 26974
rect 39340 26910 39342 26962
rect 39394 26910 39396 26962
rect 39340 25732 39396 26910
rect 39340 25666 39396 25676
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 25508 39956 26126
rect 39900 25452 40180 25508
rect 40012 25282 40068 25294
rect 40012 25230 40014 25282
rect 40066 25230 40068 25282
rect 40012 25172 40068 25230
rect 39340 25116 40068 25172
rect 39340 24946 39396 25116
rect 39340 24894 39342 24946
rect 39394 24894 39396 24946
rect 39340 24882 39396 24894
rect 39900 24724 39956 24734
rect 40124 24724 40180 25452
rect 39228 24668 39844 24724
rect 39116 24630 39172 24668
rect 37884 24098 37940 24108
rect 36204 24052 36260 24062
rect 36092 24050 36260 24052
rect 36092 23998 36206 24050
rect 36258 23998 36260 24050
rect 36092 23996 36260 23998
rect 35084 23886 35086 23938
rect 35138 23886 35140 23938
rect 35084 23874 35140 23886
rect 34972 23538 35028 23548
rect 35196 23714 35252 23726
rect 35196 23662 35198 23714
rect 35250 23662 35252 23714
rect 35084 23266 35140 23278
rect 35084 23214 35086 23266
rect 35138 23214 35140 23266
rect 34972 23156 35028 23166
rect 34412 20974 34414 21026
rect 34466 20974 34468 21026
rect 34412 20962 34468 20974
rect 34636 21586 34692 21598
rect 34636 21534 34638 21586
rect 34690 21534 34692 21586
rect 34636 21026 34692 21534
rect 34636 20974 34638 21026
rect 34690 20974 34692 21026
rect 34636 20962 34692 20974
rect 34860 20916 34916 20926
rect 34972 20916 35028 23100
rect 35084 22596 35140 23214
rect 35196 23044 35252 23662
rect 36092 23156 36148 23996
rect 36204 23986 36260 23996
rect 37772 23714 37828 23726
rect 37772 23662 37774 23714
rect 37826 23662 37828 23714
rect 36092 23062 36148 23100
rect 36764 23154 36820 23166
rect 36764 23102 36766 23154
rect 36818 23102 36820 23154
rect 35196 22988 35812 23044
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22530 35140 22540
rect 35756 22258 35812 22988
rect 35756 22206 35758 22258
rect 35810 22206 35812 22258
rect 35756 22194 35812 22206
rect 36540 22146 36596 22158
rect 36540 22094 36542 22146
rect 36594 22094 36596 22146
rect 34860 20914 35028 20916
rect 34860 20862 34862 20914
rect 34914 20862 35028 20914
rect 34860 20860 35028 20862
rect 35084 21586 35140 21598
rect 35084 21534 35086 21586
rect 35138 21534 35140 21586
rect 34860 20850 34916 20860
rect 35084 20020 35140 21534
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 21026 35252 21038
rect 35196 20974 35198 21026
rect 35250 20974 35252 21026
rect 35196 20916 35252 20974
rect 35196 20822 35252 20860
rect 35084 19954 35140 19964
rect 35868 20130 35924 20142
rect 35868 20078 35870 20130
rect 35922 20078 35924 20130
rect 33964 19294 33966 19346
rect 34018 19294 34020 19346
rect 33964 19282 34020 19294
rect 35084 19794 35140 19806
rect 35084 19742 35086 19794
rect 35138 19742 35140 19794
rect 33068 19236 33124 19246
rect 32620 19234 33124 19236
rect 32620 19182 32622 19234
rect 32674 19182 33070 19234
rect 33122 19182 33124 19234
rect 32620 19180 33124 19182
rect 32620 18340 32676 19180
rect 33068 19170 33124 19180
rect 34972 19124 35028 19134
rect 34972 19030 35028 19068
rect 32396 17668 32452 17678
rect 32284 17612 32396 17668
rect 29820 17276 30324 17332
rect 30044 17108 30100 17118
rect 30044 16770 30100 17052
rect 30044 16718 30046 16770
rect 30098 16718 30100 16770
rect 30044 16706 30100 16718
rect 30268 16324 30324 17276
rect 31052 16996 31108 17006
rect 31052 16902 31108 16940
rect 31500 16772 31556 16782
rect 30380 16324 30436 16334
rect 30268 16322 30436 16324
rect 30268 16270 30382 16322
rect 30434 16270 30436 16322
rect 30268 16268 30436 16270
rect 30380 16258 30436 16268
rect 29708 16158 29710 16210
rect 29762 16158 29764 16210
rect 29708 16146 29764 16158
rect 29932 16100 29988 16110
rect 30268 16100 30324 16110
rect 29932 16098 30324 16100
rect 29932 16046 29934 16098
rect 29986 16046 30270 16098
rect 30322 16046 30324 16098
rect 29932 16044 30324 16046
rect 27692 15250 27748 15260
rect 28588 15874 28644 15886
rect 28588 15822 28590 15874
rect 28642 15822 28644 15874
rect 28588 15316 28644 15822
rect 28700 15876 28756 15886
rect 28700 15426 28756 15820
rect 28700 15374 28702 15426
rect 28754 15374 28756 15426
rect 28700 15362 28756 15374
rect 28588 15250 28644 15260
rect 29932 15316 29988 16044
rect 30268 16034 30324 16044
rect 31500 16098 31556 16716
rect 31500 16046 31502 16098
rect 31554 16046 31556 16098
rect 31500 16034 31556 16046
rect 31948 16098 32004 16110
rect 31948 16046 31950 16098
rect 32002 16046 32004 16098
rect 29932 15222 29988 15260
rect 30716 15652 30772 15662
rect 27580 15204 27636 15214
rect 27580 15110 27636 15148
rect 30716 15202 30772 15596
rect 30716 15150 30718 15202
rect 30770 15150 30772 15202
rect 30716 15138 30772 15150
rect 29932 14644 29988 14654
rect 29708 14642 29988 14644
rect 29708 14590 29934 14642
rect 29986 14590 29988 14642
rect 29708 14588 29988 14590
rect 27244 14254 27246 14306
rect 27298 14254 27300 14306
rect 26124 13654 26180 13692
rect 26796 13746 26852 13758
rect 26796 13694 26798 13746
rect 26850 13694 26852 13746
rect 24780 13522 24836 13534
rect 24780 13470 24782 13522
rect 24834 13470 24836 13522
rect 24780 13188 24836 13470
rect 24780 13122 24836 13132
rect 23772 12962 23940 12964
rect 23772 12910 23774 12962
rect 23826 12910 23940 12962
rect 23772 12908 23940 12910
rect 23772 12898 23828 12908
rect 23884 12178 23940 12908
rect 23884 12126 23886 12178
rect 23938 12126 23940 12178
rect 23884 12114 23940 12126
rect 24332 12962 24388 12974
rect 24332 12910 24334 12962
rect 24386 12910 24388 12962
rect 24332 11508 24388 12910
rect 26796 12964 26852 13694
rect 26908 13188 26964 13198
rect 26964 13132 27076 13188
rect 26908 13122 26964 13132
rect 26796 12908 26964 12964
rect 26796 12740 26852 12750
rect 26796 12646 26852 12684
rect 25900 12290 25956 12302
rect 25900 12238 25902 12290
rect 25954 12238 25956 12290
rect 24332 11442 24388 11452
rect 25116 11954 25172 11966
rect 25116 11902 25118 11954
rect 25170 11902 25172 11954
rect 23548 11230 23550 11282
rect 23602 11230 23604 11282
rect 23548 11218 23604 11230
rect 23548 11060 23604 11070
rect 23436 11004 23548 11060
rect 23548 10994 23604 11004
rect 24332 11060 24388 11070
rect 22652 10836 22708 10846
rect 22652 10742 22708 10780
rect 22540 10518 22596 10556
rect 22316 10388 22372 10398
rect 22316 10386 22596 10388
rect 22316 10334 22318 10386
rect 22370 10334 22596 10386
rect 22316 10332 22596 10334
rect 22316 10322 22372 10332
rect 22540 10052 22596 10332
rect 22540 9996 23268 10052
rect 23212 9714 23268 9996
rect 24332 9938 24388 11004
rect 25116 10724 25172 11902
rect 25900 11620 25956 12238
rect 25900 11554 25956 11564
rect 25676 11508 25732 11518
rect 25676 11414 25732 11452
rect 25116 10658 25172 10668
rect 26236 10724 26292 10734
rect 26236 10630 26292 10668
rect 26908 10500 26964 12908
rect 27020 11282 27076 13132
rect 27244 12964 27300 14254
rect 29484 14308 29540 14318
rect 27356 13860 27412 13870
rect 29036 13860 29092 13870
rect 27356 13186 27412 13804
rect 28700 13858 29092 13860
rect 28700 13806 29038 13858
rect 29090 13806 29092 13858
rect 28700 13804 29092 13806
rect 28588 13748 28644 13758
rect 27356 13134 27358 13186
rect 27410 13134 27412 13186
rect 27356 13122 27412 13134
rect 28252 13636 28308 13646
rect 27804 12964 27860 12974
rect 27244 12962 27860 12964
rect 27244 12910 27806 12962
rect 27858 12910 27860 12962
rect 27244 12908 27860 12910
rect 27692 12740 27748 12750
rect 27692 12646 27748 12684
rect 27580 11620 27636 11630
rect 27580 11526 27636 11564
rect 27020 11230 27022 11282
rect 27074 11230 27076 11282
rect 27020 11218 27076 11230
rect 27580 11396 27636 11406
rect 27804 11396 27860 12908
rect 28252 12178 28308 13580
rect 28252 12126 28254 12178
rect 28306 12126 28308 12178
rect 28252 12114 28308 12126
rect 28588 12178 28644 13692
rect 28588 12126 28590 12178
rect 28642 12126 28644 12178
rect 28588 12114 28644 12126
rect 28700 11732 28756 13804
rect 29036 13794 29092 13804
rect 29260 12964 29316 12974
rect 29260 12870 29316 12908
rect 29484 12402 29540 14252
rect 29708 12962 29764 14588
rect 29932 14578 29988 14588
rect 31948 14644 32004 16046
rect 32284 15540 32340 17612
rect 32396 17602 32452 17612
rect 32620 16772 32676 18284
rect 33516 18452 33572 18462
rect 33516 17778 33572 18396
rect 33516 17726 33518 17778
rect 33570 17726 33572 17778
rect 33516 17714 33572 17726
rect 33628 17780 33684 17790
rect 32620 16706 32676 16716
rect 33180 16882 33236 16894
rect 33180 16830 33182 16882
rect 33234 16830 33236 16882
rect 33180 16772 33236 16830
rect 32060 15484 32340 15540
rect 32060 15426 32116 15484
rect 32060 15374 32062 15426
rect 32114 15374 32116 15426
rect 32060 15362 32116 15374
rect 31948 14578 32004 14588
rect 32396 14532 32452 14542
rect 32732 14532 32788 14542
rect 32396 14530 33012 14532
rect 32396 14478 32398 14530
rect 32450 14478 32734 14530
rect 32786 14478 33012 14530
rect 32396 14476 33012 14478
rect 32396 14466 32452 14476
rect 32732 14466 32788 14476
rect 29820 14420 29876 14430
rect 29820 13970 29876 14364
rect 30940 14420 30996 14430
rect 30940 14326 30996 14364
rect 32844 14308 32900 14318
rect 32844 14214 32900 14252
rect 29820 13918 29822 13970
rect 29874 13918 29876 13970
rect 29820 13906 29876 13918
rect 32060 13860 32116 13870
rect 32060 13766 32116 13804
rect 31052 13636 31108 13646
rect 31052 13542 31108 13580
rect 32060 13076 32116 13086
rect 29708 12910 29710 12962
rect 29762 12910 29764 12962
rect 29708 12898 29764 12910
rect 30044 12964 30100 12974
rect 29484 12350 29486 12402
rect 29538 12350 29540 12402
rect 29484 12338 29540 12350
rect 30044 12180 30100 12908
rect 27580 11394 27860 11396
rect 27580 11342 27582 11394
rect 27634 11342 27860 11394
rect 27580 11340 27860 11342
rect 28476 11676 28756 11732
rect 28924 11954 28980 11966
rect 28924 11902 28926 11954
rect 28978 11902 28980 11954
rect 27356 10500 27412 10510
rect 26908 10498 27412 10500
rect 26908 10446 27358 10498
rect 27410 10446 27412 10498
rect 26908 10444 27412 10446
rect 27356 10434 27412 10444
rect 24332 9886 24334 9938
rect 24386 9886 24388 9938
rect 24332 9874 24388 9886
rect 27580 9828 27636 11340
rect 27580 9734 27636 9772
rect 28028 10498 28084 10510
rect 28028 10446 28030 10498
rect 28082 10446 28084 10498
rect 28028 9828 28084 10446
rect 28476 10050 28532 11676
rect 28924 10724 28980 11902
rect 30044 11394 30100 12124
rect 32060 12178 32116 13020
rect 32732 12852 32788 12862
rect 32732 12758 32788 12796
rect 32060 12126 32062 12178
rect 32114 12126 32116 12178
rect 32060 12114 32116 12126
rect 32172 12738 32228 12750
rect 32172 12686 32174 12738
rect 32226 12686 32228 12738
rect 30044 11342 30046 11394
rect 30098 11342 30100 11394
rect 30044 11330 30100 11342
rect 30716 11394 30772 11406
rect 30716 11342 30718 11394
rect 30770 11342 30772 11394
rect 30044 10724 30100 10734
rect 28924 10722 30100 10724
rect 28924 10670 30046 10722
rect 30098 10670 30100 10722
rect 28924 10668 30100 10670
rect 30044 10658 30100 10668
rect 30156 10724 30212 10734
rect 30156 10052 30212 10668
rect 30716 10500 30772 11342
rect 32172 10724 32228 12686
rect 32620 12180 32676 12190
rect 32620 10834 32676 12124
rect 32620 10782 32622 10834
rect 32674 10782 32676 10834
rect 32620 10770 32676 10782
rect 32172 10658 32228 10668
rect 32956 10612 33012 14476
rect 33180 13748 33236 16716
rect 33628 13972 33684 17724
rect 34636 17780 34692 17790
rect 34636 17686 34692 17724
rect 35084 17668 35140 19742
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35868 18452 35924 20078
rect 35868 18386 35924 18396
rect 35308 18340 35364 18350
rect 35308 18246 35364 18284
rect 36204 18340 36260 18350
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 17602 35140 17612
rect 35420 17780 35476 17790
rect 35420 17668 35476 17724
rect 35420 17666 35588 17668
rect 35420 17614 35422 17666
rect 35474 17614 35588 17666
rect 35420 17612 35588 17614
rect 35420 17602 35476 17612
rect 35532 16996 35588 17612
rect 35644 17444 35700 17454
rect 35644 17442 35812 17444
rect 35644 17390 35646 17442
rect 35698 17390 35812 17442
rect 35644 17388 35812 17390
rect 35644 17378 35700 17388
rect 35756 17220 35812 17388
rect 35756 17164 36148 17220
rect 36092 17106 36148 17164
rect 36092 17054 36094 17106
rect 36146 17054 36148 17106
rect 36092 17042 36148 17054
rect 33852 16882 33908 16894
rect 33852 16830 33854 16882
rect 33906 16830 33908 16882
rect 33852 15204 33908 16830
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35532 16098 35588 16940
rect 35532 16046 35534 16098
rect 35586 16046 35588 16098
rect 35532 16034 35588 16046
rect 36204 16884 36260 18284
rect 36540 17556 36596 22094
rect 36764 21924 36820 23102
rect 37100 23156 37156 23166
rect 37100 22484 37156 23100
rect 37772 22596 37828 23662
rect 37772 22530 37828 22540
rect 39228 23378 39284 23390
rect 39228 23326 39230 23378
rect 39282 23326 39284 23378
rect 37548 22484 37604 22494
rect 37100 22482 37604 22484
rect 37100 22430 37102 22482
rect 37154 22430 37550 22482
rect 37602 22430 37604 22482
rect 37100 22428 37604 22430
rect 37100 22418 37156 22428
rect 37548 22418 37604 22428
rect 37996 22482 38052 22494
rect 37996 22430 37998 22482
rect 38050 22430 38052 22482
rect 36764 21858 36820 21868
rect 37436 21812 37492 21822
rect 37436 21718 37492 21756
rect 37996 21588 38052 22430
rect 39004 22260 39060 22270
rect 39004 22166 39060 22204
rect 37996 21522 38052 21532
rect 38220 21924 38276 21934
rect 37772 21476 37828 21486
rect 36540 17490 36596 17500
rect 37212 20916 37268 20926
rect 37212 20244 37268 20860
rect 37772 20914 37828 21420
rect 38108 21362 38164 21374
rect 38108 21310 38110 21362
rect 38162 21310 38164 21362
rect 37772 20862 37774 20914
rect 37826 20862 37828 20914
rect 37772 20850 37828 20862
rect 37996 20916 38052 20926
rect 37996 20822 38052 20860
rect 38108 20188 38164 21310
rect 34412 15876 34468 15886
rect 34412 15782 34468 15820
rect 34972 15874 35028 15886
rect 34972 15822 34974 15874
rect 35026 15822 35028 15874
rect 34972 15428 35028 15822
rect 35308 15876 35364 15886
rect 35308 15782 35364 15820
rect 36204 15652 36260 16828
rect 36428 16996 36484 17006
rect 36428 16210 36484 16940
rect 37212 16884 37268 20188
rect 37996 20132 38164 20188
rect 37884 20020 37940 20030
rect 37884 17780 37940 19964
rect 37996 19572 38052 20132
rect 37996 19506 38052 19516
rect 38108 20018 38164 20030
rect 38108 19966 38110 20018
rect 38162 19966 38164 20018
rect 37996 19348 38052 19358
rect 37996 19254 38052 19292
rect 37996 17780 38052 17790
rect 37884 17778 38052 17780
rect 37884 17726 37998 17778
rect 38050 17726 38052 17778
rect 37884 17724 38052 17726
rect 37996 17714 38052 17724
rect 37884 17444 37940 17454
rect 37212 16790 37268 16828
rect 37660 16884 37716 16894
rect 37660 16790 37716 16828
rect 36876 16660 36932 16670
rect 36876 16658 37380 16660
rect 36876 16606 36878 16658
rect 36930 16606 37380 16658
rect 36876 16604 37380 16606
rect 36876 16594 36932 16604
rect 36428 16158 36430 16210
rect 36482 16158 36484 16210
rect 36428 16146 36484 16158
rect 37100 15874 37156 15886
rect 37100 15822 37102 15874
rect 37154 15822 37156 15874
rect 35980 15596 36596 15652
rect 35980 15538 36036 15596
rect 35980 15486 35982 15538
rect 36034 15486 36036 15538
rect 35980 15474 36036 15486
rect 36540 15540 36596 15596
rect 36540 15538 36820 15540
rect 36540 15486 36542 15538
rect 36594 15486 36820 15538
rect 36540 15484 36820 15486
rect 36540 15474 36596 15484
rect 35084 15428 35140 15438
rect 34972 15426 35140 15428
rect 34972 15374 35086 15426
rect 35138 15374 35140 15426
rect 34972 15372 35140 15374
rect 35084 15362 35140 15372
rect 36764 15314 36820 15484
rect 36764 15262 36766 15314
rect 36818 15262 36820 15314
rect 34076 15204 34132 15214
rect 33852 15202 34132 15204
rect 33852 15150 34078 15202
rect 34130 15150 34132 15202
rect 33852 15148 34132 15150
rect 34076 15138 34132 15148
rect 36316 15204 36372 15214
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34972 14644 35028 14654
rect 34972 14550 35028 14588
rect 36316 14418 36372 15148
rect 36316 14366 36318 14418
rect 36370 14366 36372 14418
rect 36316 14354 36372 14366
rect 36764 14084 36820 15262
rect 37100 15204 37156 15822
rect 37100 15138 37156 15148
rect 36876 14306 36932 14318
rect 36876 14254 36878 14306
rect 36930 14254 36932 14306
rect 36876 14196 36932 14254
rect 36876 14140 37156 14196
rect 36764 14028 37044 14084
rect 33516 13916 33684 13972
rect 36988 13970 37044 14028
rect 36988 13918 36990 13970
rect 37042 13918 37044 13970
rect 33068 13746 33236 13748
rect 33068 13694 33182 13746
rect 33234 13694 33236 13746
rect 33068 13692 33236 13694
rect 33068 13074 33124 13692
rect 33180 13682 33236 13692
rect 33292 13860 33348 13870
rect 33068 13022 33070 13074
rect 33122 13022 33124 13074
rect 33068 12180 33124 13022
rect 33292 12402 33348 13804
rect 33292 12350 33294 12402
rect 33346 12350 33348 12402
rect 33292 12338 33348 12350
rect 33516 13074 33572 13916
rect 35868 13860 35924 13870
rect 35868 13766 35924 13804
rect 33516 13022 33518 13074
rect 33570 13022 33572 13074
rect 33068 12114 33124 12124
rect 33516 12178 33572 13022
rect 33516 12126 33518 12178
rect 33570 12126 33572 12178
rect 33516 12114 33572 12126
rect 33628 13746 33684 13758
rect 33628 13694 33630 13746
rect 33682 13694 33684 13746
rect 33628 11508 33684 13694
rect 36652 13522 36708 13534
rect 36652 13470 36654 13522
rect 36706 13470 36708 13522
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 33964 13076 34020 13086
rect 33964 12982 34020 13020
rect 34972 12852 35028 12862
rect 34972 12758 35028 12796
rect 34076 12180 34132 12190
rect 34132 12124 34468 12180
rect 34076 12086 34132 12124
rect 33964 11508 34020 11518
rect 33628 11506 34020 11508
rect 33628 11454 33966 11506
rect 34018 11454 34020 11506
rect 33628 11452 34020 11454
rect 33964 11442 34020 11452
rect 33180 11170 33236 11182
rect 33180 11118 33182 11170
rect 33234 11118 33236 11170
rect 33180 10834 33236 11118
rect 33740 11172 33796 11182
rect 33740 11078 33796 11116
rect 33180 10782 33182 10834
rect 33234 10782 33236 10834
rect 33180 10770 33236 10782
rect 34412 10834 34468 12124
rect 34412 10782 34414 10834
rect 34466 10782 34468 10834
rect 34412 10770 34468 10782
rect 34748 12178 34804 12190
rect 34748 12126 34750 12178
rect 34802 12126 34804 12178
rect 33068 10612 33124 10622
rect 32956 10610 33124 10612
rect 32956 10558 33070 10610
rect 33122 10558 33124 10610
rect 32956 10556 33124 10558
rect 31164 10500 31220 10510
rect 30716 10498 31220 10500
rect 30716 10446 31166 10498
rect 31218 10446 31220 10498
rect 30716 10444 31220 10446
rect 31164 10434 31220 10444
rect 32060 10500 32116 10510
rect 32956 10500 33012 10556
rect 33068 10546 33124 10556
rect 32060 10498 33012 10500
rect 32060 10446 32062 10498
rect 32114 10446 33012 10498
rect 32060 10444 33012 10446
rect 34748 10500 34804 12126
rect 36652 12068 36708 13470
rect 36988 13524 37044 13918
rect 36988 13076 37044 13468
rect 37100 13412 37156 14140
rect 37324 13972 37380 16604
rect 37884 15986 37940 17388
rect 38108 16884 38164 19966
rect 38108 16818 38164 16828
rect 38220 16772 38276 21868
rect 38444 21812 38500 21822
rect 39228 21812 39284 23326
rect 39788 23378 39844 24668
rect 39956 24668 40180 24724
rect 39900 24630 39956 24668
rect 39788 23326 39790 23378
rect 39842 23326 39844 23378
rect 39788 23314 39844 23326
rect 39900 22596 39956 22606
rect 39900 22502 39956 22540
rect 40012 22484 40068 24668
rect 40124 23940 40180 23950
rect 40348 23940 40404 31838
rect 40460 29426 40516 29438
rect 40460 29374 40462 29426
rect 40514 29374 40516 29426
rect 40460 29316 40516 29374
rect 40572 29428 40628 36540
rect 40684 36530 40740 36540
rect 41692 36372 41748 36382
rect 40684 36370 41748 36372
rect 40684 36318 41694 36370
rect 41746 36318 41748 36370
rect 40684 36316 41748 36318
rect 40684 30210 40740 36316
rect 41692 36306 41748 36316
rect 40796 32452 40852 32462
rect 40852 32396 40964 32452
rect 40796 32386 40852 32396
rect 40684 30158 40686 30210
rect 40738 30158 40740 30210
rect 40684 30146 40740 30158
rect 40908 30210 40964 32396
rect 40908 30158 40910 30210
rect 40962 30158 40964 30210
rect 40908 29652 40964 30158
rect 41020 29988 41076 29998
rect 41020 29894 41076 29932
rect 41020 29652 41076 29662
rect 40964 29650 41076 29652
rect 40964 29598 41022 29650
rect 41074 29598 41076 29650
rect 40964 29596 41076 29598
rect 40908 29558 40964 29596
rect 41020 29586 41076 29596
rect 40572 29362 40628 29372
rect 40460 28642 40516 29260
rect 40460 28590 40462 28642
rect 40514 28590 40516 28642
rect 40460 28578 40516 28590
rect 40796 25732 40852 25742
rect 40796 25638 40852 25676
rect 40124 23938 40404 23940
rect 40124 23886 40126 23938
rect 40178 23886 40404 23938
rect 40124 23884 40404 23886
rect 40460 23938 40516 23950
rect 40460 23886 40462 23938
rect 40514 23886 40516 23938
rect 40124 23874 40180 23884
rect 40124 23156 40180 23166
rect 40460 23156 40516 23886
rect 40180 23100 40516 23156
rect 40124 23062 40180 23100
rect 40012 22372 40068 22428
rect 41020 22484 41076 22494
rect 41020 22390 41076 22428
rect 39788 22370 40068 22372
rect 39788 22318 40014 22370
rect 40066 22318 40068 22370
rect 39788 22316 40068 22318
rect 39564 21812 39620 21822
rect 39228 21810 39620 21812
rect 39228 21758 39566 21810
rect 39618 21758 39620 21810
rect 39228 21756 39620 21758
rect 38444 21718 38500 21756
rect 39564 21746 39620 21756
rect 38668 21588 38724 21598
rect 38668 21494 38724 21532
rect 39788 21588 39844 22316
rect 40012 22306 40068 22316
rect 39844 21532 40068 21588
rect 39788 21494 39844 21532
rect 39004 21364 39060 21374
rect 39004 20690 39060 21308
rect 40012 20914 40068 21532
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 40012 20850 40068 20862
rect 39004 20638 39006 20690
rect 39058 20638 39060 20690
rect 39004 20626 39060 20638
rect 38556 20244 38612 20254
rect 38556 20132 38836 20188
rect 38780 20020 38836 20132
rect 39116 20020 39172 20030
rect 38780 20018 39172 20020
rect 38780 19966 38782 20018
rect 38834 19966 39118 20018
rect 39170 19966 39172 20018
rect 38780 19964 39172 19966
rect 38780 19954 38836 19964
rect 39116 19954 39172 19964
rect 39004 19796 39060 19806
rect 39004 19122 39060 19740
rect 39004 19070 39006 19122
rect 39058 19070 39060 19122
rect 39004 19058 39060 19070
rect 39564 19572 39620 19582
rect 38668 18450 38724 18462
rect 38668 18398 38670 18450
rect 38722 18398 38724 18450
rect 38668 17668 38724 18398
rect 38780 18452 38836 18462
rect 38780 18338 38836 18396
rect 38780 18286 38782 18338
rect 38834 18286 38836 18338
rect 38780 18274 38836 18286
rect 38668 16996 38724 17612
rect 39004 17556 39060 17566
rect 39004 17462 39060 17500
rect 38668 16930 38724 16940
rect 39564 16994 39620 19516
rect 39900 18338 39956 18350
rect 39900 18286 39902 18338
rect 39954 18286 39956 18338
rect 39564 16942 39566 16994
rect 39618 16942 39620 16994
rect 39564 16930 39620 16942
rect 39788 17668 39844 17678
rect 39900 17668 39956 18286
rect 39844 17612 39956 17668
rect 41020 17668 41076 17678
rect 38892 16884 38948 16894
rect 38556 16772 38612 16782
rect 38220 16770 38612 16772
rect 38220 16718 38558 16770
rect 38610 16718 38612 16770
rect 38220 16716 38612 16718
rect 38556 16706 38612 16716
rect 37884 15934 37886 15986
rect 37938 15934 37940 15986
rect 37884 15922 37940 15934
rect 37436 15314 37492 15326
rect 37436 15262 37438 15314
rect 37490 15262 37492 15314
rect 37436 14084 37492 15262
rect 37660 14306 37716 14318
rect 37660 14254 37662 14306
rect 37714 14254 37716 14306
rect 37660 14196 37716 14254
rect 37660 14140 38388 14196
rect 37436 14028 38276 14084
rect 37324 13916 37828 13972
rect 37772 13858 37828 13916
rect 37772 13806 37774 13858
rect 37826 13806 37828 13858
rect 37772 13794 37828 13806
rect 37100 13346 37156 13356
rect 38108 13524 38164 13534
rect 37100 13076 37156 13086
rect 36988 13074 37156 13076
rect 36988 13022 37102 13074
rect 37154 13022 37156 13074
rect 36988 13020 37156 13022
rect 37100 13010 37156 13020
rect 36652 12002 36708 12012
rect 37100 12402 37156 12414
rect 37100 12350 37102 12402
rect 37154 12350 37156 12402
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 36540 11732 36596 11742
rect 36540 11506 36596 11676
rect 36540 11454 36542 11506
rect 36594 11454 36596 11506
rect 36540 11442 36596 11454
rect 36988 11732 37044 11742
rect 36988 11394 37044 11676
rect 37100 11618 37156 12350
rect 38108 12402 38164 13468
rect 38220 13076 38276 14028
rect 38332 13300 38388 14140
rect 38892 13634 38948 16828
rect 39676 15428 39732 15438
rect 38892 13582 38894 13634
rect 38946 13582 38948 13634
rect 38892 13570 38948 13582
rect 39452 15426 39732 15428
rect 39452 15374 39678 15426
rect 39730 15374 39732 15426
rect 39452 15372 39732 15374
rect 38332 13234 38388 13244
rect 39340 13412 39396 13422
rect 38332 13076 38388 13086
rect 38220 13074 38388 13076
rect 38220 13022 38334 13074
rect 38386 13022 38388 13074
rect 38220 13020 38388 13022
rect 38332 13010 38388 13020
rect 38108 12350 38110 12402
rect 38162 12350 38164 12402
rect 38108 12338 38164 12350
rect 39228 12964 39284 12974
rect 39228 12178 39284 12908
rect 39340 12850 39396 13356
rect 39340 12798 39342 12850
rect 39394 12798 39396 12850
rect 39340 12786 39396 12798
rect 39340 12404 39396 12414
rect 39452 12404 39508 15372
rect 39676 15362 39732 15372
rect 39788 13970 39844 17612
rect 41020 17574 41076 17612
rect 39900 17444 39956 17454
rect 39900 17350 39956 17388
rect 40124 16100 40180 16110
rect 39788 13918 39790 13970
rect 39842 13918 39844 13970
rect 39788 12964 39844 13918
rect 39788 12898 39844 12908
rect 39900 16098 40180 16100
rect 39900 16046 40126 16098
rect 40178 16046 40180 16098
rect 39900 16044 40180 16046
rect 39340 12402 39508 12404
rect 39340 12350 39342 12402
rect 39394 12350 39508 12402
rect 39340 12348 39508 12350
rect 39340 12338 39396 12348
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 37884 12068 37940 12078
rect 37100 11566 37102 11618
rect 37154 11566 37156 11618
rect 37100 11554 37156 11566
rect 37772 11954 37828 11966
rect 37772 11902 37774 11954
rect 37826 11902 37828 11954
rect 36988 11342 36990 11394
rect 37042 11342 37044 11394
rect 36988 11330 37044 11342
rect 34972 11282 35028 11294
rect 34972 11230 34974 11282
rect 35026 11230 35028 11282
rect 34972 11172 35028 11230
rect 34972 11106 35028 11116
rect 37772 10836 37828 11902
rect 37772 10770 37828 10780
rect 37884 10722 37940 12012
rect 39228 11844 39284 12126
rect 39228 11778 39284 11788
rect 38444 11732 38500 11742
rect 38444 11506 38500 11676
rect 38444 11454 38446 11506
rect 38498 11454 38500 11506
rect 38444 11442 38500 11454
rect 39900 11508 39956 16044
rect 40124 16034 40180 16044
rect 40572 16098 40628 16110
rect 40572 16046 40574 16098
rect 40626 16046 40628 16098
rect 40460 15092 40516 15102
rect 40460 14998 40516 15036
rect 39900 11442 39956 11452
rect 40012 14530 40068 14542
rect 40012 14478 40014 14530
rect 40066 14478 40068 14530
rect 37884 10670 37886 10722
rect 37938 10670 37940 10722
rect 37884 10658 37940 10670
rect 39116 10836 39172 10846
rect 28476 9998 28478 10050
rect 28530 9998 28532 10050
rect 28476 9986 28532 9998
rect 30044 9996 30212 10052
rect 30044 9938 30100 9996
rect 30044 9886 30046 9938
rect 30098 9886 30100 9938
rect 30044 9874 30100 9886
rect 28028 9762 28084 9772
rect 28588 9828 28644 9838
rect 28588 9734 28644 9772
rect 29484 9828 29540 9838
rect 29484 9734 29540 9772
rect 30492 9828 30548 9838
rect 30492 9734 30548 9772
rect 32060 9828 32116 10444
rect 34748 10434 34804 10444
rect 36876 10500 36932 10510
rect 36876 10406 36932 10444
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 32060 9762 32116 9772
rect 23212 9662 23214 9714
rect 23266 9662 23268 9714
rect 23212 9650 23268 9662
rect 39116 9714 39172 10780
rect 40012 9940 40068 14478
rect 40348 14532 40404 14542
rect 40572 14532 40628 16046
rect 41468 15092 41524 15102
rect 41524 15036 41748 15092
rect 41468 15026 41524 15036
rect 40348 14530 40628 14532
rect 40348 14478 40350 14530
rect 40402 14478 40628 14530
rect 40348 14476 40628 14478
rect 40348 13524 40404 14476
rect 40348 13458 40404 13468
rect 40348 13300 40404 13310
rect 40348 13074 40404 13244
rect 40348 13022 40350 13074
rect 40402 13022 40404 13074
rect 40348 13010 40404 13022
rect 40124 12964 40180 12974
rect 40124 12870 40180 12908
rect 40684 11508 40740 11518
rect 40684 11414 40740 11452
rect 41692 11282 41748 15036
rect 41692 11230 41694 11282
rect 41746 11230 41748 11282
rect 41692 11218 41748 11230
rect 40236 9940 40292 9950
rect 40012 9938 40292 9940
rect 40012 9886 40238 9938
rect 40290 9886 40292 9938
rect 40012 9884 40292 9886
rect 40236 9874 40292 9884
rect 39116 9662 39118 9714
rect 39170 9662 39172 9714
rect 39116 9650 39172 9662
rect 21980 9102 21982 9154
rect 22034 9102 22036 9154
rect 21980 9090 22036 9102
rect 20972 8878 20974 8930
rect 21026 8878 21028 8930
rect 20972 8866 21028 8878
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 17276 8094 17278 8146
rect 17330 8094 17332 8146
rect 17276 8082 17332 8094
rect 18396 8372 18564 8428
rect 19516 8372 19684 8428
rect 18396 8146 18452 8372
rect 19516 8370 19572 8372
rect 19516 8318 19518 8370
rect 19570 8318 19572 8370
rect 19516 8306 19572 8318
rect 18396 8094 18398 8146
rect 18450 8094 18452 8146
rect 18396 8082 18452 8094
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 14252 7588 14308 7598
rect 14252 7494 14308 7532
rect 13244 7310 13246 7362
rect 13298 7310 13300 7362
rect 13244 7298 13300 7310
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 4284 6580 4340 6590
rect 3836 5236 3892 5246
rect 3836 5122 3892 5180
rect 3836 5070 3838 5122
rect 3890 5070 3892 5122
rect 3836 5058 3892 5070
rect 3612 4958 3614 5010
rect 3666 4958 3668 5010
rect 3612 4946 3668 4958
rect 3724 5012 3780 5022
rect 3612 4564 3668 4574
rect 3612 4470 3668 4508
rect 3388 3390 3390 3442
rect 3442 3390 3444 3442
rect 3388 3378 3444 3390
rect 3724 3442 3780 4956
rect 4284 5010 4340 6524
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 4508 5124 4564 5134
rect 6972 5124 7028 5134
rect 4508 5030 4564 5068
rect 6636 5122 7028 5124
rect 6636 5070 6974 5122
rect 7026 5070 7028 5122
rect 6636 5068 7028 5070
rect 4284 4958 4286 5010
rect 4338 4958 4340 5010
rect 4284 4946 4340 4958
rect 4844 4452 4900 4462
rect 4844 4358 4900 4396
rect 3724 3390 3726 3442
rect 3778 3390 3780 3442
rect 3724 3378 3780 3390
rect 3836 4338 3892 4350
rect 3836 4286 3838 4338
rect 3890 4286 3892 4338
rect 3836 4228 3892 4286
rect 4396 4228 4452 4238
rect 3836 4226 4452 4228
rect 3836 4174 4398 4226
rect 4450 4174 4452 4226
rect 3836 4172 4452 4174
rect 3836 2100 3892 4172
rect 4396 4162 4452 4172
rect 5292 4226 5348 4238
rect 5292 4174 5294 4226
rect 5346 4174 5348 4226
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 3948 3554 4004 3566
rect 3948 3502 3950 3554
rect 4002 3502 4004 3554
rect 3948 3444 4004 3502
rect 5292 3556 5348 4174
rect 5740 4228 5796 4238
rect 5740 4134 5796 4172
rect 5292 3490 5348 3500
rect 4508 3444 4564 3454
rect 3948 3442 4564 3444
rect 3948 3390 4510 3442
rect 4562 3390 4564 3442
rect 3948 3388 4564 3390
rect 3948 2772 4004 3388
rect 4508 3378 4564 3388
rect 4956 3444 5012 3454
rect 4956 3350 5012 3388
rect 6076 3444 6132 3454
rect 6300 3444 6356 3454
rect 6076 3442 6356 3444
rect 6076 3390 6078 3442
rect 6130 3390 6302 3442
rect 6354 3390 6356 3442
rect 6076 3388 6356 3390
rect 3948 2706 4004 2716
rect 3836 2034 3892 2044
rect 6076 800 6132 3388
rect 6300 3378 6356 3388
rect 6636 3442 6692 5068
rect 6972 5058 7028 5068
rect 10444 5124 10500 5134
rect 10444 5122 10612 5124
rect 10444 5070 10446 5122
rect 10498 5070 10612 5122
rect 10444 5068 10612 5070
rect 10444 5058 10500 5068
rect 7308 4900 7364 4910
rect 7308 4898 7588 4900
rect 7308 4846 7310 4898
rect 7362 4846 7588 4898
rect 7308 4844 7588 4846
rect 7308 4834 7364 4844
rect 7532 3554 7588 4844
rect 7980 3668 8036 3678
rect 7532 3502 7534 3554
rect 7586 3502 7588 3554
rect 7532 3490 7588 3502
rect 7644 3666 8036 3668
rect 7644 3614 7982 3666
rect 8034 3614 8036 3666
rect 7644 3612 8036 3614
rect 6636 3390 6638 3442
rect 6690 3390 6692 3442
rect 6636 3378 6692 3390
rect 6972 3332 7028 3342
rect 6748 3330 7028 3332
rect 6748 3278 6974 3330
rect 7026 3278 7028 3330
rect 6748 3276 7028 3278
rect 6748 800 6804 3276
rect 6972 3266 7028 3276
rect 7644 980 7700 3612
rect 7980 3602 8036 3612
rect 10108 3444 10164 3454
rect 10332 3444 10388 3454
rect 10108 3442 10388 3444
rect 10108 3390 10110 3442
rect 10162 3390 10334 3442
rect 10386 3390 10388 3442
rect 10108 3388 10388 3390
rect 10556 3444 10612 5068
rect 10668 4900 10724 4910
rect 10668 4898 11060 4900
rect 10668 4846 10670 4898
rect 10722 4846 11060 4898
rect 10668 4844 11060 4846
rect 10668 4834 10724 4844
rect 11004 3554 11060 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 11452 3668 11508 3678
rect 11004 3502 11006 3554
rect 11058 3502 11060 3554
rect 11004 3490 11060 3502
rect 11116 3666 11508 3668
rect 11116 3614 11454 3666
rect 11506 3614 11508 3666
rect 11116 3612 11508 3614
rect 10668 3444 10724 3454
rect 10556 3442 10724 3444
rect 10556 3390 10670 3442
rect 10722 3390 10724 3442
rect 10556 3388 10724 3390
rect 7420 924 7700 980
rect 8092 3332 8148 3342
rect 7420 800 7476 924
rect 8092 800 8148 3276
rect 9324 3332 9380 3342
rect 9324 3238 9380 3276
rect 10108 800 10164 3388
rect 10332 3378 10388 3388
rect 10668 3378 10724 3388
rect 11116 980 11172 3612
rect 11452 3602 11508 3612
rect 13132 3330 13188 3342
rect 13132 3278 13134 3330
rect 13186 3278 13188 3330
rect 10780 924 11172 980
rect 12124 1762 12180 1774
rect 12124 1710 12126 1762
rect 12178 1710 12180 1762
rect 10780 800 10836 924
rect 12124 800 12180 1710
rect 13132 1762 13188 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 13132 1710 13134 1762
rect 13186 1710 13188 1762
rect 13132 1698 13188 1710
rect 2940 18 2996 28
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
<< via2 >>
rect 28 40124 84 40180
rect 1932 43036 1988 43092
rect 1820 40626 1876 40628
rect 1820 40574 1822 40626
rect 1822 40574 1874 40626
rect 1874 40574 1876 40626
rect 1820 40572 1876 40574
rect 1372 39004 1428 39060
rect 2044 40236 2100 40292
rect 1932 38780 1988 38836
rect 1596 37660 1652 37716
rect 812 36764 868 36820
rect 1596 36428 1652 36484
rect 2156 39058 2212 39060
rect 2156 39006 2158 39058
rect 2158 39006 2210 39058
rect 2210 39006 2212 39058
rect 2156 39004 2212 39006
rect 1708 35980 1764 36036
rect 1932 36316 1988 36372
rect 3388 42364 3444 42420
rect 3388 41020 3444 41076
rect 3276 40402 3332 40404
rect 3276 40350 3278 40402
rect 3278 40350 3330 40402
rect 3330 40350 3332 40402
rect 3276 40348 3332 40350
rect 3276 39394 3332 39396
rect 3276 39342 3278 39394
rect 3278 39342 3330 39394
rect 3330 39342 3332 39394
rect 3276 39340 3332 39342
rect 2940 38946 2996 38948
rect 2940 38894 2942 38946
rect 2942 38894 2994 38946
rect 2994 38894 2996 38946
rect 2940 38892 2996 38894
rect 3724 41692 3780 41748
rect 4284 43148 4340 43204
rect 4284 41132 4340 41188
rect 4732 40572 4788 40628
rect 4956 40460 5012 40516
rect 5740 40460 5796 40516
rect 5628 40348 5684 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3948 39676 4004 39732
rect 3500 38332 3556 38388
rect 2716 37772 2772 37828
rect 2380 36764 2436 36820
rect 2380 36370 2436 36372
rect 2380 36318 2382 36370
rect 2382 36318 2434 36370
rect 2434 36318 2436 36370
rect 2380 36316 2436 36318
rect 2380 35980 2436 36036
rect 1708 34972 1764 35028
rect 2156 35196 2212 35252
rect 2044 34300 2100 34356
rect 1708 33628 1764 33684
rect 2044 33234 2100 33236
rect 2044 33182 2046 33234
rect 2046 33182 2098 33234
rect 2098 33182 2100 33234
rect 2044 33180 2100 33182
rect 1708 32956 1764 33012
rect 2492 32956 2548 33012
rect 1708 32284 1764 32340
rect 2940 37490 2996 37492
rect 2940 37438 2942 37490
rect 2942 37438 2994 37490
rect 2994 37438 2996 37490
rect 2940 37436 2996 37438
rect 2716 37100 2772 37156
rect 3276 37826 3332 37828
rect 3276 37774 3278 37826
rect 3278 37774 3330 37826
rect 3330 37774 3332 37826
rect 3276 37772 3332 37774
rect 2828 36652 2884 36708
rect 3276 35980 3332 36036
rect 3388 36316 3444 36372
rect 3276 35810 3332 35812
rect 3276 35758 3278 35810
rect 3278 35758 3330 35810
rect 3330 35758 3332 35810
rect 3276 35756 3332 35758
rect 3164 34860 3220 34916
rect 2828 34636 2884 34692
rect 1932 31612 1988 31668
rect 2044 31052 2100 31108
rect 2044 30828 2100 30884
rect 2716 30716 2772 30772
rect 2380 30268 2436 30324
rect 1708 29596 1764 29652
rect 2044 29820 2100 29876
rect 1708 28924 1764 28980
rect 2044 29260 2100 29316
rect 2492 28924 2548 28980
rect 1708 28252 1764 28308
rect 2492 28252 2548 28308
rect 2044 27970 2100 27972
rect 2044 27918 2046 27970
rect 2046 27918 2098 27970
rect 2098 27918 2100 27970
rect 2044 27916 2100 27918
rect 1708 27580 1764 27636
rect 2492 27580 2548 27636
rect 3276 35084 3332 35140
rect 2940 30994 2996 30996
rect 2940 30942 2942 30994
rect 2942 30942 2994 30994
rect 2994 30942 2996 30994
rect 2940 30940 2996 30942
rect 2268 26908 2324 26964
rect 2156 26236 2212 26292
rect 1820 26178 1876 26180
rect 1820 26126 1822 26178
rect 1822 26126 1874 26178
rect 1874 26126 1876 26178
rect 1820 26124 1876 26126
rect 3164 30716 3220 30772
rect 3276 32508 3332 32564
rect 3164 30268 3220 30324
rect 3612 37266 3668 37268
rect 3612 37214 3614 37266
rect 3614 37214 3666 37266
rect 3666 37214 3668 37266
rect 3612 37212 3668 37214
rect 3612 36988 3668 37044
rect 5740 39004 5796 39060
rect 4844 38946 4900 38948
rect 4844 38894 4846 38946
rect 4846 38894 4898 38946
rect 4898 38894 4900 38946
rect 4844 38892 4900 38894
rect 4172 38332 4228 38388
rect 4060 38108 4116 38164
rect 3948 36876 4004 36932
rect 4060 36370 4116 36372
rect 4060 36318 4062 36370
rect 4062 36318 4114 36370
rect 4114 36318 4116 36370
rect 4060 36316 4116 36318
rect 5068 38834 5124 38836
rect 5068 38782 5070 38834
rect 5070 38782 5122 38834
rect 5122 38782 5124 38834
rect 5068 38780 5124 38782
rect 4956 38668 5012 38724
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4396 37436 4452 37492
rect 4732 37938 4788 37940
rect 4732 37886 4734 37938
rect 4734 37886 4786 37938
rect 4786 37886 4788 37938
rect 4732 37884 4788 37886
rect 4844 37436 4900 37492
rect 4172 35196 4228 35252
rect 3948 35084 4004 35140
rect 3724 32508 3780 32564
rect 3612 29596 3668 29652
rect 1820 25564 1876 25620
rect 3276 26124 3332 26180
rect 2156 24892 2212 24948
rect 2940 24722 2996 24724
rect 2940 24670 2942 24722
rect 2942 24670 2994 24722
rect 2994 24670 2996 24722
rect 2940 24668 2996 24670
rect 1932 24220 1988 24276
rect 2044 23826 2100 23828
rect 2044 23774 2046 23826
rect 2046 23774 2098 23826
rect 2098 23774 2100 23826
rect 2044 23772 2100 23774
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4396 36482 4452 36484
rect 4396 36430 4398 36482
rect 4398 36430 4450 36482
rect 4450 36430 4452 36482
rect 4396 36428 4452 36430
rect 5516 38220 5572 38276
rect 5292 37884 5348 37940
rect 5628 37826 5684 37828
rect 5628 37774 5630 37826
rect 5630 37774 5682 37826
rect 5682 37774 5684 37826
rect 5628 37772 5684 37774
rect 5740 37436 5796 37492
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4956 32620 5012 32676
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5740 32674 5796 32676
rect 5740 32622 5742 32674
rect 5742 32622 5794 32674
rect 5794 32622 5796 32674
rect 5740 32620 5796 32622
rect 6188 38946 6244 38948
rect 6188 38894 6190 38946
rect 6190 38894 6242 38946
rect 6242 38894 6244 38946
rect 6188 38892 6244 38894
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5740 30156 5796 30212
rect 5516 29260 5572 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 5964 30940 6020 30996
rect 6188 31388 6244 31444
rect 6076 30828 6132 30884
rect 5852 28924 5908 28980
rect 6412 31052 6468 31108
rect 6860 39340 6916 39396
rect 6636 38108 6692 38164
rect 7308 39116 7364 39172
rect 6636 37100 6692 37156
rect 8428 40124 8484 40180
rect 7308 38556 7364 38612
rect 7868 39116 7924 39172
rect 8428 39004 8484 39060
rect 8316 38946 8372 38948
rect 8316 38894 8318 38946
rect 8318 38894 8370 38946
rect 8370 38894 8372 38946
rect 8316 38892 8372 38894
rect 8092 38834 8148 38836
rect 8092 38782 8094 38834
rect 8094 38782 8146 38834
rect 8146 38782 8148 38834
rect 8092 38780 8148 38782
rect 9548 41132 9604 41188
rect 9436 40236 9492 40292
rect 7644 38668 7700 38724
rect 8316 38220 8372 38276
rect 7980 37996 8036 38052
rect 7644 37938 7700 37940
rect 7644 37886 7646 37938
rect 7646 37886 7698 37938
rect 7698 37886 7700 37938
rect 7644 37884 7700 37886
rect 9324 38444 9380 38500
rect 9100 38332 9156 38388
rect 8652 37826 8708 37828
rect 8652 37774 8654 37826
rect 8654 37774 8706 37826
rect 8706 37774 8708 37826
rect 8652 37772 8708 37774
rect 8204 37100 8260 37156
rect 8988 37154 9044 37156
rect 8988 37102 8990 37154
rect 8990 37102 9042 37154
rect 9042 37102 9044 37154
rect 8988 37100 9044 37102
rect 9996 39340 10052 39396
rect 9660 39058 9716 39060
rect 9660 39006 9662 39058
rect 9662 39006 9714 39058
rect 9714 39006 9716 39058
rect 9660 39004 9716 39006
rect 9772 38108 9828 38164
rect 10220 38722 10276 38724
rect 10220 38670 10222 38722
rect 10222 38670 10274 38722
rect 10274 38670 10276 38722
rect 10220 38668 10276 38670
rect 10556 40236 10612 40292
rect 10668 39116 10724 39172
rect 16156 39788 16212 39844
rect 16828 39788 16884 39844
rect 16380 39394 16436 39396
rect 16380 39342 16382 39394
rect 16382 39342 16434 39394
rect 16434 39342 16436 39394
rect 16380 39340 16436 39342
rect 18172 40572 18228 40628
rect 17052 39116 17108 39172
rect 15148 38444 15204 38500
rect 19180 40626 19236 40628
rect 19180 40574 19182 40626
rect 19182 40574 19234 40626
rect 19234 40574 19236 40626
rect 19180 40572 19236 40574
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19852 40626 19908 40628
rect 19852 40574 19854 40626
rect 19854 40574 19906 40626
rect 19906 40574 19908 40626
rect 19852 40572 19908 40574
rect 20972 40572 21028 40628
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19068 38332 19124 38388
rect 20748 38220 20804 38276
rect 21756 38108 21812 38164
rect 22876 39730 22932 39732
rect 22876 39678 22878 39730
rect 22878 39678 22930 39730
rect 22930 39678 22932 39730
rect 22876 39676 22932 39678
rect 23996 39676 24052 39732
rect 22428 37996 22484 38052
rect 25116 40236 25172 40292
rect 24556 38892 24612 38948
rect 23772 37884 23828 37940
rect 18508 37772 18564 37828
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 26572 40290 26628 40292
rect 26572 40238 26574 40290
rect 26574 40238 26626 40290
rect 26626 40238 26628 40290
rect 26572 40236 26628 40238
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 26460 38668 26516 38724
rect 26124 38556 26180 38612
rect 25788 37100 25844 37156
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 9548 35756 9604 35812
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 7196 33180 7252 33236
rect 8092 31836 8148 31892
rect 6860 30828 6916 30884
rect 7756 30210 7812 30212
rect 7756 30158 7758 30210
rect 7758 30158 7810 30210
rect 7810 30158 7812 30210
rect 7756 30156 7812 30158
rect 14028 33404 14084 33460
rect 8764 31388 8820 31444
rect 8988 31218 9044 31220
rect 8988 31166 8990 31218
rect 8990 31166 9042 31218
rect 9042 31166 9044 31218
rect 8988 31164 9044 31166
rect 8316 30828 8372 30884
rect 6524 29820 6580 29876
rect 8652 30156 8708 30212
rect 8764 30044 8820 30100
rect 6972 28924 7028 28980
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6076 27132 6132 27188
rect 6860 27186 6916 27188
rect 6860 27134 6862 27186
rect 6862 27134 6914 27186
rect 6914 27134 6916 27186
rect 6860 27132 6916 27134
rect 6188 27020 6244 27076
rect 5404 26908 5460 26964
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 9660 31218 9716 31220
rect 9660 31166 9662 31218
rect 9662 31166 9714 31218
rect 9714 31166 9716 31218
rect 9660 31164 9716 31166
rect 9100 29372 9156 29428
rect 9660 29650 9716 29652
rect 9660 29598 9662 29650
rect 9662 29598 9714 29650
rect 9714 29598 9716 29650
rect 9660 29596 9716 29598
rect 9772 30492 9828 30548
rect 10108 30882 10164 30884
rect 10108 30830 10110 30882
rect 10110 30830 10162 30882
rect 10162 30830 10164 30882
rect 10108 30828 10164 30830
rect 9884 29372 9940 29428
rect 10332 30156 10388 30212
rect 11228 31164 11284 31220
rect 11676 31164 11732 31220
rect 10892 30492 10948 30548
rect 11004 30156 11060 30212
rect 11676 30210 11732 30212
rect 11676 30158 11678 30210
rect 11678 30158 11730 30210
rect 11730 30158 11732 30210
rect 11676 30156 11732 30158
rect 12572 30210 12628 30212
rect 12572 30158 12574 30210
rect 12574 30158 12626 30210
rect 12626 30158 12628 30210
rect 12572 30156 12628 30158
rect 11452 30098 11508 30100
rect 11452 30046 11454 30098
rect 11454 30046 11506 30098
rect 11506 30046 11508 30098
rect 11452 30044 11508 30046
rect 7868 26962 7924 26964
rect 7868 26910 7870 26962
rect 7870 26910 7922 26962
rect 7922 26910 7924 26962
rect 7868 26908 7924 26910
rect 7308 26796 7364 26852
rect 8652 27020 8708 27076
rect 8876 26908 8932 26964
rect 9884 28364 9940 28420
rect 9212 26850 9268 26852
rect 9212 26798 9214 26850
rect 9214 26798 9266 26850
rect 9266 26798 9268 26850
rect 9212 26796 9268 26798
rect 10668 29596 10724 29652
rect 12236 29596 12292 29652
rect 11228 28588 11284 28644
rect 11228 27020 11284 27076
rect 10108 26908 10164 26964
rect 13468 30210 13524 30212
rect 13468 30158 13470 30210
rect 13470 30158 13522 30210
rect 13522 30158 13524 30210
rect 13468 30156 13524 30158
rect 13132 30044 13188 30100
rect 12572 28700 12628 28756
rect 12236 27074 12292 27076
rect 12236 27022 12238 27074
rect 12238 27022 12290 27074
rect 12290 27022 12292 27074
rect 12236 27020 12292 27022
rect 14588 31164 14644 31220
rect 14364 30492 14420 30548
rect 13580 28700 13636 28756
rect 8316 26460 8372 26516
rect 8540 26684 8596 26740
rect 9772 26402 9828 26404
rect 9772 26350 9774 26402
rect 9774 26350 9826 26402
rect 9826 26350 9828 26402
rect 9772 26348 9828 26350
rect 10556 26796 10612 26852
rect 15148 33458 15204 33460
rect 15148 33406 15150 33458
rect 15150 33406 15202 33458
rect 15202 33406 15204 33458
rect 15148 33404 15204 33406
rect 15036 31836 15092 31892
rect 15596 31218 15652 31220
rect 15596 31166 15598 31218
rect 15598 31166 15650 31218
rect 15650 31166 15652 31218
rect 15596 31164 15652 31166
rect 15932 30492 15988 30548
rect 15708 30156 15764 30212
rect 14924 30044 14980 30100
rect 14140 28700 14196 28756
rect 13916 28028 13972 28084
rect 14924 28700 14980 28756
rect 14476 27916 14532 27972
rect 14924 27074 14980 27076
rect 14924 27022 14926 27074
rect 14926 27022 14978 27074
rect 14978 27022 14980 27074
rect 14924 27020 14980 27022
rect 15596 26572 15652 26628
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23772 4340 23828
rect 4732 23772 4788 23828
rect 1708 23548 1764 23604
rect 2492 23548 2548 23604
rect 2044 23436 2100 23492
rect 1708 22876 1764 22932
rect 1708 22428 1764 22484
rect 6188 23772 6244 23828
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5292 22764 5348 22820
rect 2492 22482 2548 22484
rect 2492 22430 2494 22482
rect 2494 22430 2546 22482
rect 2546 22430 2548 22482
rect 2492 22428 2548 22430
rect 4844 22204 4900 22260
rect 2380 21644 2436 21700
rect 3500 21644 3556 21700
rect 1820 21586 1876 21588
rect 1820 21534 1822 21586
rect 1822 21534 1874 21586
rect 1874 21534 1876 21586
rect 1820 21532 1876 21534
rect 1708 20860 1764 20916
rect 1596 20636 1652 20692
rect 2716 20690 2772 20692
rect 2716 20638 2718 20690
rect 2718 20638 2770 20690
rect 2770 20638 2772 20690
rect 2716 20636 2772 20638
rect 3388 20300 3444 20356
rect 1596 14364 1652 14420
rect 2380 17666 2436 17668
rect 2380 17614 2382 17666
rect 2382 17614 2434 17666
rect 2434 17614 2436 17666
rect 2380 17612 2436 17614
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 9548 24780 9604 24836
rect 8092 23660 8148 23716
rect 7532 22764 7588 22820
rect 7084 22258 7140 22260
rect 7084 22206 7086 22258
rect 7086 22206 7138 22258
rect 7138 22206 7140 22258
rect 7084 22204 7140 22206
rect 6972 21980 7028 22036
rect 8092 22482 8148 22484
rect 8092 22430 8094 22482
rect 8094 22430 8146 22482
rect 8146 22430 8148 22482
rect 8092 22428 8148 22430
rect 8204 22092 8260 22148
rect 9436 23660 9492 23716
rect 10444 24834 10500 24836
rect 10444 24782 10446 24834
rect 10446 24782 10498 24834
rect 10498 24782 10500 24834
rect 10444 24780 10500 24782
rect 15484 25564 15540 25620
rect 10892 24780 10948 24836
rect 11228 23548 11284 23604
rect 11900 23826 11956 23828
rect 11900 23774 11902 23826
rect 11902 23774 11954 23826
rect 11954 23774 11956 23826
rect 11900 23772 11956 23774
rect 12348 23826 12404 23828
rect 12348 23774 12350 23826
rect 12350 23774 12402 23826
rect 12402 23774 12404 23826
rect 12348 23772 12404 23774
rect 16156 31778 16212 31780
rect 16156 31726 16158 31778
rect 16158 31726 16210 31778
rect 16210 31726 16212 31778
rect 16156 31724 16212 31726
rect 17276 33068 17332 33124
rect 18396 31554 18452 31556
rect 18396 31502 18398 31554
rect 18398 31502 18450 31554
rect 18450 31502 18452 31554
rect 18396 31500 18452 31502
rect 17836 31052 17892 31108
rect 17388 30210 17444 30212
rect 17388 30158 17390 30210
rect 17390 30158 17442 30210
rect 17442 30158 17444 30210
rect 17388 30156 17444 30158
rect 16156 29484 16212 29540
rect 16716 29932 16772 29988
rect 16156 27804 16212 27860
rect 17500 29314 17556 29316
rect 17500 29262 17502 29314
rect 17502 29262 17554 29314
rect 17554 29262 17556 29314
rect 17500 29260 17556 29262
rect 16828 28364 16884 28420
rect 17948 29314 18004 29316
rect 17948 29262 17950 29314
rect 17950 29262 18002 29314
rect 18002 29262 18004 29314
rect 17948 29260 18004 29262
rect 18060 28700 18116 28756
rect 16604 27804 16660 27860
rect 16156 27074 16212 27076
rect 16156 27022 16158 27074
rect 16158 27022 16210 27074
rect 16210 27022 16212 27074
rect 16156 27020 16212 27022
rect 17164 26908 17220 26964
rect 16268 25564 16324 25620
rect 16940 26402 16996 26404
rect 16940 26350 16942 26402
rect 16942 26350 16994 26402
rect 16994 26350 16996 26402
rect 16940 26348 16996 26350
rect 16380 24892 16436 24948
rect 16604 25564 16660 25620
rect 15820 24834 15876 24836
rect 15820 24782 15822 24834
rect 15822 24782 15874 24834
rect 15874 24782 15876 24834
rect 15820 24780 15876 24782
rect 12796 23660 12852 23716
rect 13356 23548 13412 23604
rect 12572 23266 12628 23268
rect 12572 23214 12574 23266
rect 12574 23214 12626 23266
rect 12626 23214 12628 23266
rect 12572 23212 12628 23214
rect 9548 21868 9604 21924
rect 10668 22092 10724 22148
rect 10668 21868 10724 21924
rect 7980 21644 8036 21700
rect 5628 21586 5684 21588
rect 5628 21534 5630 21586
rect 5630 21534 5682 21586
rect 5682 21534 5684 21586
rect 5628 21532 5684 21534
rect 6748 21532 6804 21588
rect 4844 20748 4900 20804
rect 4060 20300 4116 20356
rect 7980 21474 8036 21476
rect 7980 21422 7982 21474
rect 7982 21422 8034 21474
rect 8034 21422 8036 21474
rect 7980 21420 8036 21422
rect 6188 20300 6244 20356
rect 3836 18844 3892 18900
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4060 19346 4116 19348
rect 4060 19294 4062 19346
rect 4062 19294 4114 19346
rect 4114 19294 4116 19346
rect 4060 19292 4116 19294
rect 7756 20076 7812 20132
rect 7084 18956 7140 19012
rect 6076 18844 6132 18900
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 3388 17666 3444 17668
rect 3388 17614 3390 17666
rect 3390 17614 3442 17666
rect 3442 17614 3444 17666
rect 3388 17612 3444 17614
rect 4732 17666 4788 17668
rect 4732 17614 4734 17666
rect 4734 17614 4786 17666
rect 4786 17614 4788 17666
rect 4732 17612 4788 17614
rect 3052 15986 3108 15988
rect 3052 15934 3054 15986
rect 3054 15934 3106 15986
rect 3106 15934 3108 15986
rect 3052 15932 3108 15934
rect 2716 14418 2772 14420
rect 2716 14366 2718 14418
rect 2718 14366 2770 14418
rect 2770 14366 2772 14418
rect 2716 14364 2772 14366
rect 4732 16716 4788 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5628 17106 5684 17108
rect 5628 17054 5630 17106
rect 5630 17054 5682 17106
rect 5682 17054 5684 17106
rect 5628 17052 5684 17054
rect 7532 18450 7588 18452
rect 7532 18398 7534 18450
rect 7534 18398 7586 18450
rect 7586 18398 7588 18450
rect 7532 18396 7588 18398
rect 9660 20076 9716 20132
rect 8092 19292 8148 19348
rect 8764 19010 8820 19012
rect 8764 18958 8766 19010
rect 8766 18958 8818 19010
rect 8818 18958 8820 19010
rect 8764 18956 8820 18958
rect 8988 18284 9044 18340
rect 8876 18172 8932 18228
rect 8092 17778 8148 17780
rect 8092 17726 8094 17778
rect 8094 17726 8146 17778
rect 8146 17726 8148 17778
rect 8092 17724 8148 17726
rect 7532 17612 7588 17668
rect 6300 17052 6356 17108
rect 4956 16380 5012 16436
rect 3948 16044 4004 16100
rect 5516 15986 5572 15988
rect 5516 15934 5518 15986
rect 5518 15934 5570 15986
rect 5570 15934 5572 15986
rect 5516 15932 5572 15934
rect 4060 15260 4116 15316
rect 5068 15314 5124 15316
rect 5068 15262 5070 15314
rect 5070 15262 5122 15314
rect 5122 15262 5124 15314
rect 5068 15260 5124 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3388 13692 3444 13748
rect 4620 13746 4676 13748
rect 4620 13694 4622 13746
rect 4622 13694 4674 13746
rect 4674 13694 4676 13746
rect 4620 13692 4676 13694
rect 4172 13468 4228 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 10332 17836 10388 17892
rect 9884 17666 9940 17668
rect 9884 17614 9886 17666
rect 9886 17614 9938 17666
rect 9938 17614 9940 17666
rect 9884 17612 9940 17614
rect 9548 16940 9604 16996
rect 7532 16770 7588 16772
rect 7532 16718 7534 16770
rect 7534 16718 7586 16770
rect 7586 16718 7588 16770
rect 7532 16716 7588 16718
rect 7420 16380 7476 16436
rect 8540 16098 8596 16100
rect 8540 16046 8542 16098
rect 8542 16046 8594 16098
rect 8594 16046 8596 16098
rect 8540 16044 8596 16046
rect 11788 22204 11844 22260
rect 12460 22204 12516 22260
rect 13020 22146 13076 22148
rect 13020 22094 13022 22146
rect 13022 22094 13074 22146
rect 13074 22094 13076 22146
rect 13020 22092 13076 22094
rect 13804 22428 13860 22484
rect 14252 22428 14308 22484
rect 14588 23212 14644 23268
rect 14924 22876 14980 22932
rect 13916 22258 13972 22260
rect 13916 22206 13918 22258
rect 13918 22206 13970 22258
rect 13970 22206 13972 22258
rect 13916 22204 13972 22206
rect 14252 22258 14308 22260
rect 14252 22206 14254 22258
rect 14254 22206 14306 22258
rect 14306 22206 14308 22258
rect 14252 22204 14308 22206
rect 14924 22204 14980 22260
rect 12460 21586 12516 21588
rect 12460 21534 12462 21586
rect 12462 21534 12514 21586
rect 12514 21534 12516 21586
rect 12460 21532 12516 21534
rect 13580 20188 13636 20244
rect 11340 18396 11396 18452
rect 10556 16994 10612 16996
rect 10556 16942 10558 16994
rect 10558 16942 10610 16994
rect 10610 16942 10612 16994
rect 10556 16940 10612 16942
rect 11900 18284 11956 18340
rect 12572 18226 12628 18228
rect 12572 18174 12574 18226
rect 12574 18174 12626 18226
rect 12626 18174 12628 18226
rect 12572 18172 12628 18174
rect 13020 17890 13076 17892
rect 13020 17838 13022 17890
rect 13022 17838 13074 17890
rect 13074 17838 13076 17890
rect 13020 17836 13076 17838
rect 13244 17836 13300 17892
rect 12796 16940 12852 16996
rect 13580 16940 13636 16996
rect 12460 16268 12516 16324
rect 13580 16322 13636 16324
rect 13580 16270 13582 16322
rect 13582 16270 13634 16322
rect 13634 16270 13636 16322
rect 13580 16268 13636 16270
rect 6412 14588 6468 14644
rect 8540 14588 8596 14644
rect 13244 15538 13300 15540
rect 13244 15486 13246 15538
rect 13246 15486 13298 15538
rect 13298 15486 13300 15538
rect 13244 15484 13300 15486
rect 9548 14588 9604 14644
rect 10108 14418 10164 14420
rect 10108 14366 10110 14418
rect 10110 14366 10162 14418
rect 10162 14366 10164 14418
rect 10108 14364 10164 14366
rect 6076 13468 6132 13524
rect 9324 13132 9380 13188
rect 6972 12962 7028 12964
rect 6972 12910 6974 12962
rect 6974 12910 7026 12962
rect 7026 12910 7028 12962
rect 6972 12908 7028 12910
rect 8540 12908 8596 12964
rect 6860 12738 6916 12740
rect 6860 12686 6862 12738
rect 6862 12686 6914 12738
rect 6914 12686 6916 12738
rect 6860 12684 6916 12686
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 6076 11452 6132 11508
rect 7756 12738 7812 12740
rect 7756 12686 7758 12738
rect 7758 12686 7810 12738
rect 7810 12686 7812 12738
rect 7756 12684 7812 12686
rect 7644 11506 7700 11508
rect 7644 11454 7646 11506
rect 7646 11454 7698 11506
rect 7698 11454 7700 11506
rect 7644 11452 7700 11454
rect 7196 11228 7252 11284
rect 8652 11282 8708 11284
rect 8652 11230 8654 11282
rect 8654 11230 8706 11282
rect 8706 11230 8708 11282
rect 8652 11228 8708 11230
rect 9884 12908 9940 12964
rect 9772 12684 9828 12740
rect 9100 10668 9156 10724
rect 10444 14588 10500 14644
rect 12348 14418 12404 14420
rect 12348 14366 12350 14418
rect 12350 14366 12402 14418
rect 12402 14366 12404 14418
rect 12348 14364 12404 14366
rect 13804 21308 13860 21364
rect 15372 23660 15428 23716
rect 15708 23436 15764 23492
rect 15932 22876 15988 22932
rect 16268 23212 16324 23268
rect 15260 22316 15316 22372
rect 15036 21420 15092 21476
rect 15260 19906 15316 19908
rect 15260 19854 15262 19906
rect 15262 19854 15314 19906
rect 15314 19854 15316 19906
rect 15260 19852 15316 19854
rect 14028 17890 14084 17892
rect 14028 17838 14030 17890
rect 14030 17838 14082 17890
rect 14082 17838 14084 17890
rect 14028 17836 14084 17838
rect 13804 15484 13860 15540
rect 16492 23436 16548 23492
rect 24780 33516 24836 33572
rect 19740 33068 19796 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 23996 32956 24052 33012
rect 19180 32620 19236 32676
rect 20076 32674 20132 32676
rect 20076 32622 20078 32674
rect 20078 32622 20130 32674
rect 20130 32622 20132 32674
rect 20076 32620 20132 32622
rect 18732 31052 18788 31108
rect 19404 29932 19460 29988
rect 19404 29538 19460 29540
rect 19404 29486 19406 29538
rect 19406 29486 19458 29538
rect 19458 29486 19460 29538
rect 19404 29484 19460 29486
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20300 31554 20356 31556
rect 20300 31502 20302 31554
rect 20302 31502 20354 31554
rect 20354 31502 20356 31554
rect 20300 31500 20356 31502
rect 20188 29932 20244 29988
rect 20300 30044 20356 30100
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19516 29260 19572 29316
rect 21756 30828 21812 30884
rect 21532 30098 21588 30100
rect 21532 30046 21534 30098
rect 21534 30046 21586 30098
rect 21586 30046 21588 30098
rect 21532 30044 21588 30046
rect 21756 30044 21812 30100
rect 22204 30210 22260 30212
rect 22204 30158 22206 30210
rect 22206 30158 22258 30210
rect 22258 30158 22260 30210
rect 22204 30156 22260 30158
rect 19852 28754 19908 28756
rect 19852 28702 19854 28754
rect 19854 28702 19906 28754
rect 19906 28702 19908 28754
rect 19852 28700 19908 28702
rect 20524 28700 20580 28756
rect 19516 28642 19572 28644
rect 19516 28590 19518 28642
rect 19518 28590 19570 28642
rect 19570 28590 19572 28642
rect 19516 28588 19572 28590
rect 20636 28642 20692 28644
rect 20636 28590 20638 28642
rect 20638 28590 20690 28642
rect 20690 28590 20692 28642
rect 20636 28588 20692 28590
rect 20188 28530 20244 28532
rect 20188 28478 20190 28530
rect 20190 28478 20242 28530
rect 20242 28478 20244 28530
rect 20188 28476 20244 28478
rect 21196 29932 21252 29988
rect 21084 29036 21140 29092
rect 20860 28476 20916 28532
rect 24556 31724 24612 31780
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 23324 30156 23380 30212
rect 22764 29708 22820 29764
rect 26236 32956 26292 33012
rect 26348 33404 26404 33460
rect 26012 32450 26068 32452
rect 26012 32398 26014 32450
rect 26014 32398 26066 32450
rect 26066 32398 26068 32450
rect 26012 32396 26068 32398
rect 25676 31164 25732 31220
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 27244 33516 27300 33572
rect 27132 33458 27188 33460
rect 27132 33406 27134 33458
rect 27134 33406 27186 33458
rect 27186 33406 27188 33458
rect 27132 33404 27188 33406
rect 29596 33404 29652 33460
rect 24668 30044 24724 30100
rect 23548 29484 23604 29540
rect 24332 29538 24388 29540
rect 24332 29486 24334 29538
rect 24334 29486 24386 29538
rect 24386 29486 24388 29538
rect 24332 29484 24388 29486
rect 24108 29426 24164 29428
rect 24108 29374 24110 29426
rect 24110 29374 24162 29426
rect 24162 29374 24164 29426
rect 24108 29372 24164 29374
rect 22204 28700 22260 28756
rect 22316 29036 22372 29092
rect 24668 28700 24724 28756
rect 24780 30268 24836 30324
rect 24332 28642 24388 28644
rect 24332 28590 24334 28642
rect 24334 28590 24386 28642
rect 24386 28590 24388 28642
rect 24332 28588 24388 28590
rect 23548 28530 23604 28532
rect 23548 28478 23550 28530
rect 23550 28478 23602 28530
rect 23602 28478 23604 28530
rect 23548 28476 23604 28478
rect 21196 28364 21252 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18396 28028 18452 28084
rect 19740 27970 19796 27972
rect 19740 27918 19742 27970
rect 19742 27918 19794 27970
rect 19794 27918 19796 27970
rect 19740 27916 19796 27918
rect 20188 27858 20244 27860
rect 20188 27806 20190 27858
rect 20190 27806 20242 27858
rect 20242 27806 20244 27858
rect 20188 27804 20244 27806
rect 18284 26908 18340 26964
rect 25004 27916 25060 27972
rect 25788 30098 25844 30100
rect 25788 30046 25790 30098
rect 25790 30046 25842 30098
rect 25842 30046 25844 30098
rect 25788 30044 25844 30046
rect 25340 29314 25396 29316
rect 25340 29262 25342 29314
rect 25342 29262 25394 29314
rect 25394 29262 25396 29314
rect 25340 29260 25396 29262
rect 26124 29260 26180 29316
rect 26236 29708 26292 29764
rect 25340 28588 25396 28644
rect 18396 26684 18452 26740
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19404 26402 19460 26404
rect 19404 26350 19406 26402
rect 19406 26350 19458 26402
rect 19458 26350 19460 26402
rect 19404 26348 19460 26350
rect 20188 26402 20244 26404
rect 20188 26350 20190 26402
rect 20190 26350 20242 26402
rect 20242 26350 20244 26402
rect 20188 26348 20244 26350
rect 19628 26124 19684 26180
rect 17388 24892 17444 24948
rect 17052 23772 17108 23828
rect 17612 24780 17668 24836
rect 18284 24780 18340 24836
rect 18844 24834 18900 24836
rect 18844 24782 18846 24834
rect 18846 24782 18898 24834
rect 18898 24782 18900 24834
rect 18844 24780 18900 24782
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20076 24722 20132 24724
rect 20076 24670 20078 24722
rect 20078 24670 20130 24722
rect 20130 24670 20132 24722
rect 20076 24668 20132 24670
rect 17500 23436 17556 23492
rect 16716 22876 16772 22932
rect 16828 22428 16884 22484
rect 16940 21362 16996 21364
rect 16940 21310 16942 21362
rect 16942 21310 16994 21362
rect 16994 21310 16996 21362
rect 16940 21308 16996 21310
rect 17836 23436 17892 23492
rect 21084 26124 21140 26180
rect 20524 25618 20580 25620
rect 20524 25566 20526 25618
rect 20526 25566 20578 25618
rect 20578 25566 20580 25618
rect 20524 25564 20580 25566
rect 20412 24556 20468 24612
rect 21532 23996 21588 24052
rect 22204 25228 22260 25284
rect 18060 23212 18116 23268
rect 19180 23660 19236 23716
rect 17948 21308 18004 21364
rect 18732 22370 18788 22372
rect 18732 22318 18734 22370
rect 18734 22318 18786 22370
rect 18786 22318 18788 22370
rect 18732 22316 18788 22318
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18732 21474 18788 21476
rect 18732 21422 18734 21474
rect 18734 21422 18786 21474
rect 18786 21422 18788 21474
rect 18732 21420 18788 21422
rect 18284 20860 18340 20916
rect 19068 20914 19124 20916
rect 19068 20862 19070 20914
rect 19070 20862 19122 20914
rect 19122 20862 19124 20914
rect 19068 20860 19124 20862
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21420 23714 21476 23716
rect 21420 23662 21422 23714
rect 21422 23662 21474 23714
rect 21474 23662 21476 23714
rect 21420 23660 21476 23662
rect 21420 23378 21476 23380
rect 21420 23326 21422 23378
rect 21422 23326 21474 23378
rect 21474 23326 21476 23378
rect 21420 23324 21476 23326
rect 20972 23212 21028 23268
rect 20412 22370 20468 22372
rect 20412 22318 20414 22370
rect 20414 22318 20466 22370
rect 20466 22318 20468 22370
rect 20412 22316 20468 22318
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 17388 20188 17444 20244
rect 17164 19852 17220 19908
rect 15596 18450 15652 18452
rect 15596 18398 15598 18450
rect 15598 18398 15650 18450
rect 15650 18398 15652 18450
rect 15596 18396 15652 18398
rect 16604 16828 16660 16884
rect 16156 15820 16212 15876
rect 17164 19010 17220 19012
rect 17164 18958 17166 19010
rect 17166 18958 17218 19010
rect 17218 18958 17220 19010
rect 17164 18956 17220 18958
rect 19068 19740 19124 19796
rect 17836 18396 17892 18452
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 20076 19740 20132 19796
rect 21644 22370 21700 22372
rect 21644 22318 21646 22370
rect 21646 22318 21698 22370
rect 21698 22318 21700 22370
rect 21644 22316 21700 22318
rect 22428 26348 22484 26404
rect 23772 26402 23828 26404
rect 23772 26350 23774 26402
rect 23774 26350 23826 26402
rect 23826 26350 23828 26402
rect 23772 26348 23828 26350
rect 23436 26124 23492 26180
rect 22988 25506 23044 25508
rect 22988 25454 22990 25506
rect 22990 25454 23042 25506
rect 23042 25454 23044 25506
rect 22988 25452 23044 25454
rect 22316 24050 22372 24052
rect 22316 23998 22318 24050
rect 22318 23998 22370 24050
rect 22370 23998 22372 24050
rect 22316 23996 22372 23998
rect 22316 23266 22372 23268
rect 22316 23214 22318 23266
rect 22318 23214 22370 23266
rect 22370 23214 22372 23266
rect 22316 23212 22372 23214
rect 22204 22316 22260 22372
rect 25564 28588 25620 28644
rect 27468 32956 27524 33012
rect 29372 32844 29428 32900
rect 29036 31948 29092 32004
rect 28588 31778 28644 31780
rect 28588 31726 28590 31778
rect 28590 31726 28642 31778
rect 28642 31726 28644 31778
rect 28588 31724 28644 31726
rect 27356 31554 27412 31556
rect 27356 31502 27358 31554
rect 27358 31502 27410 31554
rect 27410 31502 27412 31554
rect 27356 31500 27412 31502
rect 27020 30322 27076 30324
rect 27020 30270 27022 30322
rect 27022 30270 27074 30322
rect 27074 30270 27076 30322
rect 27020 30268 27076 30270
rect 27244 29372 27300 29428
rect 29036 31500 29092 31556
rect 29484 32508 29540 32564
rect 29484 31724 29540 31780
rect 32956 33458 33012 33460
rect 32956 33406 32958 33458
rect 32958 33406 33010 33458
rect 33010 33406 33012 33458
rect 32956 33404 33012 33406
rect 30156 32956 30212 33012
rect 30492 33180 30548 33236
rect 30156 32732 30212 32788
rect 33964 33234 34020 33236
rect 33964 33182 33966 33234
rect 33966 33182 34018 33234
rect 34018 33182 34020 33234
rect 33964 33180 34020 33182
rect 31164 32844 31220 32900
rect 32396 32786 32452 32788
rect 32396 32734 32398 32786
rect 32398 32734 32450 32786
rect 32450 32734 32452 32786
rect 32396 32732 32452 32734
rect 31164 32562 31220 32564
rect 31164 32510 31166 32562
rect 31166 32510 31218 32562
rect 31218 32510 31220 32562
rect 31164 32508 31220 32510
rect 31948 32562 32004 32564
rect 31948 32510 31950 32562
rect 31950 32510 32002 32562
rect 32002 32510 32004 32562
rect 31948 32508 32004 32510
rect 32732 32508 32788 32564
rect 32956 33068 33012 33124
rect 30156 31948 30212 32004
rect 31388 31500 31444 31556
rect 31836 32284 31892 32340
rect 30268 31164 30324 31220
rect 28028 30098 28084 30100
rect 28028 30046 28030 30098
rect 28030 30046 28082 30098
rect 28082 30046 28084 30098
rect 28028 30044 28084 30046
rect 31948 31554 32004 31556
rect 31948 31502 31950 31554
rect 31950 31502 32002 31554
rect 32002 31502 32004 31554
rect 31948 31500 32004 31502
rect 30604 30882 30660 30884
rect 30604 30830 30606 30882
rect 30606 30830 30658 30882
rect 30658 30830 30660 30882
rect 30604 30828 30660 30830
rect 31724 30044 31780 30100
rect 31052 29986 31108 29988
rect 31052 29934 31054 29986
rect 31054 29934 31106 29986
rect 31106 29934 31108 29986
rect 31052 29932 31108 29934
rect 29596 29596 29652 29652
rect 27356 29260 27412 29316
rect 28140 29314 28196 29316
rect 28140 29262 28142 29314
rect 28142 29262 28194 29314
rect 28194 29262 28196 29314
rect 28140 29260 28196 29262
rect 28252 28700 28308 28756
rect 28028 28642 28084 28644
rect 28028 28590 28030 28642
rect 28030 28590 28082 28642
rect 28082 28590 28084 28642
rect 28028 28588 28084 28590
rect 27804 28418 27860 28420
rect 27804 28366 27806 28418
rect 27806 28366 27858 28418
rect 27858 28366 27860 28418
rect 27804 28364 27860 28366
rect 26124 26908 26180 26964
rect 25340 26178 25396 26180
rect 25340 26126 25342 26178
rect 25342 26126 25394 26178
rect 25394 26126 25396 26178
rect 25340 26124 25396 26126
rect 23436 25452 23492 25508
rect 23436 23996 23492 24052
rect 24556 23772 24612 23828
rect 24892 25564 24948 25620
rect 20636 21084 20692 21140
rect 23884 20860 23940 20916
rect 20860 20802 20916 20804
rect 20860 20750 20862 20802
rect 20862 20750 20914 20802
rect 20914 20750 20916 20802
rect 20860 20748 20916 20750
rect 20412 19740 20468 19796
rect 21196 20524 21252 20580
rect 19516 18956 19572 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 17052 17164 17108 17220
rect 20300 18284 20356 18340
rect 20748 19180 20804 19236
rect 20748 18060 20804 18116
rect 20076 17724 20132 17780
rect 20748 17778 20804 17780
rect 20748 17726 20750 17778
rect 20750 17726 20802 17778
rect 20802 17726 20804 17778
rect 20748 17724 20804 17726
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19180 17164 19236 17220
rect 17948 16828 18004 16884
rect 18396 16828 18452 16884
rect 18956 16882 19012 16884
rect 18956 16830 18958 16882
rect 18958 16830 19010 16882
rect 19010 16830 19012 16882
rect 18956 16828 19012 16830
rect 16716 15090 16772 15092
rect 16716 15038 16718 15090
rect 16718 15038 16770 15090
rect 16770 15038 16772 15090
rect 16716 15036 16772 15038
rect 13692 14924 13748 14980
rect 15820 14588 15876 14644
rect 10668 13132 10724 13188
rect 11788 12908 11844 12964
rect 10668 12684 10724 12740
rect 11228 12738 11284 12740
rect 11228 12686 11230 12738
rect 11230 12686 11282 12738
rect 11282 12686 11284 12738
rect 11228 12684 11284 12686
rect 9884 12178 9940 12180
rect 9884 12126 9886 12178
rect 9886 12126 9938 12178
rect 9938 12126 9940 12178
rect 9884 12124 9940 12126
rect 10108 12348 10164 12404
rect 10444 12124 10500 12180
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2044 9714 2100 9716
rect 2044 9662 2046 9714
rect 2046 9662 2098 9714
rect 2098 9662 2100 9714
rect 2044 9660 2100 9662
rect 1932 8930 1988 8932
rect 1932 8878 1934 8930
rect 1934 8878 1986 8930
rect 1986 8878 1988 8930
rect 1932 8876 1988 8878
rect 8204 9772 8260 9828
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 2044 8146 2100 8148
rect 2044 8094 2046 8146
rect 2046 8094 2098 8146
rect 2098 8094 2100 8146
rect 2044 8092 2100 8094
rect 1932 6748 1988 6804
rect 2716 6524 2772 6580
rect 2044 6076 2100 6132
rect 1932 5404 1988 5460
rect 2044 5068 2100 5124
rect 1708 4450 1764 4452
rect 1708 4398 1710 4450
rect 1710 4398 1762 4450
rect 1762 4398 1764 4450
rect 1708 4396 1764 4398
rect 1708 4172 1764 4228
rect 1708 3554 1764 3556
rect 1708 3502 1710 3554
rect 1710 3502 1762 3554
rect 1762 3502 1764 3554
rect 1708 3500 1764 3502
rect 2716 5180 2772 5236
rect 2380 4060 2436 4116
rect 2380 3500 2436 3556
rect 1820 1708 1876 1764
rect 3276 7420 3332 7476
rect 3276 5010 3332 5012
rect 3276 4958 3278 5010
rect 3278 4958 3330 5010
rect 3330 4958 3332 5010
rect 3276 4956 3332 4958
rect 3276 4508 3332 4564
rect 3052 3442 3108 3444
rect 3052 3390 3054 3442
rect 3054 3390 3106 3442
rect 3106 3390 3108 3442
rect 3052 3388 3108 3390
rect 2380 700 2436 756
rect 9548 9826 9604 9828
rect 9548 9774 9550 9826
rect 9550 9774 9602 9826
rect 9602 9774 9604 9826
rect 9548 9772 9604 9774
rect 8652 9436 8708 9492
rect 9996 9324 10052 9380
rect 12236 12348 12292 12404
rect 11788 12178 11844 12180
rect 11788 12126 11790 12178
rect 11790 12126 11842 12178
rect 11842 12126 11844 12178
rect 11788 12124 11844 12126
rect 12460 12962 12516 12964
rect 12460 12910 12462 12962
rect 12462 12910 12514 12962
rect 12514 12910 12516 12962
rect 12460 12908 12516 12910
rect 11564 10722 11620 10724
rect 11564 10670 11566 10722
rect 11566 10670 11618 10722
rect 11618 10670 11620 10722
rect 11564 10668 11620 10670
rect 13468 12908 13524 12964
rect 13580 11170 13636 11172
rect 13580 11118 13582 11170
rect 13582 11118 13634 11170
rect 13634 11118 13636 11170
rect 13580 11116 13636 11118
rect 12460 9996 12516 10052
rect 10556 9436 10612 9492
rect 12012 9324 12068 9380
rect 11676 9100 11732 9156
rect 9548 8876 9604 8932
rect 13020 9154 13076 9156
rect 13020 9102 13022 9154
rect 13022 9102 13074 9154
rect 13074 9102 13076 9154
rect 13020 9100 13076 9102
rect 12124 8876 12180 8932
rect 13132 7532 13188 7588
rect 16828 14476 16884 14532
rect 16604 12124 16660 12180
rect 17500 14588 17556 14644
rect 19404 16882 19460 16884
rect 19404 16830 19406 16882
rect 19406 16830 19458 16882
rect 19458 16830 19460 16882
rect 19404 16828 19460 16830
rect 18396 14924 18452 14980
rect 18508 15036 18564 15092
rect 18284 14588 18340 14644
rect 17948 12908 18004 12964
rect 18732 12908 18788 12964
rect 17500 12124 17556 12180
rect 16492 11340 16548 11396
rect 14588 11170 14644 11172
rect 14588 11118 14590 11170
rect 14590 11118 14642 11170
rect 14642 11118 14644 11170
rect 14588 11116 14644 11118
rect 15036 10780 15092 10836
rect 14364 10668 14420 10724
rect 16604 11170 16660 11172
rect 16604 11118 16606 11170
rect 16606 11118 16658 11170
rect 16658 11118 16660 11170
rect 16604 11116 16660 11118
rect 16492 10834 16548 10836
rect 16492 10782 16494 10834
rect 16494 10782 16546 10834
rect 16546 10782 16548 10834
rect 16492 10780 16548 10782
rect 21756 19234 21812 19236
rect 21756 19182 21758 19234
rect 21758 19182 21810 19234
rect 21810 19182 21812 19234
rect 21756 19180 21812 19182
rect 24444 21586 24500 21588
rect 24444 21534 24446 21586
rect 24446 21534 24498 21586
rect 24498 21534 24500 21586
rect 24444 21532 24500 21534
rect 23996 19292 24052 19348
rect 24108 21084 24164 21140
rect 25676 25228 25732 25284
rect 25116 24050 25172 24052
rect 25116 23998 25118 24050
rect 25118 23998 25170 24050
rect 25170 23998 25172 24050
rect 25116 23996 25172 23998
rect 26124 23826 26180 23828
rect 26124 23774 26126 23826
rect 26126 23774 26178 23826
rect 26178 23774 26180 23826
rect 26124 23772 26180 23774
rect 26460 27356 26516 27412
rect 29036 28700 29092 28756
rect 29036 28476 29092 28532
rect 26908 26908 26964 26964
rect 26796 26124 26852 26180
rect 26348 23324 26404 23380
rect 27244 26236 27300 26292
rect 28364 26290 28420 26292
rect 28364 26238 28366 26290
rect 28366 26238 28418 26290
rect 28418 26238 28420 26290
rect 28364 26236 28420 26238
rect 27244 25618 27300 25620
rect 27244 25566 27246 25618
rect 27246 25566 27298 25618
rect 27298 25566 27300 25618
rect 27244 25564 27300 25566
rect 28924 26178 28980 26180
rect 28924 26126 28926 26178
rect 28926 26126 28978 26178
rect 28978 26126 28980 26178
rect 28924 26124 28980 26126
rect 31388 29650 31444 29652
rect 31388 29598 31390 29650
rect 31390 29598 31442 29650
rect 31442 29598 31444 29650
rect 31388 29596 31444 29598
rect 31836 29932 31892 29988
rect 33292 32956 33348 33012
rect 32732 29484 32788 29540
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35644 33068 35700 33124
rect 36540 33068 36596 33124
rect 34412 32956 34468 33012
rect 33516 32562 33572 32564
rect 33516 32510 33518 32562
rect 33518 32510 33570 32562
rect 33570 32510 33572 32562
rect 33516 32508 33572 32510
rect 34412 32338 34468 32340
rect 34412 32286 34414 32338
rect 34414 32286 34466 32338
rect 34466 32286 34468 32338
rect 34412 32284 34468 32286
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35084 31836 35140 31892
rect 37324 33068 37380 33124
rect 37548 33964 37604 34020
rect 38444 34018 38500 34020
rect 38444 33966 38446 34018
rect 38446 33966 38498 34018
rect 38498 33966 38500 34018
rect 38444 33964 38500 33966
rect 37212 32396 37268 32452
rect 37436 31948 37492 32004
rect 37100 31890 37156 31892
rect 37100 31838 37102 31890
rect 37102 31838 37154 31890
rect 37154 31838 37156 31890
rect 37100 31836 37156 31838
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 36092 30828 36148 30884
rect 36876 30380 36932 30436
rect 36764 30268 36820 30324
rect 33404 29708 33460 29764
rect 33852 29650 33908 29652
rect 33852 29598 33854 29650
rect 33854 29598 33906 29650
rect 33906 29598 33908 29650
rect 33852 29596 33908 29598
rect 33516 29260 33572 29316
rect 30268 27356 30324 27412
rect 28812 24610 28868 24612
rect 28812 24558 28814 24610
rect 28814 24558 28866 24610
rect 28866 24558 28868 24610
rect 28812 24556 28868 24558
rect 26348 22258 26404 22260
rect 26348 22206 26350 22258
rect 26350 22206 26402 22258
rect 26402 22206 26404 22258
rect 26348 22204 26404 22206
rect 25116 21586 25172 21588
rect 25116 21534 25118 21586
rect 25118 21534 25170 21586
rect 25170 21534 25172 21586
rect 25116 21532 25172 21534
rect 24892 20914 24948 20916
rect 24892 20862 24894 20914
rect 24894 20862 24946 20914
rect 24946 20862 24948 20914
rect 24892 20860 24948 20862
rect 24444 20524 24500 20580
rect 25788 21586 25844 21588
rect 25788 21534 25790 21586
rect 25790 21534 25842 21586
rect 25842 21534 25844 21586
rect 25788 21532 25844 21534
rect 25676 19740 25732 19796
rect 26124 19346 26180 19348
rect 26124 19294 26126 19346
rect 26126 19294 26178 19346
rect 26178 19294 26180 19346
rect 26124 19292 26180 19294
rect 24892 19122 24948 19124
rect 24892 19070 24894 19122
rect 24894 19070 24946 19122
rect 24946 19070 24948 19122
rect 24892 19068 24948 19070
rect 23772 18956 23828 19012
rect 23212 18338 23268 18340
rect 23212 18286 23214 18338
rect 23214 18286 23266 18338
rect 23266 18286 23268 18338
rect 23212 18284 23268 18286
rect 21756 18172 21812 18228
rect 22876 18172 22932 18228
rect 20860 16828 20916 16884
rect 23548 16716 23604 16772
rect 22876 16658 22932 16660
rect 22876 16606 22878 16658
rect 22878 16606 22930 16658
rect 22930 16606 22932 16658
rect 22876 16604 22932 16606
rect 20524 15874 20580 15876
rect 20524 15822 20526 15874
rect 20526 15822 20578 15874
rect 20578 15822 20580 15874
rect 20524 15820 20580 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20524 15202 20580 15204
rect 20524 15150 20526 15202
rect 20526 15150 20578 15202
rect 20578 15150 20580 15202
rect 20524 15148 20580 15150
rect 21308 14812 21364 14868
rect 20748 14642 20804 14644
rect 20748 14590 20750 14642
rect 20750 14590 20802 14642
rect 20802 14590 20804 14642
rect 20748 14588 20804 14590
rect 21420 14642 21476 14644
rect 21420 14590 21422 14642
rect 21422 14590 21474 14642
rect 21474 14590 21476 14642
rect 21420 14588 21476 14590
rect 20300 14530 20356 14532
rect 20300 14478 20302 14530
rect 20302 14478 20354 14530
rect 20354 14478 20356 14530
rect 20300 14476 20356 14478
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21644 14476 21700 14532
rect 25788 19010 25844 19012
rect 25788 18958 25790 19010
rect 25790 18958 25842 19010
rect 25842 18958 25844 19010
rect 25788 18956 25844 18958
rect 24556 18562 24612 18564
rect 24556 18510 24558 18562
rect 24558 18510 24610 18562
rect 24610 18510 24612 18562
rect 24556 18508 24612 18510
rect 25788 18396 25844 18452
rect 24108 18172 24164 18228
rect 25340 16882 25396 16884
rect 25340 16830 25342 16882
rect 25342 16830 25394 16882
rect 25394 16830 25396 16882
rect 25340 16828 25396 16830
rect 24220 16716 24276 16772
rect 23772 15820 23828 15876
rect 23996 15596 24052 15652
rect 23548 15148 23604 15204
rect 22316 14812 22372 14868
rect 22204 14530 22260 14532
rect 22204 14478 22206 14530
rect 22206 14478 22258 14530
rect 22258 14478 22260 14530
rect 22204 14476 22260 14478
rect 23212 13804 23268 13860
rect 21644 12962 21700 12964
rect 21644 12910 21646 12962
rect 21646 12910 21698 12962
rect 21698 12910 21700 12962
rect 21644 12908 21700 12910
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 17948 11340 18004 11396
rect 18620 11340 18676 11396
rect 15372 10722 15428 10724
rect 15372 10670 15374 10722
rect 15374 10670 15426 10722
rect 15426 10670 15428 10722
rect 15372 10668 15428 10670
rect 17724 10610 17780 10612
rect 17724 10558 17726 10610
rect 17726 10558 17778 10610
rect 17778 10558 17780 10610
rect 17724 10556 17780 10558
rect 15372 9996 15428 10052
rect 13916 8930 13972 8932
rect 13916 8878 13918 8930
rect 13918 8878 13970 8930
rect 13970 8878 13972 8930
rect 13916 8876 13972 8878
rect 16156 9324 16212 9380
rect 17276 9324 17332 9380
rect 16716 9154 16772 9156
rect 16716 9102 16718 9154
rect 16718 9102 16770 9154
rect 16770 9102 16772 9154
rect 16716 9100 16772 9102
rect 19516 9996 19572 10052
rect 20076 11394 20132 11396
rect 20076 11342 20078 11394
rect 20078 11342 20130 11394
rect 20130 11342 20132 11394
rect 20076 11340 20132 11342
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 21196 10780 21252 10836
rect 22540 12908 22596 12964
rect 21980 11116 22036 11172
rect 20412 9100 20468 9156
rect 20972 9996 21028 10052
rect 25452 16604 25508 16660
rect 25788 15148 25844 15204
rect 26124 16828 26180 16884
rect 23996 13858 24052 13860
rect 23996 13806 23998 13858
rect 23998 13806 24050 13858
rect 24050 13806 24052 13858
rect 23996 13804 24052 13806
rect 23772 13692 23828 13748
rect 29708 27020 29764 27076
rect 31500 28530 31556 28532
rect 31500 28478 31502 28530
rect 31502 28478 31554 28530
rect 31554 28478 31556 28530
rect 31500 28476 31556 28478
rect 30492 27020 30548 27076
rect 33404 28700 33460 28756
rect 29820 26796 29876 26852
rect 30716 26796 30772 26852
rect 30156 25228 30212 25284
rect 33180 26290 33236 26292
rect 33180 26238 33182 26290
rect 33182 26238 33234 26290
rect 33234 26238 33236 26290
rect 33180 26236 33236 26238
rect 33964 29260 34020 29316
rect 34188 29708 34244 29764
rect 34300 28530 34356 28532
rect 34300 28478 34302 28530
rect 34302 28478 34354 28530
rect 34354 28478 34356 28530
rect 34300 28476 34356 28478
rect 34412 26908 34468 26964
rect 32844 25282 32900 25284
rect 32844 25230 32846 25282
rect 32846 25230 32898 25282
rect 32898 25230 32900 25282
rect 32844 25228 32900 25230
rect 33180 24946 33236 24948
rect 33180 24894 33182 24946
rect 33182 24894 33234 24946
rect 33234 24894 33236 24946
rect 33180 24892 33236 24894
rect 32732 24780 32788 24836
rect 30604 24722 30660 24724
rect 30604 24670 30606 24722
rect 30606 24670 30658 24722
rect 30658 24670 30660 24722
rect 30604 24668 30660 24670
rect 31724 24722 31780 24724
rect 31724 24670 31726 24722
rect 31726 24670 31778 24722
rect 31778 24670 31780 24722
rect 31724 24668 31780 24670
rect 31276 24220 31332 24276
rect 29260 22316 29316 22372
rect 28252 22146 28308 22148
rect 28252 22094 28254 22146
rect 28254 22094 28306 22146
rect 28306 22094 28308 22146
rect 28252 22092 28308 22094
rect 29036 21980 29092 22036
rect 33628 25394 33684 25396
rect 33628 25342 33630 25394
rect 33630 25342 33682 25394
rect 33682 25342 33684 25394
rect 33628 25340 33684 25342
rect 33740 25116 33796 25172
rect 33516 23548 33572 23604
rect 30940 22316 30996 22372
rect 29596 22146 29652 22148
rect 29596 22094 29598 22146
rect 29598 22094 29650 22146
rect 29650 22094 29652 22146
rect 29596 22092 29652 22094
rect 32060 21810 32116 21812
rect 32060 21758 32062 21810
rect 32062 21758 32114 21810
rect 32114 21758 32116 21810
rect 32060 21756 32116 21758
rect 29596 21586 29652 21588
rect 29596 21534 29598 21586
rect 29598 21534 29650 21586
rect 29650 21534 29652 21586
rect 29596 21532 29652 21534
rect 27020 20524 27076 20580
rect 27020 19740 27076 19796
rect 27132 19122 27188 19124
rect 27132 19070 27134 19122
rect 27134 19070 27186 19122
rect 27186 19070 27188 19122
rect 27132 19068 27188 19070
rect 26796 18172 26852 18228
rect 26348 17388 26404 17444
rect 26908 17442 26964 17444
rect 26908 17390 26910 17442
rect 26910 17390 26962 17442
rect 26962 17390 26964 17442
rect 26908 17388 26964 17390
rect 27580 17442 27636 17444
rect 27580 17390 27582 17442
rect 27582 17390 27634 17442
rect 27634 17390 27636 17442
rect 27580 17388 27636 17390
rect 27244 16828 27300 16884
rect 27020 15874 27076 15876
rect 27020 15822 27022 15874
rect 27022 15822 27074 15874
rect 27074 15822 27076 15874
rect 27020 15820 27076 15822
rect 27244 15260 27300 15316
rect 27804 17052 27860 17108
rect 32284 22316 32340 22372
rect 34076 24220 34132 24276
rect 34300 24162 34356 24164
rect 34300 24110 34302 24162
rect 34302 24110 34354 24162
rect 34354 24110 34356 24162
rect 34300 24108 34356 24110
rect 33180 21810 33236 21812
rect 33180 21758 33182 21810
rect 33182 21758 33234 21810
rect 33234 21758 33236 21810
rect 33180 21756 33236 21758
rect 34076 21644 34132 21700
rect 32620 21362 32676 21364
rect 32620 21310 32622 21362
rect 32622 21310 32674 21362
rect 32674 21310 32676 21362
rect 32620 21308 32676 21310
rect 32172 21196 32228 21252
rect 28812 19068 28868 19124
rect 29036 18508 29092 18564
rect 28588 18172 28644 18228
rect 28812 16994 28868 16996
rect 28812 16942 28814 16994
rect 28814 16942 28866 16994
rect 28866 16942 28868 16994
rect 28812 16940 28868 16942
rect 31388 20802 31444 20804
rect 31388 20750 31390 20802
rect 31390 20750 31442 20802
rect 31442 20750 31444 20802
rect 31388 20748 31444 20750
rect 33964 21196 34020 21252
rect 30940 20076 30996 20132
rect 32620 20076 32676 20132
rect 32508 20018 32564 20020
rect 32508 19966 32510 20018
rect 32510 19966 32562 20018
rect 32562 19966 32564 20018
rect 32508 19964 32564 19966
rect 30828 19794 30884 19796
rect 30828 19742 30830 19794
rect 30830 19742 30882 19794
rect 30882 19742 30884 19794
rect 30828 19740 30884 19742
rect 32172 19292 32228 19348
rect 30716 18450 30772 18452
rect 30716 18398 30718 18450
rect 30718 18398 30770 18450
rect 30770 18398 30772 18450
rect 30716 18396 30772 18398
rect 32508 17778 32564 17780
rect 32508 17726 32510 17778
rect 32510 17726 32562 17778
rect 32562 17726 32564 17778
rect 32508 17724 32564 17726
rect 33516 20018 33572 20020
rect 33516 19966 33518 20018
rect 33518 19966 33570 20018
rect 33570 19966 33572 20018
rect 33516 19964 33572 19966
rect 35868 30044 35924 30100
rect 34748 29596 34804 29652
rect 35308 29538 35364 29540
rect 35308 29486 35310 29538
rect 35310 29486 35362 29538
rect 35362 29486 35364 29538
rect 35308 29484 35364 29486
rect 36540 29314 36596 29316
rect 36540 29262 36542 29314
rect 36542 29262 36594 29314
rect 36594 29262 36596 29314
rect 36540 29260 36596 29262
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 38108 32562 38164 32564
rect 38108 32510 38110 32562
rect 38110 32510 38162 32562
rect 38162 32510 38164 32562
rect 38108 32508 38164 32510
rect 38108 31948 38164 32004
rect 39116 32396 39172 32452
rect 39900 32562 39956 32564
rect 39900 32510 39902 32562
rect 39902 32510 39954 32562
rect 39954 32510 39956 32562
rect 39900 32508 39956 32510
rect 40460 32396 40516 32452
rect 37884 30882 37940 30884
rect 37884 30830 37886 30882
rect 37886 30830 37938 30882
rect 37938 30830 37940 30882
rect 37884 30828 37940 30830
rect 37324 30044 37380 30100
rect 37548 29932 37604 29988
rect 36988 29260 37044 29316
rect 35308 28754 35364 28756
rect 35308 28702 35310 28754
rect 35310 28702 35362 28754
rect 35362 28702 35364 28754
rect 35308 28700 35364 28702
rect 35084 28642 35140 28644
rect 35084 28590 35086 28642
rect 35086 28590 35138 28642
rect 35138 28590 35140 28642
rect 35084 28588 35140 28590
rect 34636 27132 34692 27188
rect 34524 25340 34580 25396
rect 36316 28642 36372 28644
rect 36316 28590 36318 28642
rect 36318 28590 36370 28642
rect 36370 28590 36372 28642
rect 36316 28588 36372 28590
rect 37660 28418 37716 28420
rect 37660 28366 37662 28418
rect 37662 28366 37714 28418
rect 37714 28366 37716 28418
rect 37660 28364 37716 28366
rect 39116 30380 39172 30436
rect 38892 30268 38948 30324
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35980 26962 36036 26964
rect 35980 26910 35982 26962
rect 35982 26910 36034 26962
rect 36034 26910 36036 26962
rect 35980 26908 36036 26910
rect 36876 26460 36932 26516
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 36988 25788 37044 25844
rect 35644 25116 35700 25172
rect 35084 24892 35140 24948
rect 35308 24834 35364 24836
rect 35308 24782 35310 24834
rect 35310 24782 35362 24834
rect 35362 24782 35364 24834
rect 35308 24780 35364 24782
rect 36316 25506 36372 25508
rect 36316 25454 36318 25506
rect 36318 25454 36370 25506
rect 36370 25454 36372 25506
rect 36316 25452 36372 25454
rect 36092 25116 36148 25172
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35084 23996 35140 24052
rect 35756 24050 35812 24052
rect 35756 23998 35758 24050
rect 35758 23998 35810 24050
rect 35810 23998 35812 24050
rect 35756 23996 35812 23998
rect 37100 25506 37156 25508
rect 37100 25454 37102 25506
rect 37102 25454 37154 25506
rect 37154 25454 37156 25506
rect 37100 25452 37156 25454
rect 37996 27186 38052 27188
rect 37996 27134 37998 27186
rect 37998 27134 38050 27186
rect 38050 27134 38052 27186
rect 37996 27132 38052 27134
rect 38780 26514 38836 26516
rect 38780 26462 38782 26514
rect 38782 26462 38834 26514
rect 38834 26462 38836 26514
rect 38780 26460 38836 26462
rect 38892 25788 38948 25844
rect 38668 24892 38724 24948
rect 39116 24722 39172 24724
rect 39116 24670 39118 24722
rect 39118 24670 39170 24722
rect 39170 24670 39172 24722
rect 39116 24668 39172 24670
rect 39900 29426 39956 29428
rect 39900 29374 39902 29426
rect 39902 29374 39954 29426
rect 39954 29374 39956 29426
rect 39900 29372 39956 29374
rect 39788 29260 39844 29316
rect 40236 29596 40292 29652
rect 39900 28364 39956 28420
rect 39340 25676 39396 25732
rect 37884 24108 37940 24164
rect 34972 23548 35028 23604
rect 34972 23100 35028 23156
rect 36092 23154 36148 23156
rect 36092 23102 36094 23154
rect 36094 23102 36146 23154
rect 36146 23102 36148 23154
rect 36092 23100 36148 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22540 35140 22596
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 20914 35252 20916
rect 35196 20862 35198 20914
rect 35198 20862 35250 20914
rect 35250 20862 35252 20914
rect 35196 20860 35252 20862
rect 35084 19964 35140 20020
rect 34972 19122 35028 19124
rect 34972 19070 34974 19122
rect 34974 19070 35026 19122
rect 35026 19070 35028 19122
rect 34972 19068 35028 19070
rect 32620 18284 32676 18340
rect 32396 17612 32452 17668
rect 30044 17052 30100 17108
rect 31052 16994 31108 16996
rect 31052 16942 31054 16994
rect 31054 16942 31106 16994
rect 31106 16942 31108 16994
rect 31052 16940 31108 16942
rect 31500 16716 31556 16772
rect 27692 15260 27748 15316
rect 28700 15820 28756 15876
rect 28588 15260 28644 15316
rect 29932 15314 29988 15316
rect 29932 15262 29934 15314
rect 29934 15262 29986 15314
rect 29986 15262 29988 15314
rect 29932 15260 29988 15262
rect 30716 15596 30772 15652
rect 27580 15202 27636 15204
rect 27580 15150 27582 15202
rect 27582 15150 27634 15202
rect 27634 15150 27636 15202
rect 27580 15148 27636 15150
rect 26124 13746 26180 13748
rect 26124 13694 26126 13746
rect 26126 13694 26178 13746
rect 26178 13694 26180 13746
rect 26124 13692 26180 13694
rect 24780 13132 24836 13188
rect 26908 13132 26964 13188
rect 26796 12738 26852 12740
rect 26796 12686 26798 12738
rect 26798 12686 26850 12738
rect 26850 12686 26852 12738
rect 26796 12684 26852 12686
rect 24332 11452 24388 11508
rect 23548 11004 23604 11060
rect 24332 11004 24388 11060
rect 22652 10834 22708 10836
rect 22652 10782 22654 10834
rect 22654 10782 22706 10834
rect 22706 10782 22708 10834
rect 22652 10780 22708 10782
rect 22540 10610 22596 10612
rect 22540 10558 22542 10610
rect 22542 10558 22594 10610
rect 22594 10558 22596 10610
rect 22540 10556 22596 10558
rect 25900 11564 25956 11620
rect 25676 11506 25732 11508
rect 25676 11454 25678 11506
rect 25678 11454 25730 11506
rect 25730 11454 25732 11506
rect 25676 11452 25732 11454
rect 25116 10668 25172 10724
rect 26236 10722 26292 10724
rect 26236 10670 26238 10722
rect 26238 10670 26290 10722
rect 26290 10670 26292 10722
rect 26236 10668 26292 10670
rect 29484 14252 29540 14308
rect 27356 13804 27412 13860
rect 28588 13692 28644 13748
rect 28252 13580 28308 13636
rect 27692 12738 27748 12740
rect 27692 12686 27694 12738
rect 27694 12686 27746 12738
rect 27746 12686 27748 12738
rect 27692 12684 27748 12686
rect 27580 11618 27636 11620
rect 27580 11566 27582 11618
rect 27582 11566 27634 11618
rect 27634 11566 27636 11618
rect 27580 11564 27636 11566
rect 29260 12962 29316 12964
rect 29260 12910 29262 12962
rect 29262 12910 29314 12962
rect 29314 12910 29316 12962
rect 29260 12908 29316 12910
rect 33516 18450 33572 18452
rect 33516 18398 33518 18450
rect 33518 18398 33570 18450
rect 33570 18398 33572 18450
rect 33516 18396 33572 18398
rect 33628 17724 33684 17780
rect 32620 16716 32676 16772
rect 33180 16716 33236 16772
rect 31948 14588 32004 14644
rect 29820 14364 29876 14420
rect 30940 14418 30996 14420
rect 30940 14366 30942 14418
rect 30942 14366 30994 14418
rect 30994 14366 30996 14418
rect 30940 14364 30996 14366
rect 32844 14306 32900 14308
rect 32844 14254 32846 14306
rect 32846 14254 32898 14306
rect 32898 14254 32900 14306
rect 32844 14252 32900 14254
rect 32060 13858 32116 13860
rect 32060 13806 32062 13858
rect 32062 13806 32114 13858
rect 32114 13806 32116 13858
rect 32060 13804 32116 13806
rect 31052 13634 31108 13636
rect 31052 13582 31054 13634
rect 31054 13582 31106 13634
rect 31106 13582 31108 13634
rect 31052 13580 31108 13582
rect 32060 13020 32116 13076
rect 30044 12908 30100 12964
rect 30044 12124 30100 12180
rect 27580 9826 27636 9828
rect 27580 9774 27582 9826
rect 27582 9774 27634 9826
rect 27634 9774 27636 9826
rect 27580 9772 27636 9774
rect 32732 12850 32788 12852
rect 32732 12798 32734 12850
rect 32734 12798 32786 12850
rect 32786 12798 32788 12850
rect 32732 12796 32788 12798
rect 30156 10668 30212 10724
rect 32620 12178 32676 12180
rect 32620 12126 32622 12178
rect 32622 12126 32674 12178
rect 32674 12126 32676 12178
rect 32620 12124 32676 12126
rect 32172 10668 32228 10724
rect 34636 17778 34692 17780
rect 34636 17726 34638 17778
rect 34638 17726 34690 17778
rect 34690 17726 34692 17778
rect 34636 17724 34692 17726
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35868 18396 35924 18452
rect 35308 18338 35364 18340
rect 35308 18286 35310 18338
rect 35310 18286 35362 18338
rect 35362 18286 35364 18338
rect 35308 18284 35364 18286
rect 36204 18284 36260 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 17612 35140 17668
rect 35420 17724 35476 17780
rect 35532 16940 35588 16996
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37100 23100 37156 23156
rect 37772 22540 37828 22596
rect 36764 21868 36820 21924
rect 37436 21810 37492 21812
rect 37436 21758 37438 21810
rect 37438 21758 37490 21810
rect 37490 21758 37492 21810
rect 37436 21756 37492 21758
rect 39004 22258 39060 22260
rect 39004 22206 39006 22258
rect 39006 22206 39058 22258
rect 39058 22206 39060 22258
rect 39004 22204 39060 22206
rect 37996 21532 38052 21588
rect 38220 21868 38276 21924
rect 37772 21420 37828 21476
rect 36540 17500 36596 17556
rect 37212 20914 37268 20916
rect 37212 20862 37214 20914
rect 37214 20862 37266 20914
rect 37266 20862 37268 20914
rect 37212 20860 37268 20862
rect 37996 20914 38052 20916
rect 37996 20862 37998 20914
rect 37998 20862 38050 20914
rect 38050 20862 38052 20914
rect 37996 20860 38052 20862
rect 37212 20188 37268 20244
rect 36204 16828 36260 16884
rect 34412 15874 34468 15876
rect 34412 15822 34414 15874
rect 34414 15822 34466 15874
rect 34466 15822 34468 15874
rect 34412 15820 34468 15822
rect 35308 15874 35364 15876
rect 35308 15822 35310 15874
rect 35310 15822 35362 15874
rect 35362 15822 35364 15874
rect 35308 15820 35364 15822
rect 36428 16940 36484 16996
rect 37884 19964 37940 20020
rect 37996 19516 38052 19572
rect 37996 19346 38052 19348
rect 37996 19294 37998 19346
rect 37998 19294 38050 19346
rect 38050 19294 38052 19346
rect 37996 19292 38052 19294
rect 37884 17388 37940 17444
rect 37212 16882 37268 16884
rect 37212 16830 37214 16882
rect 37214 16830 37266 16882
rect 37266 16830 37268 16882
rect 37212 16828 37268 16830
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 36316 15148 36372 15204
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34972 14642 35028 14644
rect 34972 14590 34974 14642
rect 34974 14590 35026 14642
rect 35026 14590 35028 14642
rect 34972 14588 35028 14590
rect 37100 15148 37156 15204
rect 33292 13804 33348 13860
rect 35868 13858 35924 13860
rect 35868 13806 35870 13858
rect 35870 13806 35922 13858
rect 35922 13806 35924 13858
rect 35868 13804 35924 13806
rect 33068 12124 33124 12180
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 33964 13074 34020 13076
rect 33964 13022 33966 13074
rect 33966 13022 34018 13074
rect 34018 13022 34020 13074
rect 33964 13020 34020 13022
rect 34972 12850 35028 12852
rect 34972 12798 34974 12850
rect 34974 12798 35026 12850
rect 35026 12798 35028 12850
rect 34972 12796 35028 12798
rect 34076 12178 34132 12180
rect 34076 12126 34078 12178
rect 34078 12126 34130 12178
rect 34130 12126 34132 12178
rect 34076 12124 34132 12126
rect 33740 11170 33796 11172
rect 33740 11118 33742 11170
rect 33742 11118 33794 11170
rect 33794 11118 33796 11170
rect 33740 11116 33796 11118
rect 36988 13468 37044 13524
rect 38108 16828 38164 16884
rect 38444 21810 38500 21812
rect 38444 21758 38446 21810
rect 38446 21758 38498 21810
rect 38498 21758 38500 21810
rect 38444 21756 38500 21758
rect 39900 24722 39956 24724
rect 39900 24670 39902 24722
rect 39902 24670 39954 24722
rect 39954 24670 39956 24722
rect 39900 24668 39956 24670
rect 39900 22594 39956 22596
rect 39900 22542 39902 22594
rect 39902 22542 39954 22594
rect 39954 22542 39956 22594
rect 39900 22540 39956 22542
rect 40796 32396 40852 32452
rect 41020 29986 41076 29988
rect 41020 29934 41022 29986
rect 41022 29934 41074 29986
rect 41074 29934 41076 29986
rect 41020 29932 41076 29934
rect 40908 29596 40964 29652
rect 40572 29372 40628 29428
rect 40460 29260 40516 29316
rect 40796 25730 40852 25732
rect 40796 25678 40798 25730
rect 40798 25678 40850 25730
rect 40850 25678 40852 25730
rect 40796 25676 40852 25678
rect 40124 23154 40180 23156
rect 40124 23102 40126 23154
rect 40126 23102 40178 23154
rect 40178 23102 40180 23154
rect 40124 23100 40180 23102
rect 40012 22428 40068 22484
rect 41020 22482 41076 22484
rect 41020 22430 41022 22482
rect 41022 22430 41074 22482
rect 41074 22430 41076 22482
rect 41020 22428 41076 22430
rect 38668 21586 38724 21588
rect 38668 21534 38670 21586
rect 38670 21534 38722 21586
rect 38722 21534 38724 21586
rect 38668 21532 38724 21534
rect 39788 21586 39844 21588
rect 39788 21534 39790 21586
rect 39790 21534 39842 21586
rect 39842 21534 39844 21586
rect 39788 21532 39844 21534
rect 39004 21308 39060 21364
rect 38556 20188 38612 20244
rect 39004 19740 39060 19796
rect 39564 19516 39620 19572
rect 38780 18396 38836 18452
rect 38668 17612 38724 17668
rect 39004 17554 39060 17556
rect 39004 17502 39006 17554
rect 39006 17502 39058 17554
rect 39058 17502 39060 17554
rect 39004 17500 39060 17502
rect 38668 16940 38724 16996
rect 39788 17666 39844 17668
rect 39788 17614 39790 17666
rect 39790 17614 39842 17666
rect 39842 17614 39844 17666
rect 39788 17612 39844 17614
rect 41020 17666 41076 17668
rect 41020 17614 41022 17666
rect 41022 17614 41074 17666
rect 41074 17614 41076 17666
rect 41020 17612 41076 17614
rect 38892 16828 38948 16884
rect 37100 13356 37156 13412
rect 38108 13468 38164 13524
rect 36652 12012 36708 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36540 11676 36596 11732
rect 36988 11676 37044 11732
rect 38332 13244 38388 13300
rect 39340 13356 39396 13412
rect 39228 12908 39284 12964
rect 39900 17442 39956 17444
rect 39900 17390 39902 17442
rect 39902 17390 39954 17442
rect 39954 17390 39956 17442
rect 39900 17388 39956 17390
rect 39788 12908 39844 12964
rect 37884 12012 37940 12068
rect 34972 11116 35028 11172
rect 37772 10780 37828 10836
rect 39228 11788 39284 11844
rect 38444 11676 38500 11732
rect 40460 15090 40516 15092
rect 40460 15038 40462 15090
rect 40462 15038 40514 15090
rect 40514 15038 40516 15090
rect 40460 15036 40516 15038
rect 39900 11452 39956 11508
rect 39116 10780 39172 10836
rect 34748 10444 34804 10500
rect 28028 9772 28084 9828
rect 28588 9826 28644 9828
rect 28588 9774 28590 9826
rect 28590 9774 28642 9826
rect 28642 9774 28644 9826
rect 28588 9772 28644 9774
rect 29484 9826 29540 9828
rect 29484 9774 29486 9826
rect 29486 9774 29538 9826
rect 29538 9774 29540 9826
rect 29484 9772 29540 9774
rect 30492 9826 30548 9828
rect 30492 9774 30494 9826
rect 30494 9774 30546 9826
rect 30546 9774 30548 9826
rect 30492 9772 30548 9774
rect 36876 10498 36932 10500
rect 36876 10446 36878 10498
rect 36878 10446 36930 10498
rect 36930 10446 36932 10498
rect 36876 10444 36932 10446
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 32060 9772 32116 9828
rect 41468 15036 41524 15092
rect 40348 13468 40404 13524
rect 40348 13244 40404 13300
rect 40124 12962 40180 12964
rect 40124 12910 40126 12962
rect 40126 12910 40178 12962
rect 40178 12910 40180 12962
rect 40124 12908 40180 12910
rect 40684 11506 40740 11508
rect 40684 11454 40686 11506
rect 40686 11454 40738 11506
rect 40738 11454 40740 11506
rect 40684 11452 40740 11454
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 14252 7586 14308 7588
rect 14252 7534 14254 7586
rect 14254 7534 14306 7586
rect 14306 7534 14308 7586
rect 14252 7532 14308 7534
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 4284 6524 4340 6580
rect 3836 5180 3892 5236
rect 3724 4956 3780 5012
rect 3612 4562 3668 4564
rect 3612 4510 3614 4562
rect 3614 4510 3666 4562
rect 3666 4510 3668 4562
rect 3612 4508 3668 4510
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 4508 5122 4564 5124
rect 4508 5070 4510 5122
rect 4510 5070 4562 5122
rect 4562 5070 4564 5122
rect 4508 5068 4564 5070
rect 4844 4450 4900 4452
rect 4844 4398 4846 4450
rect 4846 4398 4898 4450
rect 4898 4398 4900 4450
rect 4844 4396 4900 4398
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5740 4226 5796 4228
rect 5740 4174 5742 4226
rect 5742 4174 5794 4226
rect 5794 4174 5796 4226
rect 5740 4172 5796 4174
rect 5292 3500 5348 3556
rect 4956 3442 5012 3444
rect 4956 3390 4958 3442
rect 4958 3390 5010 3442
rect 5010 3390 5012 3442
rect 4956 3388 5012 3390
rect 3948 2716 4004 2772
rect 3836 2044 3892 2100
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 8092 3276 8148 3332
rect 9324 3330 9380 3332
rect 9324 3278 9326 3330
rect 9326 3278 9378 3330
rect 9378 3278 9380 3330
rect 9324 3276 9380 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 2940 28 2996 84
<< metal3 >>
rect 0 43764 800 43792
rect 0 43708 4340 43764
rect 0 43680 800 43708
rect 4284 43204 4340 43708
rect 4274 43148 4284 43204
rect 4340 43148 4350 43204
rect 0 43092 800 43120
rect 0 43036 1932 43092
rect 1988 43036 1998 43092
rect 0 43008 800 43036
rect 0 42420 800 42448
rect 0 42364 3388 42420
rect 3444 42364 3454 42420
rect 0 42336 800 42364
rect 0 41748 800 41776
rect 0 41692 3724 41748
rect 3780 41692 3790 41748
rect 0 41664 800 41692
rect 4274 41132 4284 41188
rect 4340 41132 9548 41188
rect 9604 41132 9614 41188
rect 0 41076 800 41104
rect 0 41020 3388 41076
rect 3444 41020 3454 41076
rect 0 40992 800 41020
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 1810 40572 1820 40628
rect 1876 40572 4732 40628
rect 4788 40572 4798 40628
rect 18162 40572 18172 40628
rect 18228 40572 19180 40628
rect 19236 40572 19246 40628
rect 19842 40572 19852 40628
rect 19908 40572 20972 40628
rect 21028 40572 21038 40628
rect 4946 40460 4956 40516
rect 5012 40460 5740 40516
rect 5796 40460 5806 40516
rect 0 40404 800 40432
rect 0 40348 2100 40404
rect 3266 40348 3276 40404
rect 3332 40348 5628 40404
rect 5684 40348 5694 40404
rect 0 40320 800 40348
rect 2044 40292 2100 40348
rect 2034 40236 2044 40292
rect 2100 40236 2110 40292
rect 9426 40236 9436 40292
rect 9492 40236 10556 40292
rect 10612 40236 10622 40292
rect 25106 40236 25116 40292
rect 25172 40236 26572 40292
rect 26628 40236 26638 40292
rect 18 40124 28 40180
rect 84 40124 8428 40180
rect 8484 40124 8494 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 16146 39788 16156 39844
rect 16212 39788 16828 39844
rect 16884 39788 16894 39844
rect 0 39732 800 39760
rect 0 39676 3948 39732
rect 4004 39676 4014 39732
rect 22866 39676 22876 39732
rect 22932 39676 23996 39732
rect 24052 39676 24062 39732
rect 0 39648 800 39676
rect 3266 39340 3276 39396
rect 3332 39340 6860 39396
rect 6916 39340 6926 39396
rect 9986 39340 9996 39396
rect 10052 39340 16380 39396
rect 16436 39340 16446 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 1148 39116 7308 39172
rect 7364 39116 7868 39172
rect 7924 39116 7934 39172
rect 10658 39116 10668 39172
rect 10724 39116 17052 39172
rect 17108 39116 17118 39172
rect 0 39060 800 39088
rect 1148 39060 1204 39116
rect 0 39004 1204 39060
rect 1362 39004 1372 39060
rect 1428 39004 2156 39060
rect 2212 39004 2222 39060
rect 5730 39004 5740 39060
rect 5796 39004 5806 39060
rect 8418 39004 8428 39060
rect 8484 39004 9660 39060
rect 9716 39004 9726 39060
rect 0 38976 800 39004
rect 5740 38948 5796 39004
rect 2930 38892 2940 38948
rect 2996 38892 4844 38948
rect 4900 38892 4910 38948
rect 5740 38892 6188 38948
rect 6244 38892 6254 38948
rect 8306 38892 8316 38948
rect 8372 38892 24556 38948
rect 24612 38892 24622 38948
rect 1922 38780 1932 38836
rect 1988 38780 5068 38836
rect 5124 38780 5134 38836
rect 8082 38780 8092 38836
rect 8148 38780 8428 38836
rect 8372 38724 8428 38780
rect 4946 38668 4956 38724
rect 5012 38668 7644 38724
rect 7700 38668 7710 38724
rect 8372 38668 10220 38724
rect 10276 38668 26460 38724
rect 26516 38668 26526 38724
rect 7298 38556 7308 38612
rect 7364 38556 26124 38612
rect 26180 38556 26190 38612
rect 9314 38444 9324 38500
rect 9380 38444 15148 38500
rect 15204 38444 15214 38500
rect 0 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 0 38332 3388 38388
rect 3490 38332 3500 38388
rect 3556 38332 4172 38388
rect 4228 38332 4238 38388
rect 9090 38332 9100 38388
rect 9156 38332 19068 38388
rect 19124 38332 19134 38388
rect 0 38304 800 38332
rect 3332 38276 3388 38332
rect 3332 38220 5516 38276
rect 5572 38220 5582 38276
rect 8306 38220 8316 38276
rect 8372 38220 20748 38276
rect 20804 38220 20814 38276
rect 4050 38108 4060 38164
rect 4116 38108 6636 38164
rect 6692 38108 6702 38164
rect 9762 38108 9772 38164
rect 9828 38108 21756 38164
rect 21812 38108 21822 38164
rect 7970 37996 7980 38052
rect 8036 37996 22428 38052
rect 22484 37996 22494 38052
rect 4722 37884 4732 37940
rect 4788 37884 5292 37940
rect 5348 37884 5358 37940
rect 7634 37884 7644 37940
rect 7700 37884 23772 37940
rect 23828 37884 23838 37940
rect 2706 37772 2716 37828
rect 2772 37772 3276 37828
rect 3332 37772 3342 37828
rect 5590 37772 5628 37828
rect 5684 37772 5694 37828
rect 8642 37772 8652 37828
rect 8708 37772 18508 37828
rect 18564 37772 18574 37828
rect 0 37716 800 37744
rect 0 37660 1596 37716
rect 1652 37660 1662 37716
rect 0 37632 800 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 2930 37436 2940 37492
rect 2996 37436 4396 37492
rect 4452 37436 4462 37492
rect 4834 37436 4844 37492
rect 4900 37436 5740 37492
rect 5796 37436 5806 37492
rect 3574 37212 3612 37268
rect 3668 37212 3678 37268
rect 2706 37100 2716 37156
rect 2772 37100 6636 37156
rect 6692 37100 6702 37156
rect 8194 37100 8204 37156
rect 8260 37100 8988 37156
rect 9044 37100 25788 37156
rect 25844 37100 25854 37156
rect 0 37044 800 37072
rect 0 36988 3612 37044
rect 3668 36988 3678 37044
rect 0 36960 800 36988
rect 3332 36876 3948 36932
rect 4004 36876 4014 36932
rect 802 36764 812 36820
rect 868 36764 2380 36820
rect 2436 36764 2446 36820
rect 3332 36708 3388 36876
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 2818 36652 2828 36708
rect 2884 36652 3388 36708
rect 1586 36428 1596 36484
rect 1652 36428 4396 36484
rect 4452 36428 4462 36484
rect 0 36372 800 36400
rect 0 36316 1932 36372
rect 1988 36316 2380 36372
rect 2436 36316 2446 36372
rect 3378 36316 3388 36372
rect 3444 36316 4060 36372
rect 4116 36316 4126 36372
rect 0 36288 800 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 1698 35980 1708 36036
rect 1764 35980 1774 36036
rect 2370 35980 2380 36036
rect 2436 35980 3276 36036
rect 3332 35980 3342 36036
rect 0 35700 800 35728
rect 1708 35700 1764 35980
rect 3266 35756 3276 35812
rect 3332 35756 9548 35812
rect 9604 35756 9614 35812
rect 0 35644 1764 35700
rect 0 35616 800 35644
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 2146 35196 2156 35252
rect 2212 35196 4172 35252
rect 4228 35196 4238 35252
rect 3266 35084 3276 35140
rect 3332 35084 3948 35140
rect 4004 35084 4014 35140
rect 0 35028 800 35056
rect 0 34972 1708 35028
rect 1764 34972 1774 35028
rect 0 34944 800 34972
rect 2828 34860 3164 34916
rect 3220 34860 3230 34916
rect 2828 34692 2884 34860
rect 2818 34636 2828 34692
rect 2884 34636 2894 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 0 34356 800 34384
rect 0 34300 2044 34356
rect 2100 34300 2110 34356
rect 0 34272 800 34300
rect 37538 33964 37548 34020
rect 37604 33964 38444 34020
rect 38500 33964 38510 34020
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 0 33628 1708 33684
rect 1764 33628 1774 33684
rect 0 33600 800 33628
rect 24770 33516 24780 33572
rect 24836 33516 27244 33572
rect 27300 33516 27310 33572
rect 14018 33404 14028 33460
rect 14084 33404 15148 33460
rect 15204 33404 15214 33460
rect 26338 33404 26348 33460
rect 26404 33404 27132 33460
rect 27188 33404 27198 33460
rect 29586 33404 29596 33460
rect 29652 33404 32956 33460
rect 33012 33404 33022 33460
rect 2034 33180 2044 33236
rect 2100 33180 7196 33236
rect 7252 33180 7262 33236
rect 30482 33180 30492 33236
rect 30548 33180 33964 33236
rect 34020 33180 34030 33236
rect 17266 33068 17276 33124
rect 17332 33068 19740 33124
rect 19796 33068 19806 33124
rect 32946 33068 32956 33124
rect 33012 33068 35644 33124
rect 35700 33068 35710 33124
rect 36530 33068 36540 33124
rect 36596 33068 37324 33124
rect 37380 33068 37390 33124
rect 0 33012 800 33040
rect 0 32956 1708 33012
rect 1764 32956 2492 33012
rect 2548 32956 2558 33012
rect 23986 32956 23996 33012
rect 24052 32956 26236 33012
rect 26292 32956 26302 33012
rect 27458 32956 27468 33012
rect 27524 32956 30156 33012
rect 30212 32956 30222 33012
rect 33282 32956 33292 33012
rect 33348 32956 34412 33012
rect 34468 32956 34478 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 29362 32844 29372 32900
rect 29428 32844 31164 32900
rect 31220 32844 31230 32900
rect 30146 32732 30156 32788
rect 30212 32732 32396 32788
rect 32452 32732 32462 32788
rect 4946 32620 4956 32676
rect 5012 32620 5740 32676
rect 5796 32620 5806 32676
rect 19170 32620 19180 32676
rect 19236 32620 20076 32676
rect 20132 32620 20142 32676
rect 3266 32508 3276 32564
rect 3332 32508 3724 32564
rect 3780 32508 3790 32564
rect 29474 32508 29484 32564
rect 29540 32508 31164 32564
rect 31220 32508 31948 32564
rect 32004 32508 32732 32564
rect 32788 32508 33516 32564
rect 33572 32508 33582 32564
rect 38098 32508 38108 32564
rect 38164 32508 39900 32564
rect 39956 32508 39966 32564
rect 24658 32396 24668 32452
rect 24724 32396 26012 32452
rect 26068 32396 26078 32452
rect 37202 32396 37212 32452
rect 37268 32396 39116 32452
rect 39172 32396 40460 32452
rect 40516 32396 40796 32452
rect 40852 32396 40862 32452
rect 0 32340 800 32368
rect 0 32284 1708 32340
rect 1764 32284 1774 32340
rect 31826 32284 31836 32340
rect 31892 32284 34412 32340
rect 34468 32284 34478 32340
rect 0 32256 800 32284
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 29026 31948 29036 32004
rect 29092 31948 30156 32004
rect 30212 31948 30222 32004
rect 37426 31948 37436 32004
rect 37492 31948 38108 32004
rect 38164 31948 38174 32004
rect 8082 31836 8092 31892
rect 8148 31836 15036 31892
rect 15092 31836 15102 31892
rect 35074 31836 35084 31892
rect 35140 31836 37100 31892
rect 37156 31836 37166 31892
rect 16146 31724 16156 31780
rect 16212 31724 24556 31780
rect 24612 31724 24622 31780
rect 28578 31724 28588 31780
rect 28644 31724 29484 31780
rect 29540 31724 29550 31780
rect 0 31668 800 31696
rect 0 31612 1932 31668
rect 1988 31612 1998 31668
rect 0 31584 800 31612
rect 18386 31500 18396 31556
rect 18452 31500 20300 31556
rect 20356 31500 20366 31556
rect 27346 31500 27356 31556
rect 27412 31500 29036 31556
rect 29092 31500 29102 31556
rect 31378 31500 31388 31556
rect 31444 31500 31948 31556
rect 32004 31500 32014 31556
rect 6178 31388 6188 31444
rect 6244 31388 8764 31444
rect 8820 31388 8830 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 8978 31164 8988 31220
rect 9044 31164 9660 31220
rect 9716 31164 11228 31220
rect 11284 31164 11676 31220
rect 11732 31164 14588 31220
rect 14644 31164 15596 31220
rect 15652 31164 15662 31220
rect 25666 31164 25676 31220
rect 25732 31164 30268 31220
rect 30324 31164 30334 31220
rect 2034 31052 2044 31108
rect 2100 31052 2110 31108
rect 3332 31052 6412 31108
rect 6468 31052 6478 31108
rect 17826 31052 17836 31108
rect 17892 31052 18732 31108
rect 18788 31052 18798 31108
rect 0 30996 800 31024
rect 2044 30996 2100 31052
rect 3332 30996 3388 31052
rect 0 30940 2100 30996
rect 2930 30940 2940 30996
rect 2996 30940 3388 30996
rect 4620 30940 5964 30996
rect 6020 30940 6030 30996
rect 0 30912 800 30940
rect 4620 30884 4676 30940
rect 2034 30828 2044 30884
rect 2100 30828 4676 30884
rect 6066 30828 6076 30884
rect 6132 30828 6860 30884
rect 6916 30828 6926 30884
rect 8306 30828 8316 30884
rect 8372 30828 10108 30884
rect 10164 30828 10174 30884
rect 21746 30828 21756 30884
rect 21812 30828 30604 30884
rect 30660 30828 30670 30884
rect 36082 30828 36092 30884
rect 36148 30828 37884 30884
rect 37940 30828 37950 30884
rect 2706 30716 2716 30772
rect 2772 30716 3164 30772
rect 3220 30716 3230 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 9762 30492 9772 30548
rect 9828 30492 10892 30548
rect 10948 30492 10958 30548
rect 14354 30492 14364 30548
rect 14420 30492 15932 30548
rect 15988 30492 15998 30548
rect 36866 30380 36876 30436
rect 36932 30380 39116 30436
rect 39172 30380 39182 30436
rect 0 30324 800 30352
rect 0 30268 2380 30324
rect 2436 30268 3164 30324
rect 3220 30268 3230 30324
rect 24770 30268 24780 30324
rect 24836 30268 27020 30324
rect 27076 30268 27086 30324
rect 36754 30268 36764 30324
rect 36820 30268 38892 30324
rect 38948 30268 38958 30324
rect 0 30240 800 30268
rect 5730 30156 5740 30212
rect 5796 30156 7756 30212
rect 7812 30156 8652 30212
rect 8708 30156 8718 30212
rect 10322 30156 10332 30212
rect 10388 30156 11004 30212
rect 11060 30156 11676 30212
rect 11732 30156 12572 30212
rect 12628 30156 12638 30212
rect 13458 30156 13468 30212
rect 13524 30156 15708 30212
rect 15764 30156 17388 30212
rect 17444 30156 17454 30212
rect 22194 30156 22204 30212
rect 22260 30156 23324 30212
rect 23380 30156 23390 30212
rect 8754 30044 8764 30100
rect 8820 30044 11452 30100
rect 11508 30044 11518 30100
rect 13122 30044 13132 30100
rect 13188 30044 14924 30100
rect 14980 30044 14990 30100
rect 20290 30044 20300 30100
rect 20356 30044 21532 30100
rect 21588 30044 21598 30100
rect 21746 30044 21756 30100
rect 21812 30044 24668 30100
rect 24724 30044 24734 30100
rect 25778 30044 25788 30100
rect 25844 30044 28028 30100
rect 28084 30044 28094 30100
rect 31714 30044 31724 30100
rect 31780 30044 35868 30100
rect 35924 30044 37324 30100
rect 37380 30044 37390 30100
rect 21756 29988 21812 30044
rect 16706 29932 16716 29988
rect 16772 29932 19404 29988
rect 19460 29932 19470 29988
rect 20178 29932 20188 29988
rect 20244 29932 21196 29988
rect 21252 29932 21812 29988
rect 31042 29932 31052 29988
rect 31108 29932 31836 29988
rect 31892 29932 31902 29988
rect 37538 29932 37548 29988
rect 37604 29932 41020 29988
rect 41076 29932 41086 29988
rect 2034 29820 2044 29876
rect 2100 29820 6524 29876
rect 6580 29820 6590 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 22754 29708 22764 29764
rect 22820 29708 26236 29764
rect 26292 29708 26302 29764
rect 33394 29708 33404 29764
rect 33460 29708 34188 29764
rect 34244 29708 34254 29764
rect 0 29652 800 29680
rect 0 29596 1708 29652
rect 1764 29596 3612 29652
rect 3668 29596 3678 29652
rect 9650 29596 9660 29652
rect 9716 29596 10668 29652
rect 10724 29596 12236 29652
rect 12292 29596 12302 29652
rect 29586 29596 29596 29652
rect 29652 29596 31388 29652
rect 31444 29596 31454 29652
rect 33842 29596 33852 29652
rect 33908 29596 34748 29652
rect 34804 29596 34814 29652
rect 40226 29596 40236 29652
rect 40292 29596 40908 29652
rect 40964 29596 40974 29652
rect 0 29568 800 29596
rect 16146 29484 16156 29540
rect 16212 29484 19404 29540
rect 19460 29484 19470 29540
rect 23538 29484 23548 29540
rect 23604 29484 24332 29540
rect 24388 29484 24398 29540
rect 32722 29484 32732 29540
rect 32788 29484 35308 29540
rect 35364 29484 35374 29540
rect 9090 29372 9100 29428
rect 9156 29372 9884 29428
rect 9940 29372 9950 29428
rect 24098 29372 24108 29428
rect 24164 29372 27244 29428
rect 27300 29372 27310 29428
rect 39890 29372 39900 29428
rect 39956 29372 40572 29428
rect 40628 29372 40638 29428
rect 2034 29260 2044 29316
rect 2100 29260 5516 29316
rect 5572 29260 5582 29316
rect 17490 29260 17500 29316
rect 17556 29260 17948 29316
rect 18004 29260 19516 29316
rect 19572 29260 19582 29316
rect 25330 29260 25340 29316
rect 25396 29260 26124 29316
rect 26180 29260 27356 29316
rect 27412 29260 28140 29316
rect 28196 29260 28206 29316
rect 33506 29260 33516 29316
rect 33572 29260 33964 29316
rect 34020 29260 36540 29316
rect 36596 29260 36988 29316
rect 37044 29260 39788 29316
rect 39844 29260 40460 29316
rect 40516 29260 40526 29316
rect 21074 29036 21084 29092
rect 21140 29036 22316 29092
rect 22372 29036 22382 29092
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 1708 28980
rect 1764 28924 2492 28980
rect 2548 28924 2558 28980
rect 5842 28924 5852 28980
rect 5908 28924 6972 28980
rect 7028 28924 7038 28980
rect 0 28896 800 28924
rect 12562 28700 12572 28756
rect 12628 28700 13580 28756
rect 13636 28700 14140 28756
rect 14196 28700 14924 28756
rect 14980 28700 14990 28756
rect 18050 28700 18060 28756
rect 18116 28700 19852 28756
rect 19908 28700 19918 28756
rect 20514 28700 20524 28756
rect 20580 28700 22204 28756
rect 22260 28700 24388 28756
rect 24658 28700 24668 28756
rect 24724 28700 25620 28756
rect 28242 28700 28252 28756
rect 28308 28700 29036 28756
rect 29092 28700 29102 28756
rect 33394 28700 33404 28756
rect 33460 28700 35308 28756
rect 35364 28700 35374 28756
rect 24332 28644 24388 28700
rect 25564 28644 25620 28700
rect 9884 28588 11228 28644
rect 11284 28588 11294 28644
rect 19506 28588 19516 28644
rect 19572 28588 20636 28644
rect 20692 28588 20702 28644
rect 24322 28588 24332 28644
rect 24388 28588 25340 28644
rect 25396 28588 25406 28644
rect 25554 28588 25564 28644
rect 25620 28588 28028 28644
rect 28084 28588 28094 28644
rect 35074 28588 35084 28644
rect 35140 28588 36316 28644
rect 36372 28588 36382 28644
rect 9884 28420 9940 28588
rect 20132 28420 20188 28532
rect 20244 28476 20254 28532
rect 20850 28476 20860 28532
rect 20916 28476 23548 28532
rect 23604 28476 23614 28532
rect 29026 28476 29036 28532
rect 29092 28476 31500 28532
rect 31556 28476 31566 28532
rect 31892 28476 34300 28532
rect 34356 28476 34366 28532
rect 31892 28420 31948 28476
rect 9874 28364 9884 28420
rect 9940 28364 9950 28420
rect 16818 28364 16828 28420
rect 16884 28364 21196 28420
rect 21252 28364 21262 28420
rect 27794 28364 27804 28420
rect 27860 28364 31948 28420
rect 37650 28364 37660 28420
rect 37716 28364 39900 28420
rect 39956 28364 39966 28420
rect 0 28308 800 28336
rect 0 28252 1708 28308
rect 1764 28252 2492 28308
rect 2548 28252 2558 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 13906 28028 13916 28084
rect 13972 28028 18396 28084
rect 18452 28028 18462 28084
rect 2034 27916 2044 27972
rect 2100 27916 14476 27972
rect 14532 27916 14542 27972
rect 19730 27916 19740 27972
rect 19796 27916 25004 27972
rect 25060 27916 25070 27972
rect 16146 27804 16156 27860
rect 16212 27804 16604 27860
rect 16660 27804 20188 27860
rect 20244 27804 20254 27860
rect 0 27636 800 27664
rect 0 27580 1708 27636
rect 1764 27580 2492 27636
rect 2548 27580 2558 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 26450 27356 26460 27412
rect 26516 27356 30268 27412
rect 30324 27356 30334 27412
rect 6066 27132 6076 27188
rect 6132 27132 6860 27188
rect 6916 27132 6926 27188
rect 34626 27132 34636 27188
rect 34692 27132 37996 27188
rect 38052 27132 38062 27188
rect 6178 27020 6188 27076
rect 6244 27020 8652 27076
rect 8708 27020 8718 27076
rect 11218 27020 11228 27076
rect 11284 27020 12236 27076
rect 12292 27020 12302 27076
rect 14914 27020 14924 27076
rect 14980 27020 16156 27076
rect 16212 27020 16222 27076
rect 29698 27020 29708 27076
rect 29764 27020 30492 27076
rect 30548 27020 30558 27076
rect 0 26964 800 26992
rect 0 26908 2268 26964
rect 2324 26908 2334 26964
rect 5394 26908 5404 26964
rect 5460 26908 7868 26964
rect 7924 26908 7934 26964
rect 8372 26908 8876 26964
rect 8932 26908 10108 26964
rect 10164 26908 10174 26964
rect 17154 26908 17164 26964
rect 17220 26908 18284 26964
rect 18340 26908 26124 26964
rect 26180 26908 26908 26964
rect 26964 26908 26974 26964
rect 34402 26908 34412 26964
rect 34468 26908 35980 26964
rect 36036 26908 36046 26964
rect 0 26880 800 26908
rect 8372 26852 8428 26908
rect 7298 26796 7308 26852
rect 7364 26796 8428 26852
rect 9202 26796 9212 26852
rect 9268 26796 10556 26852
rect 10612 26796 10622 26852
rect 29810 26796 29820 26852
rect 29876 26796 30716 26852
rect 30772 26796 30782 26852
rect 8530 26684 8540 26740
rect 8596 26684 18396 26740
rect 18452 26684 18462 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 15586 26572 15596 26628
rect 15652 26572 15662 26628
rect 15596 26516 15652 26572
rect 8306 26460 8316 26516
rect 8372 26404 8428 26516
rect 15596 26460 20188 26516
rect 36866 26460 36876 26516
rect 36932 26460 38780 26516
rect 38836 26460 38846 26516
rect 8372 26348 9772 26404
rect 9828 26348 9838 26404
rect 16930 26348 16940 26404
rect 16996 26348 19404 26404
rect 19460 26348 19470 26404
rect 20132 26348 20188 26460
rect 20244 26348 20254 26404
rect 22418 26348 22428 26404
rect 22484 26348 23772 26404
rect 23828 26348 23838 26404
rect 0 26292 800 26320
rect 0 26236 2156 26292
rect 2212 26236 2222 26292
rect 27234 26236 27244 26292
rect 27300 26236 28364 26292
rect 28420 26236 33180 26292
rect 33236 26236 33246 26292
rect 0 26208 800 26236
rect 1810 26124 1820 26180
rect 1876 26124 3276 26180
rect 3332 26124 3342 26180
rect 19618 26124 19628 26180
rect 19684 26124 21084 26180
rect 21140 26124 23436 26180
rect 23492 26124 25340 26180
rect 25396 26124 26796 26180
rect 26852 26124 28924 26180
rect 28980 26124 28990 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 36978 25788 36988 25844
rect 37044 25788 38892 25844
rect 38948 25788 38958 25844
rect 39330 25676 39340 25732
rect 39396 25676 40796 25732
rect 40852 25676 40862 25732
rect 0 25620 800 25648
rect 0 25564 1820 25620
rect 1876 25564 1886 25620
rect 15474 25564 15484 25620
rect 15540 25564 16268 25620
rect 16324 25564 16604 25620
rect 16660 25564 20524 25620
rect 20580 25564 24892 25620
rect 24948 25564 27244 25620
rect 27300 25564 27310 25620
rect 0 25536 800 25564
rect 22978 25452 22988 25508
rect 23044 25452 23436 25508
rect 23492 25452 23502 25508
rect 36306 25452 36316 25508
rect 36372 25452 37100 25508
rect 37156 25452 37166 25508
rect 33618 25340 33628 25396
rect 33684 25340 34524 25396
rect 34580 25340 34590 25396
rect 22194 25228 22204 25284
rect 22260 25228 25676 25284
rect 25732 25228 25742 25284
rect 30146 25228 30156 25284
rect 30212 25228 32844 25284
rect 32900 25228 32910 25284
rect 33730 25116 33740 25172
rect 33796 25116 35644 25172
rect 35700 25116 36092 25172
rect 36148 25116 36158 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 0 24892 2156 24948
rect 2212 24892 2222 24948
rect 16370 24892 16380 24948
rect 16436 24892 17388 24948
rect 17444 24892 17454 24948
rect 31892 24892 33180 24948
rect 33236 24892 35084 24948
rect 35140 24892 38668 24948
rect 38724 24892 38734 24948
rect 0 24864 800 24892
rect 9538 24780 9548 24836
rect 9604 24780 10444 24836
rect 10500 24780 10892 24836
rect 10948 24780 10958 24836
rect 15810 24780 15820 24836
rect 15876 24780 17612 24836
rect 17668 24780 18284 24836
rect 18340 24780 18844 24836
rect 18900 24780 18910 24836
rect 2930 24668 2940 24724
rect 2996 24668 5628 24724
rect 5684 24668 5694 24724
rect 18844 24612 18900 24780
rect 31892 24724 31948 24892
rect 32722 24780 32732 24836
rect 32788 24780 35308 24836
rect 35364 24780 35374 24836
rect 20066 24668 20076 24724
rect 20132 24668 28868 24724
rect 30594 24668 30604 24724
rect 30660 24668 31724 24724
rect 31780 24668 31948 24724
rect 39106 24668 39116 24724
rect 39172 24668 39900 24724
rect 39956 24668 39966 24724
rect 28812 24612 28868 24668
rect 18844 24556 20412 24612
rect 20468 24556 20478 24612
rect 28802 24556 28812 24612
rect 28868 24556 28878 24612
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1932 24276
rect 1988 24220 1998 24276
rect 31266 24220 31276 24276
rect 31332 24220 34076 24276
rect 34132 24220 34142 24276
rect 0 24192 800 24220
rect 34290 24108 34300 24164
rect 34356 24108 37884 24164
rect 37940 24108 37950 24164
rect 21522 23996 21532 24052
rect 21588 23996 22316 24052
rect 22372 23996 22382 24052
rect 23426 23996 23436 24052
rect 23492 23996 25116 24052
rect 25172 23996 25182 24052
rect 35074 23996 35084 24052
rect 35140 23996 35756 24052
rect 35812 23996 35822 24052
rect 2034 23772 2044 23828
rect 2100 23772 4284 23828
rect 4340 23772 4350 23828
rect 4722 23772 4732 23828
rect 4788 23772 6188 23828
rect 6244 23772 6254 23828
rect 11890 23772 11900 23828
rect 11956 23772 12348 23828
rect 12404 23772 17052 23828
rect 17108 23772 17118 23828
rect 24546 23772 24556 23828
rect 24612 23772 26124 23828
rect 26180 23772 26190 23828
rect 8082 23660 8092 23716
rect 8148 23660 9436 23716
rect 9492 23660 9502 23716
rect 12786 23660 12796 23716
rect 12852 23660 15372 23716
rect 15428 23660 15438 23716
rect 18508 23660 19180 23716
rect 19236 23660 21420 23716
rect 21476 23660 21486 23716
rect 0 23604 800 23632
rect 18508 23604 18564 23660
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 11218 23548 11228 23604
rect 11284 23548 13356 23604
rect 13412 23548 13422 23604
rect 18396 23548 18564 23604
rect 33506 23548 33516 23604
rect 33572 23548 34972 23604
rect 35028 23548 35038 23604
rect 0 23520 800 23548
rect 18396 23492 18452 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 2034 23436 2044 23492
rect 2100 23436 3612 23492
rect 3668 23436 3678 23492
rect 15698 23436 15708 23492
rect 15764 23436 16492 23492
rect 16548 23436 17500 23492
rect 17556 23436 17836 23492
rect 17892 23436 18452 23492
rect 21410 23324 21420 23380
rect 21476 23324 26348 23380
rect 26404 23324 26414 23380
rect 12562 23212 12572 23268
rect 12628 23212 14588 23268
rect 14644 23212 14654 23268
rect 16258 23212 16268 23268
rect 16324 23212 18060 23268
rect 18116 23212 18126 23268
rect 20962 23212 20972 23268
rect 21028 23212 22316 23268
rect 22372 23212 22382 23268
rect 34962 23100 34972 23156
rect 35028 23100 36092 23156
rect 36148 23100 37100 23156
rect 37156 23100 40124 23156
rect 40180 23100 40190 23156
rect 0 22932 800 22960
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 14914 22876 14924 22932
rect 14980 22876 15932 22932
rect 15988 22876 16716 22932
rect 16772 22876 16782 22932
rect 0 22848 800 22876
rect 5282 22764 5292 22820
rect 5348 22764 7532 22820
rect 7588 22764 7598 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 35074 22540 35084 22596
rect 35140 22540 35150 22596
rect 37762 22540 37772 22596
rect 37828 22540 39900 22596
rect 39956 22540 39966 22596
rect 1698 22428 1708 22484
rect 1764 22428 2492 22484
rect 2548 22428 2558 22484
rect 8082 22428 8092 22484
rect 8148 22428 13804 22484
rect 13860 22428 13870 22484
rect 14242 22428 14252 22484
rect 14308 22428 16828 22484
rect 16884 22428 16894 22484
rect 15250 22316 15260 22372
rect 15316 22316 18732 22372
rect 18788 22316 18798 22372
rect 20402 22316 20412 22372
rect 20468 22316 21644 22372
rect 21700 22316 22204 22372
rect 22260 22316 22270 22372
rect 29250 22316 29260 22372
rect 29316 22316 30940 22372
rect 30996 22316 32284 22372
rect 32340 22316 32350 22372
rect 0 22260 800 22288
rect 35084 22260 35140 22540
rect 40002 22428 40012 22484
rect 40068 22428 41020 22484
rect 41076 22428 41086 22484
rect 0 22204 4844 22260
rect 4900 22204 4910 22260
rect 7074 22204 7084 22260
rect 7140 22204 11788 22260
rect 11844 22204 11854 22260
rect 12450 22204 12460 22260
rect 12516 22204 13916 22260
rect 13972 22204 13982 22260
rect 14242 22204 14252 22260
rect 14308 22204 14924 22260
rect 14980 22204 14990 22260
rect 26338 22204 26348 22260
rect 26404 22204 35140 22260
rect 38994 22204 39004 22260
rect 39060 22204 39070 22260
rect 0 22176 800 22204
rect 8194 22092 8204 22148
rect 8260 22092 10668 22148
rect 10724 22092 10734 22148
rect 13010 22092 13020 22148
rect 13076 22092 13086 22148
rect 28242 22092 28252 22148
rect 28308 22092 29596 22148
rect 29652 22092 29662 22148
rect 13020 22036 13076 22092
rect 39004 22036 39060 22204
rect 6962 21980 6972 22036
rect 7028 21980 13076 22036
rect 29026 21980 29036 22036
rect 29092 21980 39060 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 6748 21868 9548 21924
rect 9604 21868 10668 21924
rect 10724 21868 10734 21924
rect 36754 21868 36764 21924
rect 36820 21868 38220 21924
rect 38276 21868 38286 21924
rect 2370 21644 2380 21700
rect 2436 21644 3500 21700
rect 3556 21644 3566 21700
rect 6748 21588 6804 21868
rect 32050 21756 32060 21812
rect 32116 21756 33180 21812
rect 33236 21756 33246 21812
rect 37426 21756 37436 21812
rect 37492 21756 38444 21812
rect 38500 21756 38510 21812
rect 7970 21644 7980 21700
rect 8036 21644 8428 21700
rect 8372 21588 8428 21644
rect 25788 21644 34076 21700
rect 34132 21644 34142 21700
rect 25788 21588 25844 21644
rect 1810 21532 1820 21588
rect 1876 21532 5628 21588
rect 5684 21532 6748 21588
rect 6804 21532 6814 21588
rect 8372 21532 12460 21588
rect 12516 21532 12526 21588
rect 24434 21532 24444 21588
rect 24500 21532 25116 21588
rect 25172 21532 25182 21588
rect 25778 21532 25788 21588
rect 25844 21532 25854 21588
rect 29586 21532 29596 21588
rect 29652 21532 37996 21588
rect 38052 21532 38062 21588
rect 38658 21532 38668 21588
rect 38724 21532 39788 21588
rect 39844 21532 39854 21588
rect 38668 21476 38724 21532
rect 7970 21420 7980 21476
rect 8036 21420 8428 21476
rect 15026 21420 15036 21476
rect 15092 21420 18732 21476
rect 18788 21420 18798 21476
rect 37762 21420 37772 21476
rect 37828 21420 38724 21476
rect 8372 21364 8428 21420
rect 8372 21308 13804 21364
rect 13860 21308 13870 21364
rect 16930 21308 16940 21364
rect 16996 21308 17948 21364
rect 18004 21308 18014 21364
rect 32610 21308 32620 21364
rect 32676 21308 39004 21364
rect 39060 21308 39070 21364
rect 32162 21196 32172 21252
rect 32228 21196 33964 21252
rect 34020 21196 34030 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 20626 21084 20636 21140
rect 20692 21084 24108 21140
rect 24164 21084 24174 21140
rect 0 20916 800 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 18274 20860 18284 20916
rect 18340 20860 19068 20916
rect 19124 20860 19134 20916
rect 23874 20860 23884 20916
rect 23940 20860 24892 20916
rect 24948 20860 24958 20916
rect 35186 20860 35196 20916
rect 35252 20860 37212 20916
rect 37268 20860 37278 20916
rect 37986 20860 37996 20916
rect 38052 20860 38062 20916
rect 0 20832 800 20860
rect 37996 20804 38052 20860
rect 4834 20748 4844 20804
rect 4900 20748 20860 20804
rect 20916 20748 20926 20804
rect 31378 20748 31388 20804
rect 31444 20748 38052 20804
rect 1586 20636 1596 20692
rect 1652 20636 2716 20692
rect 2772 20636 2782 20692
rect 21186 20524 21196 20580
rect 21252 20524 24444 20580
rect 24500 20524 27020 20580
rect 27076 20524 27086 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 3378 20300 3388 20356
rect 3444 20300 4060 20356
rect 4116 20300 6188 20356
rect 6244 20300 6254 20356
rect 13570 20188 13580 20244
rect 13636 20188 17388 20244
rect 17444 20188 17454 20244
rect 37202 20188 37212 20244
rect 37268 20188 38556 20244
rect 38612 20188 38622 20244
rect 7746 20076 7756 20132
rect 7812 20076 9660 20132
rect 9716 20076 9726 20132
rect 30930 20076 30940 20132
rect 30996 20076 32620 20132
rect 32676 20076 32686 20132
rect 32498 19964 32508 20020
rect 32564 19964 33516 20020
rect 33572 19964 33582 20020
rect 35074 19964 35084 20020
rect 35140 19964 37884 20020
rect 37940 19964 37950 20020
rect 15250 19852 15260 19908
rect 15316 19852 17164 19908
rect 17220 19852 17230 19908
rect 19058 19740 19068 19796
rect 19124 19740 20076 19796
rect 20132 19740 20412 19796
rect 20468 19740 25676 19796
rect 25732 19740 27020 19796
rect 27076 19740 27086 19796
rect 30818 19740 30828 19796
rect 30884 19740 39004 19796
rect 39060 19740 39070 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 37986 19516 37996 19572
rect 38052 19516 39564 19572
rect 39620 19516 39630 19572
rect 4050 19292 4060 19348
rect 4116 19292 8092 19348
rect 8148 19292 8158 19348
rect 23986 19292 23996 19348
rect 24052 19292 26124 19348
rect 26180 19292 26190 19348
rect 32162 19292 32172 19348
rect 32228 19292 37996 19348
rect 38052 19292 38062 19348
rect 20738 19180 20748 19236
rect 20804 19180 21756 19236
rect 21812 19180 21822 19236
rect 24882 19068 24892 19124
rect 24948 19068 27132 19124
rect 27188 19068 27198 19124
rect 28802 19068 28812 19124
rect 28868 19068 34972 19124
rect 35028 19068 35038 19124
rect 7074 18956 7084 19012
rect 7140 18956 8764 19012
rect 8820 18956 8830 19012
rect 17154 18956 17164 19012
rect 17220 18956 19516 19012
rect 19572 18956 19582 19012
rect 23762 18956 23772 19012
rect 23828 18956 25788 19012
rect 25844 18956 25854 19012
rect 3826 18844 3836 18900
rect 3892 18844 6076 18900
rect 6132 18844 6142 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 24546 18508 24556 18564
rect 24612 18508 29036 18564
rect 29092 18508 29102 18564
rect 7522 18396 7532 18452
rect 7588 18396 8428 18452
rect 11330 18396 11340 18452
rect 11396 18396 15596 18452
rect 15652 18396 15662 18452
rect 17826 18396 17836 18452
rect 17892 18396 18508 18452
rect 18564 18396 18574 18452
rect 25778 18396 25788 18452
rect 25844 18396 30716 18452
rect 30772 18396 33516 18452
rect 33572 18396 33582 18452
rect 35858 18396 35868 18452
rect 35924 18396 38780 18452
rect 38836 18396 38846 18452
rect 8372 18340 8428 18396
rect 8372 18284 8988 18340
rect 9044 18284 11900 18340
rect 11956 18284 11966 18340
rect 20290 18284 20300 18340
rect 20356 18284 23212 18340
rect 23268 18284 23278 18340
rect 32610 18284 32620 18340
rect 32676 18284 35308 18340
rect 35364 18284 36204 18340
rect 36260 18284 36270 18340
rect 8866 18172 8876 18228
rect 8932 18172 12572 18228
rect 12628 18172 12638 18228
rect 20748 18172 21756 18228
rect 21812 18172 22876 18228
rect 22932 18172 24108 18228
rect 24164 18172 26796 18228
rect 26852 18172 28588 18228
rect 28644 18172 28654 18228
rect 20748 18116 20804 18172
rect 20738 18060 20748 18116
rect 20804 18060 20814 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 10322 17836 10332 17892
rect 10388 17836 13020 17892
rect 13076 17836 13086 17892
rect 13234 17836 13244 17892
rect 13300 17836 14028 17892
rect 14084 17836 14094 17892
rect 8082 17724 8092 17780
rect 8148 17724 8428 17780
rect 20066 17724 20076 17780
rect 20132 17724 20748 17780
rect 20804 17724 20814 17780
rect 32498 17724 32508 17780
rect 32564 17724 33628 17780
rect 33684 17724 34636 17780
rect 34692 17724 35420 17780
rect 35476 17724 35486 17780
rect 8372 17668 8428 17724
rect 2370 17612 2380 17668
rect 2436 17612 3388 17668
rect 3444 17612 4732 17668
rect 4788 17612 7532 17668
rect 7588 17612 7598 17668
rect 8372 17612 9884 17668
rect 9940 17612 9950 17668
rect 32386 17612 32396 17668
rect 32452 17612 35084 17668
rect 35140 17612 35150 17668
rect 38658 17612 38668 17668
rect 38724 17612 39788 17668
rect 39844 17612 41020 17668
rect 41076 17612 41086 17668
rect 36530 17500 36540 17556
rect 36596 17500 39004 17556
rect 39060 17500 39070 17556
rect 26338 17388 26348 17444
rect 26404 17388 26908 17444
rect 26964 17388 27580 17444
rect 27636 17388 27646 17444
rect 37874 17388 37884 17444
rect 37940 17388 39900 17444
rect 39956 17388 39966 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 17042 17164 17052 17220
rect 17108 17164 19180 17220
rect 19236 17164 19246 17220
rect 5618 17052 5628 17108
rect 5684 17052 6300 17108
rect 6356 17052 6366 17108
rect 27794 17052 27804 17108
rect 27860 17052 30044 17108
rect 30100 17052 30110 17108
rect 9538 16940 9548 16996
rect 9604 16940 10556 16996
rect 10612 16940 12796 16996
rect 12852 16940 13580 16996
rect 13636 16940 13646 16996
rect 28802 16940 28812 16996
rect 28868 16940 31052 16996
rect 31108 16940 31118 16996
rect 35522 16940 35532 16996
rect 35588 16940 36428 16996
rect 36484 16940 38668 16996
rect 38724 16940 38734 16996
rect 16594 16828 16604 16884
rect 16660 16828 17948 16884
rect 18004 16828 18396 16884
rect 18452 16828 18956 16884
rect 19012 16828 19404 16884
rect 19460 16828 20860 16884
rect 20916 16828 20926 16884
rect 25330 16828 25340 16884
rect 25396 16828 26124 16884
rect 26180 16828 27244 16884
rect 27300 16828 27310 16884
rect 36194 16828 36204 16884
rect 36260 16828 37212 16884
rect 37268 16828 37660 16884
rect 37716 16828 37726 16884
rect 38098 16828 38108 16884
rect 38164 16828 38892 16884
rect 38948 16828 38958 16884
rect 25340 16772 25396 16828
rect 4722 16716 4732 16772
rect 4788 16716 7532 16772
rect 7588 16716 7598 16772
rect 23538 16716 23548 16772
rect 23604 16716 24220 16772
rect 24276 16716 25396 16772
rect 31490 16716 31500 16772
rect 31556 16716 32620 16772
rect 32676 16716 33180 16772
rect 33236 16716 33246 16772
rect 22866 16604 22876 16660
rect 22932 16604 25452 16660
rect 25508 16604 25518 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 4946 16380 4956 16436
rect 5012 16380 7420 16436
rect 7476 16380 7486 16436
rect 12450 16268 12460 16324
rect 12516 16268 13580 16324
rect 13636 16268 13646 16324
rect 3938 16044 3948 16100
rect 4004 16044 8540 16100
rect 8596 16044 8606 16100
rect 3042 15932 3052 15988
rect 3108 15932 5516 15988
rect 5572 15932 5582 15988
rect 16146 15820 16156 15876
rect 16212 15820 20524 15876
rect 20580 15820 23772 15876
rect 23828 15820 23838 15876
rect 27010 15820 27020 15876
rect 27076 15820 28700 15876
rect 28756 15820 28766 15876
rect 34402 15820 34412 15876
rect 34468 15820 35308 15876
rect 35364 15820 35374 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23986 15596 23996 15652
rect 24052 15596 30716 15652
rect 30772 15596 30782 15652
rect 13234 15484 13244 15540
rect 13300 15484 13804 15540
rect 13860 15484 13870 15540
rect 4050 15260 4060 15316
rect 4116 15260 5068 15316
rect 5124 15260 5134 15316
rect 27234 15260 27244 15316
rect 27300 15260 27692 15316
rect 27748 15260 28588 15316
rect 28644 15260 29932 15316
rect 29988 15260 29998 15316
rect 20514 15148 20524 15204
rect 20580 15148 23548 15204
rect 23604 15148 23614 15204
rect 25778 15148 25788 15204
rect 25844 15148 27580 15204
rect 27636 15148 27646 15204
rect 36306 15148 36316 15204
rect 36372 15148 37100 15204
rect 37156 15148 37166 15204
rect 16706 15036 16716 15092
rect 16772 15036 18508 15092
rect 18564 15036 18574 15092
rect 40450 15036 40460 15092
rect 40516 15036 41468 15092
rect 41524 15036 41534 15092
rect 13682 14924 13692 14980
rect 13748 14924 18396 14980
rect 18452 14924 18462 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 21298 14812 21308 14868
rect 21364 14812 22316 14868
rect 22372 14812 22382 14868
rect 6402 14588 6412 14644
rect 6468 14588 8540 14644
rect 8596 14588 9548 14644
rect 9604 14588 10444 14644
rect 10500 14588 10510 14644
rect 15810 14588 15820 14644
rect 15876 14588 17500 14644
rect 17556 14588 18284 14644
rect 18340 14588 20748 14644
rect 20804 14588 21420 14644
rect 21476 14588 21486 14644
rect 31938 14588 31948 14644
rect 32004 14588 34972 14644
rect 35028 14588 35038 14644
rect 16818 14476 16828 14532
rect 16884 14476 20300 14532
rect 20356 14476 21644 14532
rect 21700 14476 22204 14532
rect 22260 14476 22270 14532
rect 1586 14364 1596 14420
rect 1652 14364 2716 14420
rect 2772 14364 2782 14420
rect 10098 14364 10108 14420
rect 10164 14364 12348 14420
rect 12404 14364 12414 14420
rect 29810 14364 29820 14420
rect 29876 14364 30940 14420
rect 30996 14364 31006 14420
rect 29474 14252 29484 14308
rect 29540 14252 32844 14308
rect 32900 14252 32910 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 23202 13804 23212 13860
rect 23268 13804 23996 13860
rect 24052 13804 24062 13860
rect 27346 13804 27356 13860
rect 27412 13804 32060 13860
rect 32116 13804 32126 13860
rect 33282 13804 33292 13860
rect 33348 13804 35868 13860
rect 35924 13804 35934 13860
rect 3378 13692 3388 13748
rect 3444 13692 4620 13748
rect 4676 13692 4686 13748
rect 23762 13692 23772 13748
rect 23828 13692 26124 13748
rect 26180 13692 28588 13748
rect 28644 13692 28654 13748
rect 28242 13580 28252 13636
rect 28308 13580 31052 13636
rect 31108 13580 31118 13636
rect 4162 13468 4172 13524
rect 4228 13468 6076 13524
rect 6132 13468 6142 13524
rect 36978 13468 36988 13524
rect 37044 13468 38108 13524
rect 38164 13468 40348 13524
rect 40404 13468 40414 13524
rect 37090 13356 37100 13412
rect 37156 13356 39340 13412
rect 39396 13356 39406 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 38322 13244 38332 13300
rect 38388 13244 40348 13300
rect 40404 13244 40414 13300
rect 9314 13132 9324 13188
rect 9380 13132 10668 13188
rect 10724 13132 10734 13188
rect 24770 13132 24780 13188
rect 24836 13132 26908 13188
rect 26964 13132 26974 13188
rect 32050 13020 32060 13076
rect 32116 13020 33964 13076
rect 34020 13020 34030 13076
rect 6962 12908 6972 12964
rect 7028 12908 8540 12964
rect 8596 12908 9884 12964
rect 9940 12908 9950 12964
rect 11778 12908 11788 12964
rect 11844 12908 12460 12964
rect 12516 12908 13468 12964
rect 13524 12908 13534 12964
rect 17938 12908 17948 12964
rect 18004 12908 18732 12964
rect 18788 12908 18798 12964
rect 21634 12908 21644 12964
rect 21700 12908 22540 12964
rect 22596 12908 22606 12964
rect 29250 12908 29260 12964
rect 29316 12908 30044 12964
rect 30100 12908 30110 12964
rect 39218 12908 39228 12964
rect 39284 12908 39788 12964
rect 39844 12908 40124 12964
rect 40180 12908 40190 12964
rect 32722 12796 32732 12852
rect 32788 12796 34972 12852
rect 35028 12796 35038 12852
rect 6850 12684 6860 12740
rect 6916 12684 7756 12740
rect 7812 12684 7822 12740
rect 9762 12684 9772 12740
rect 9828 12684 10668 12740
rect 10724 12684 11228 12740
rect 11284 12684 11294 12740
rect 26786 12684 26796 12740
rect 26852 12684 27692 12740
rect 27748 12684 27758 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 10098 12348 10108 12404
rect 10164 12348 12236 12404
rect 12292 12348 12302 12404
rect 9874 12124 9884 12180
rect 9940 12124 10444 12180
rect 10500 12124 11788 12180
rect 11844 12124 11854 12180
rect 16594 12124 16604 12180
rect 16660 12124 17500 12180
rect 17556 12124 17566 12180
rect 30034 12124 30044 12180
rect 30100 12124 32620 12180
rect 32676 12124 33068 12180
rect 33124 12124 34076 12180
rect 34132 12124 34142 12180
rect 36642 12012 36652 12068
rect 36708 12012 37884 12068
rect 37940 12012 37950 12068
rect 38668 11788 39228 11844
rect 39284 11788 39294 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 38668 11732 38724 11788
rect 36530 11676 36540 11732
rect 36596 11676 36988 11732
rect 37044 11676 38444 11732
rect 38500 11676 38724 11732
rect 25890 11564 25900 11620
rect 25956 11564 27580 11620
rect 27636 11564 27646 11620
rect 6066 11452 6076 11508
rect 6132 11452 7644 11508
rect 7700 11452 7710 11508
rect 24322 11452 24332 11508
rect 24388 11452 25676 11508
rect 25732 11452 25742 11508
rect 39890 11452 39900 11508
rect 39956 11452 40684 11508
rect 40740 11452 40750 11508
rect 16482 11340 16492 11396
rect 16548 11340 17948 11396
rect 18004 11340 18620 11396
rect 18676 11340 20076 11396
rect 20132 11340 20142 11396
rect 7186 11228 7196 11284
rect 7252 11228 8652 11284
rect 8708 11228 8718 11284
rect 13570 11116 13580 11172
rect 13636 11116 14588 11172
rect 14644 11116 14654 11172
rect 16594 11116 16604 11172
rect 16660 11116 21980 11172
rect 22036 11116 22046 11172
rect 33730 11116 33740 11172
rect 33796 11116 34972 11172
rect 35028 11116 35038 11172
rect 23538 11004 23548 11060
rect 23604 11004 24332 11060
rect 24388 11004 24398 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 15026 10780 15036 10836
rect 15092 10780 16492 10836
rect 16548 10780 16558 10836
rect 21186 10780 21196 10836
rect 21252 10780 22652 10836
rect 22708 10780 22718 10836
rect 37762 10780 37772 10836
rect 37828 10780 39116 10836
rect 39172 10780 39182 10836
rect 9090 10668 9100 10724
rect 9156 10668 11564 10724
rect 11620 10668 11630 10724
rect 14354 10668 14364 10724
rect 14420 10668 15372 10724
rect 15428 10668 15438 10724
rect 25106 10668 25116 10724
rect 25172 10668 26236 10724
rect 26292 10668 26302 10724
rect 30146 10668 30156 10724
rect 30212 10668 32172 10724
rect 32228 10668 32238 10724
rect 17714 10556 17724 10612
rect 17780 10556 22540 10612
rect 22596 10556 22606 10612
rect 34738 10444 34748 10500
rect 34804 10444 36876 10500
rect 36932 10444 36942 10500
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 12450 9996 12460 10052
rect 12516 9996 15372 10052
rect 15428 9996 15438 10052
rect 19506 9996 19516 10052
rect 19572 9996 20972 10052
rect 21028 9996 21038 10052
rect 8194 9772 8204 9828
rect 8260 9772 9548 9828
rect 9604 9772 9614 9828
rect 27570 9772 27580 9828
rect 27636 9772 28028 9828
rect 28084 9772 28588 9828
rect 28644 9772 29484 9828
rect 29540 9772 30492 9828
rect 30548 9772 32060 9828
rect 32116 9772 32126 9828
rect 2034 9660 2044 9716
rect 2100 9660 2110 9716
rect 0 9492 800 9520
rect 2044 9492 2100 9660
rect 0 9436 2100 9492
rect 8642 9436 8652 9492
rect 8708 9436 10556 9492
rect 10612 9436 10622 9492
rect 0 9408 800 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 9986 9324 9996 9380
rect 10052 9324 12012 9380
rect 12068 9324 12078 9380
rect 16146 9324 16156 9380
rect 16212 9324 17276 9380
rect 17332 9324 17342 9380
rect 11666 9100 11676 9156
rect 11732 9100 13020 9156
rect 13076 9100 13086 9156
rect 16706 9100 16716 9156
rect 16772 9100 20412 9156
rect 20468 9100 20478 9156
rect 1922 8876 1932 8932
rect 1988 8876 1998 8932
rect 9538 8876 9548 8932
rect 9604 8876 12124 8932
rect 12180 8876 13916 8932
rect 13972 8876 13982 8932
rect 0 8820 800 8848
rect 1932 8820 1988 8876
rect 0 8764 1988 8820
rect 0 8736 800 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 0 8148 800 8176
rect 0 8092 2044 8148
rect 2100 8092 2110 8148
rect 0 8064 800 8092
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 13122 7532 13132 7588
rect 13188 7532 14252 7588
rect 14308 7532 14318 7588
rect 0 7476 800 7504
rect 0 7420 3276 7476
rect 3332 7420 3342 7476
rect 0 7392 800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 0 6804 800 6832
rect 0 6748 1932 6804
rect 1988 6748 1998 6804
rect 0 6720 800 6748
rect 2706 6524 2716 6580
rect 2772 6524 4284 6580
rect 4340 6524 4350 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 0 6132 800 6160
rect 0 6076 2044 6132
rect 2100 6076 2110 6132
rect 0 6048 800 6076
rect 0 5460 800 5488
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 0 5404 1932 5460
rect 1988 5404 1998 5460
rect 0 5376 800 5404
rect 2706 5180 2716 5236
rect 2772 5180 3836 5236
rect 3892 5180 3902 5236
rect 2034 5068 2044 5124
rect 2100 5068 4508 5124
rect 4564 5068 4574 5124
rect 3266 4956 3276 5012
rect 3332 4956 3724 5012
rect 3780 4956 3790 5012
rect 0 4788 800 4816
rect 0 4732 980 4788
rect 0 4704 800 4732
rect 924 4564 980 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 924 4508 1764 4564
rect 3266 4508 3276 4564
rect 3332 4508 3612 4564
rect 3668 4508 3678 4564
rect 1708 4452 1764 4508
rect 1698 4396 1708 4452
rect 1764 4396 4844 4452
rect 4900 4396 4910 4452
rect 1698 4172 1708 4228
rect 1764 4172 5740 4228
rect 5796 4172 5806 4228
rect 0 4116 800 4144
rect 0 4060 2380 4116
rect 2436 4060 2446 4116
rect 0 4032 800 4060
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 1698 3500 1708 3556
rect 1764 3500 1774 3556
rect 2370 3500 2380 3556
rect 2436 3500 5292 3556
rect 5348 3500 5358 3556
rect 0 3444 800 3472
rect 1708 3444 1764 3500
rect 0 3388 1764 3444
rect 3042 3388 3052 3444
rect 3108 3388 4956 3444
rect 5012 3388 5022 3444
rect 0 3360 800 3388
rect 8082 3276 8092 3332
rect 8148 3276 9324 3332
rect 9380 3276 9390 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 2772 800 2800
rect 0 2716 3948 2772
rect 4004 2716 4014 2772
rect 0 2688 800 2716
rect 0 2100 800 2128
rect 0 2044 3836 2100
rect 3892 2044 3902 2100
rect 0 2016 800 2044
rect 1810 1708 1820 1764
rect 1876 1708 1886 1764
rect 0 1428 800 1456
rect 1820 1428 1876 1708
rect 0 1372 1876 1428
rect 0 1344 800 1372
rect 0 756 800 784
rect 0 700 2380 756
rect 2436 700 2446 756
rect 0 672 800 700
rect 0 84 800 112
rect 0 28 2940 84
rect 2996 28 3006 84
rect 0 0 800 28
<< via3 >>
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 5628 37772 5684 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 3612 37212 3668 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 5628 24668 5684 24724
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 3612 23436 3668 23492
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 40012 4768 40828
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 3612 37268 3668 37278
rect 3612 23492 3668 37212
rect 3612 23426 3668 23436
rect 4448 36876 4768 38388
rect 19808 40796 20128 40828
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 5628 37828 5684 37838
rect 5628 24724 5684 37772
rect 5628 24658 5684 24668
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 40012 35488 40828
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14336 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _127_
timestamp 1698431365
transform -1 0 15008 0 -1 20384
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8064 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _129_
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _130_
timestamp 1698431365
transform 1 0 3920 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _131_
timestamp 1698431365
transform -1 0 6720 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _132_
timestamp 1698431365
transform 1 0 3024 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _133_
timestamp 1698431365
transform -1 0 3920 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _134_
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _135_
timestamp 1698431365
transform -1 0 4480 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _136_
timestamp 1698431365
transform 1 0 1904 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _137_
timestamp 1698431365
transform 1 0 1904 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _138_
timestamp 1698431365
transform -1 0 15344 0 -1 15680
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _139_
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _140_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _141_
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _142_
timestamp 1698431365
transform -1 0 11984 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _143_
timestamp 1698431365
transform -1 0 10640 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _144_
timestamp 1698431365
transform 1 0 8064 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _145_
timestamp 1698431365
transform -1 0 7168 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _146_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _147_
timestamp 1698431365
transform 1 0 13440 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _148_
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _149_
timestamp 1698431365
transform -1 0 20496 0 1 17248
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _150_
timestamp 1698431365
transform 1 0 22400 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _151_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _152_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _153_
timestamp 1698431365
transform -1 0 18368 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _154_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _155_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _156_
timestamp 1698431365
transform -1 0 22288 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _157_
timestamp 1698431365
transform -1 0 20496 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _158_
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _159_
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _160_
timestamp 1698431365
transform 1 0 23072 0 1 17248
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _161_
timestamp 1698431365
transform 1 0 27328 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _162_
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _163_
timestamp 1698431365
transform -1 0 30688 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _164_
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _165_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _166_
timestamp 1698431365
transform 1 0 32592 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _167_
timestamp 1698431365
transform -1 0 28000 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _168_
timestamp 1698431365
transform -1 0 26544 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _169_
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _170_
timestamp 1698431365
transform -1 0 30128 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _171_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _172_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _173_
timestamp 1698431365
transform -1 0 34048 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _174_
timestamp 1698431365
transform -1 0 39648 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _175_
timestamp 1698431365
transform 1 0 39984 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _176_
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _177_
timestamp 1698431365
transform 1 0 39648 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _178_
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _179_
timestamp 1698431365
transform -1 0 35952 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _180_
timestamp 1698431365
transform -1 0 34048 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _181_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _182_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _183_
timestamp 1698431365
transform 1 0 27552 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _184_
timestamp 1698431365
transform -1 0 27552 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _185_
timestamp 1698431365
transform -1 0 26208 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _186_
timestamp 1698431365
transform 1 0 21504 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _187_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _188_
timestamp 1698431365
transform -1 0 19264 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _189_
timestamp 1698431365
transform 1 0 25648 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _190_
timestamp 1698431365
transform -1 0 26208 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _191_
timestamp 1698431365
transform -1 0 22736 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _192_
timestamp 1698431365
transform -1 0 22288 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _193_
timestamp 1698431365
transform 1 0 27104 0 -1 23520
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _194_
timestamp 1698431365
transform -1 0 35280 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _195_
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _196_
timestamp 1698431365
transform 1 0 31584 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _197_
timestamp 1698431365
transform 1 0 30464 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _198_
timestamp 1698431365
transform 1 0 38528 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _199_
timestamp 1698431365
transform -1 0 39648 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _200_
timestamp 1698431365
transform 1 0 39648 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _201_
timestamp 1698431365
transform 1 0 39312 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _202_
timestamp 1698431365
transform 1 0 38192 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _203_
timestamp 1698431365
transform -1 0 35504 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _204_
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _205_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _206_
timestamp 1698431365
transform -1 0 36400 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _207_
timestamp 1698431365
transform -1 0 34048 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _208_
timestamp 1698431365
transform 1 0 40768 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _209_
timestamp 1698431365
transform -1 0 39648 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _210_
timestamp 1698431365
transform 1 0 39648 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _211_
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _212_
timestamp 1698431365
transform -1 0 31696 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _213_
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _214_
timestamp 1698431365
transform -1 0 28784 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _215_
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _216_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _217_
timestamp 1698431365
transform -1 0 24864 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _218_
timestamp 1698431365
transform 1 0 27888 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _219_
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _220_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _221_
timestamp 1698431365
transform -1 0 22064 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _222_
timestamp 1698431365
transform -1 0 20384 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _223_
timestamp 1698431365
transform -1 0 20608 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _224_
timestamp 1698431365
transform -1 0 19936 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _225_
timestamp 1698431365
transform -1 0 17024 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _226_
timestamp 1698431365
transform -1 0 15120 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _227_
timestamp 1698431365
transform 1 0 14784 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _228_
timestamp 1698431365
transform -1 0 12880 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _229_
timestamp 1698431365
transform -1 0 10304 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _230_
timestamp 1698431365
transform -1 0 9184 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _231_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _232_
timestamp 1698431365
transform -1 0 10640 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _233_
timestamp 1698431365
transform -1 0 11312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _234_
timestamp 1698431365
transform -1 0 11984 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _235_
timestamp 1698431365
transform -1 0 10640 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _236_
timestamp 1698431365
transform -1 0 7504 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _237_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _238_
timestamp 1698431365
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _239_
timestamp 1698431365
transform 1 0 15792 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _240_
timestamp 1698431365
transform -1 0 15120 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _241_
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _242_
timestamp 1698431365
transform -1 0 17920 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _243_
timestamp 1698431365
transform -1 0 20720 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _244_
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _245_
timestamp 1698431365
transform -1 0 18592 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _246_
timestamp 1698431365
transform 1 0 15680 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _247_
timestamp 1698431365
transform -1 0 14448 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _248_
timestamp 1698431365
transform -1 0 12096 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _249_
timestamp 1698431365
transform -1 0 11200 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _250_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6720 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _251_
timestamp 1698431365
transform -1 0 12544 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _252_
timestamp 1698431365
transform -1 0 6832 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _253_
timestamp 1698431365
transform -1 0 8848 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _254_
timestamp 1698431365
transform -1 0 5376 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _255_
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _256_
timestamp 1698431365
transform 1 0 4480 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _257_
timestamp 1698431365
transform -1 0 9296 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _258_
timestamp 1698431365
transform -1 0 5376 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _259_
timestamp 1698431365
transform -1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _260_
timestamp 1698431365
transform -1 0 16352 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _261_
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _262_
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _263_
timestamp 1698431365
transform 1 0 9296 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _264_
timestamp 1698431365
transform 1 0 7952 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _265_
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _266_
timestamp 1698431365
transform -1 0 10976 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _267_
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _268_
timestamp 1698431365
transform 1 0 11984 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _269_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _270_
timestamp 1698431365
transform -1 0 24192 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _271_
timestamp 1698431365
transform 1 0 18592 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _272_
timestamp 1698431365
transform -1 0 20384 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _273_
timestamp 1698431365
transform 1 0 14784 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _274_
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _275_
timestamp 1698431365
transform 1 0 13216 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _276_
timestamp 1698431365
transform 1 0 19152 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _277_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _278_
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _279_
timestamp 1698431365
transform -1 0 24304 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _280_
timestamp 1698431365
transform -1 0 28896 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _281_
timestamp 1698431365
transform 1 0 23632 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _282_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _283_
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _284_
timestamp 1698431365
transform 1 0 30016 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _285_
timestamp 1698431365
transform -1 0 32704 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _286_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _287_
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _288_
timestamp 1698431365
transform -1 0 32816 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _289_
timestamp 1698431365
transform 1 0 27104 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _290_
timestamp 1698431365
transform 1 0 34048 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _291_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _292_
timestamp 1698431365
transform 1 0 36736 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _293_
timestamp 1698431365
transform -1 0 40656 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _294_
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _295_
timestamp 1698431365
transform -1 0 40880 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _296_
timestamp 1698431365
transform -1 0 38864 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _297_
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _298_
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _299_
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _300_
timestamp 1698431365
transform -1 0 32816 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _301_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _302_
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _303_
timestamp 1698431365
transform -1 0 24752 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _304_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _305_
timestamp 1698431365
transform -1 0 20944 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _306_
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _307_
timestamp 1698431365
transform 1 0 22736 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _308_
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _309_
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _310_
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _311_
timestamp 1698431365
transform 1 0 30576 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _312_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _313_
timestamp 1698431365
transform -1 0 32816 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _314_
timestamp 1698431365
transform 1 0 33936 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _315_
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _316_
timestamp 1698431365
transform -1 0 40768 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _317_
timestamp 1698431365
transform 1 0 36064 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _318_
timestamp 1698431365
transform 1 0 34384 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _319_
timestamp 1698431365
transform 1 0 32816 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _320_
timestamp 1698431365
transform -1 0 38192 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _321_
timestamp 1698431365
transform 1 0 32816 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _322_
timestamp 1698431365
transform -1 0 36736 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _323_
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _324_
timestamp 1698431365
transform 1 0 36960 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _325_
timestamp 1698431365
transform -1 0 40656 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _326_
timestamp 1698431365
transform -1 0 34048 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _327_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _328_
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _329_
timestamp 1698431365
transform 1 0 25648 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _330_
timestamp 1698431365
transform 1 0 23296 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _331_
timestamp 1698431365
transform 1 0 21056 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _332_
timestamp 1698431365
transform 1 0 24080 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _333_
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _334_
timestamp 1698431365
transform 1 0 20384 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _335_
timestamp 1698431365
transform 1 0 17136 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _336_
timestamp 1698431365
transform -1 0 21056 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _337_
timestamp 1698431365
transform 1 0 15456 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _338_
timestamp 1698431365
transform -1 0 19712 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _339_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _340_
timestamp 1698431365
transform 1 0 11536 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _341_
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _342_
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _343_
timestamp 1698431365
transform -1 0 9184 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _344_
timestamp 1698431365
transform 1 0 10640 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _345_
timestamp 1698431365
transform -1 0 12992 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _346_
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _347_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _348_
timestamp 1698431365
transform 1 0 5376 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _349_
timestamp 1698431365
transform -1 0 8736 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _350_
timestamp 1698431365
transform -1 0 19488 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _351_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _352_
timestamp 1698431365
transform -1 0 15568 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _353_
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _354_
timestamp 1698431365
transform 1 0 13216 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _355_
timestamp 1698431365
transform 1 0 12432 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _356_
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _357_
timestamp 1698431365
transform 1 0 13216 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _358_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _359_
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _360_
timestamp 1698431365
transform -1 0 13216 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _361_
timestamp 1698431365
transform -1 0 11200 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1698431365
transform -1 0 4144 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _391_
timestamp 1698431365
transform -1 0 6160 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1698431365
transform 1 0 10192 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _393_
timestamp 1698431365
transform -1 0 7392 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1698431365
transform -1 0 4480 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _395_
timestamp 1698431365
transform 1 0 7840 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1698431365
transform -1 0 6160 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1698431365
transform -1 0 6832 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1698431365
transform -1 0 3472 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _400_
timestamp 1698431365
transform 1 0 6832 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1698431365
transform 1 0 2128 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _402_
timestamp 1698431365
transform -1 0 6832 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _403_
timestamp 1698431365
transform -1 0 6720 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1698431365
transform -1 0 5376 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _406_
timestamp 1698431365
transform -1 0 3472 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1698431365
transform -1 0 10864 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _408_
timestamp 1698431365
transform -1 0 3472 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1698431365
transform -1 0 3584 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1698431365
transform -1 0 3808 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1698431365
transform -1 0 4816 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _412_
timestamp 1698431365
transform -1 0 4928 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1698431365
transform -1 0 6048 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _414_
timestamp 1698431365
transform 1 0 7504 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1698431365
transform -1 0 5152 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _416_
timestamp 1698431365
transform 1 0 6832 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _417_
timestamp 1698431365
transform -1 0 3808 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _418_
timestamp 1698431365
transform 1 0 9520 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _419_
timestamp 1698431365
transform -1 0 3808 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _420_
timestamp 1698431365
transform 1 0 8176 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _421_
timestamp 1698431365
transform -1 0 4256 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__I
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1698431365
transform 1 0 28000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__I
timestamp 1698431365
transform -1 0 29568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__I
timestamp 1698431365
transform -1 0 27664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__I
timestamp 1698431365
transform 1 0 32032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__I
timestamp 1698431365
transform 1 0 32368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__I
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__I
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__I
timestamp 1698431365
transform 1 0 33488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I
timestamp 1698431365
transform -1 0 38528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1698431365
transform 1 0 40992 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1698431365
transform 1 0 39872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1698431365
transform 1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1698431365
transform -1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1698431365
transform 1 0 21728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1698431365
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1698431365
transform 1 0 30240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__I
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1698431365
transform 1 0 40992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I
timestamp 1698431365
transform -1 0 40096 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1698431365
transform -1 0 37856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1698431365
transform 1 0 35728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I
timestamp 1698431365
transform -1 0 26208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1698431365
transform -1 0 37296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1698431365
transform 1 0 36064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__I
timestamp 1698431365
transform -1 0 32816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I
timestamp 1698431365
transform 1 0 40992 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__I
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I
timestamp 1698431365
transform 1 0 31360 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__I
timestamp 1698431365
transform 1 0 31920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__I
timestamp 1698431365
transform 1 0 29680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I
timestamp 1698431365
transform -1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__I
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698431365
transform -1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698431365
transform -1 0 9856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698431365
transform 1 0 14560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698431365
transform 1 0 13888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__CLK
timestamp 1698431365
transform -1 0 12208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__CLK
timestamp 1698431365
transform 1 0 11200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__CLK
timestamp 1698431365
transform 1 0 10416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__CLK
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__CLK
timestamp 1698431365
transform -1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__CLK
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__CLK
timestamp 1698431365
transform -1 0 19488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__CLK
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__CLK
timestamp 1698431365
transform 1 0 16128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__CLK
timestamp 1698431365
transform 1 0 18928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__277__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__CLK
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__CLK
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__CLK
timestamp 1698431365
transform -1 0 34496 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__CLK
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__CLK
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__CLK
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__CLK
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__CLK
timestamp 1698431365
transform 1 0 36960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__CLK
timestamp 1698431365
transform 1 0 35952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__CLK
timestamp 1698431365
transform 1 0 37632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__CLK
timestamp 1698431365
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__CLK
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__CLK
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__CLK
timestamp 1698431365
transform -1 0 34944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__CLK
timestamp 1698431365
transform 1 0 26432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__CLK
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__CLK
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__CLK
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__CLK
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__CLK
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__CLK
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__CLK
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__CLK
timestamp 1698431365
transform 1 0 39760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__CLK
timestamp 1698431365
transform 1 0 36064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__CLK
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__CLK
timestamp 1698431365
transform 1 0 37184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__CLK
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__CLK
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__CLK
timestamp 1698431365
transform -1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__CLK
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__CLK
timestamp 1698431365
transform 1 0 36960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__CLK
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__CLK
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__CLK
timestamp 1698431365
transform 1 0 33376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__CLK
timestamp 1698431365
transform -1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__CLK
timestamp 1698431365
transform 1 0 32368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__CLK
timestamp 1698431365
transform 1 0 30128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__CLK
timestamp 1698431365
transform 1 0 27328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__CLK
timestamp 1698431365
transform 1 0 26096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__CLK
timestamp 1698431365
transform 1 0 21392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__CLK
timestamp 1698431365
transform -1 0 19488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__CLK
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__CLK
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__CLK
timestamp 1698431365
transform 1 0 12208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__CLK
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__CLK
timestamp 1698431365
transform -1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__CLK
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__CLK
timestamp 1698431365
transform -1 0 11312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__CLK
timestamp 1698431365
transform -1 0 8512 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__CLK
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__CLK
timestamp 1698431365
transform 1 0 17360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__CLK
timestamp 1698431365
transform 1 0 15680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__CLK
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__CLK
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__CLK
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__CLK
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__I
timestamp 1698431365
transform -1 0 9072 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__I
timestamp 1698431365
transform -1 0 10304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_prog_clk_I
timestamp 1698431365
transform 1 0 15904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_prog_clk_I
timestamp 1698431365
transform -1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_prog_clk_I
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_prog_clk_I
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_prog_clk_I
timestamp 1698431365
transform 1 0 25760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_prog_clk_I
timestamp 1698431365
transform 1 0 33488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_prog_clk_I
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_prog_clk_I
timestamp 1698431365
transform -1 0 33264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 21616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 4928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 1792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 10192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 19936 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 4368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 9632 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 1792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 3136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 1792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 7056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 7504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 22960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 4368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 5712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 4816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 26320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 10192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 5264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 25648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 2016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 5712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 6160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 18928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 3808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 3584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1698431365
transform 1 0 26768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output62_I
timestamp 1698431365
transform 1 0 25760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1698431365
transform -1 0 15680 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1698431365
transform 1 0 14560 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1698431365
transform -1 0 15680 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1698431365
transform 1 0 14672 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1698431365
transform -1 0 32368 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1698431365
transform 1 0 26768 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_30
timestamp 1698431365
transform 1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_40 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_53
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_64
timestamp 1698431365
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_76
timestamp 1698431365
transform 1 0 9856 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_95
timestamp 1698431365
transform 1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_108 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_124 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_132
timestamp 1698431365
transform 1 0 16128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_358
timestamp 1698431365
transform 1 0 41440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_12
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_25
timestamp 1698431365
transform 1 0 4144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_29
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_33
timestamp 1698431365
transform 1 0 5040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_37
timestamp 1698431365
transform 1 0 5488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_41
timestamp 1698431365
transform 1 0 5936 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_57
timestamp 1698431365
transform 1 0 7728 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_65
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_360
timestamp 1698431365
transform 1 0 41664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_364
timestamp 1698431365
transform 1 0 42112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_6
timestamp 1698431365
transform 1 0 2016 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_31
timestamp 1698431365
transform 1 0 4816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_45
timestamp 1698431365
transform 1 0 6384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_55
timestamp 1698431365
transform 1 0 7504 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_71
timestamp 1698431365
transform 1 0 9296 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_85
timestamp 1698431365
transform 1 0 10864 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_349
timestamp 1698431365
transform 1 0 40432 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_365
timestamp 1698431365
transform 1 0 42224 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_22
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_54
timestamp 1698431365
transform 1 0 7392 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_360
timestamp 1698431365
transform 1 0 41664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_364
timestamp 1698431365
transform 1 0 42112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_16
timestamp 1698431365
transform 1 0 3136 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_349
timestamp 1698431365
transform 1 0 40432 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_365
timestamp 1698431365
transform 1 0 42224 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_16
timestamp 1698431365
transform 1 0 3136 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_48
timestamp 1698431365
transform 1 0 6720 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_104
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_121
timestamp 1698431365
transform 1 0 14896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_137
timestamp 1698431365
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_360
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_364
timestamp 1698431365
transform 1 0 42112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_20
timestamp 1698431365
transform 1 0 3584 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_57
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_93
timestamp 1698431365
transform 1 0 11760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_97
timestamp 1698431365
transform 1 0 12208 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_123
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_164
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_349
timestamp 1698431365
transform 1 0 40432 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_365
timestamp 1698431365
transform 1 0 42224 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_16
timestamp 1698431365
transform 1 0 3136 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_48
timestamp 1698431365
transform 1 0 6720 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_83
timestamp 1698431365
transform 1 0 10640 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_91
timestamp 1698431365
transform 1 0 11536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_93
timestamp 1698431365
transform 1 0 11760 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_110
timestamp 1698431365
transform 1 0 13664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_114
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_122
timestamp 1698431365
transform 1 0 15008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_152
timestamp 1698431365
transform 1 0 18368 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_168
timestamp 1698431365
transform 1 0 20160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_172
timestamp 1698431365
transform 1 0 20608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_360
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_364
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_16
timestamp 1698431365
transform 1 0 3136 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_154
timestamp 1698431365
transform 1 0 18592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_162
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_209
timestamp 1698431365
transform 1 0 24752 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_225
timestamp 1698431365
transform 1 0 26544 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_249
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_262
timestamp 1698431365
transform 1 0 30688 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_333
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_351
timestamp 1698431365
transform 1 0 40656 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_359
timestamp 1698431365
transform 1 0 41552 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_363
timestamp 1698431365
transform 1 0 42000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_365
timestamp 1698431365
transform 1 0 42224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_97
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_152
timestamp 1698431365
transform 1 0 18368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_198
timestamp 1698431365
transform 1 0 23520 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_240
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_248
timestamp 1698431365
transform 1 0 29120 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_252
timestamp 1698431365
transform 1 0 29568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_270
timestamp 1698431365
transform 1 0 31584 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_296
timestamp 1698431365
transform 1 0 34496 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_312
timestamp 1698431365
transform 1 0 36288 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_332
timestamp 1698431365
transform 1 0 38528 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_348
timestamp 1698431365
transform 1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_364
timestamp 1698431365
transform 1 0 42112 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_117
timestamp 1698431365
transform 1 0 14448 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_202
timestamp 1698431365
transform 1 0 23968 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_210
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_214
timestamp 1698431365
transform 1 0 25312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_306
timestamp 1698431365
transform 1 0 35616 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_312
timestamp 1698431365
transform 1 0 36288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_327
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_332
timestamp 1698431365
transform 1 0 38528 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_348
timestamp 1698431365
transform 1 0 40320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_82
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_129
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_326
timestamp 1698431365
transform 1 0 37856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_342
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_364
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_86
timestamp 1698431365
transform 1 0 10976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_90
timestamp 1698431365
transform 1 0 11424 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_118
timestamp 1698431365
transform 1 0 14560 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_126
timestamp 1698431365
transform 1 0 15456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_130
timestamp 1698431365
transform 1 0 15904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_158
timestamp 1698431365
transform 1 0 19040 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_281
timestamp 1698431365
transform 1 0 32816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_285
timestamp 1698431365
transform 1 0 33264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_289
timestamp 1698431365
transform 1 0 33712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_306
timestamp 1698431365
transform 1 0 35616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_355
timestamp 1698431365
transform 1 0 41104 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_363
timestamp 1698431365
transform 1 0 42000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_365
timestamp 1698431365
transform 1 0 42224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_48
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_52
timestamp 1698431365
transform 1 0 7168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_97
timestamp 1698431365
transform 1 0 12208 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_105
timestamp 1698431365
transform 1 0 13104 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_255
timestamp 1698431365
transform 1 0 29904 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_263
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_316
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_320
timestamp 1698431365
transform 1 0 37184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_322
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_339
timestamp 1698431365
transform 1 0 39312 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_345
timestamp 1698431365
transform 1 0 39984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_360
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_364
timestamp 1698431365
transform 1 0 42112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_79
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_87
timestamp 1698431365
transform 1 0 11088 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_195
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_203
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_221
timestamp 1698431365
transform 1 0 26096 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_229
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_253
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_270
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_274
timestamp 1698431365
transform 1 0 32032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_276
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_289
timestamp 1698431365
transform 1 0 33712 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_351
timestamp 1698431365
transform 1 0 40656 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_359
timestamp 1698431365
transform 1 0 41552 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_363
timestamp 1698431365
transform 1 0 42000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_365
timestamp 1698431365
transform 1 0 42224 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_19
timestamp 1698431365
transform 1 0 3472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_27
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_62
timestamp 1698431365
transform 1 0 8288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_125
timestamp 1698431365
transform 1 0 15344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_167
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698431365
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_228
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_232
timestamp 1698431365
transform 1 0 27328 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_249
timestamp 1698431365
transform 1 0 29232 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_253
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_257
timestamp 1698431365
transform 1 0 30128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_307
timestamp 1698431365
transform 1 0 35728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_311
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_313
timestamp 1698431365
transform 1 0 36400 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_360
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_364
timestamp 1698431365
transform 1 0 42112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_75
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_79
timestamp 1698431365
transform 1 0 10192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_96
timestamp 1698431365
transform 1 0 12096 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_117
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698431365
transform 1 0 23184 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_230
timestamp 1698431365
transform 1 0 27104 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_353
timestamp 1698431365
transform 1 0 40880 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_361
timestamp 1698431365
transform 1 0 41776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_365
timestamp 1698431365
transform 1 0 42224 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_36
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_40
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_52
timestamp 1698431365
transform 1 0 7168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_128
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_132
timestamp 1698431365
transform 1 0 16128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698431365
transform 1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_156
timestamp 1698431365
transform 1 0 18816 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1698431365
transform 1 0 22960 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_254
timestamp 1698431365
transform 1 0 29792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_271
timestamp 1698431365
transform 1 0 31696 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_318
timestamp 1698431365
transform 1 0 36960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_322
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_326
timestamp 1698431365
transform 1 0 37856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_330
timestamp 1698431365
transform 1 0 38304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_347
timestamp 1698431365
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_364
timestamp 1698431365
transform 1 0 42112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_4
timestamp 1698431365
transform 1 0 1792 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_41
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_43
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_62
timestamp 1698431365
transform 1 0 8288 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_70
timestamp 1698431365
transform 1 0 9184 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_121
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_129
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_189
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_232
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_285
timestamp 1698431365
transform 1 0 33264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_289
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_309
timestamp 1698431365
transform 1 0 35952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_352
timestamp 1698431365
transform 1 0 40768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_356
timestamp 1698431365
transform 1 0 41216 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_364
timestamp 1698431365
transform 1 0 42112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_4
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_49
timestamp 1698431365
transform 1 0 6832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_74
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_91
timestamp 1698431365
transform 1 0 11536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_99
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_134
timestamp 1698431365
transform 1 0 16352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_176
timestamp 1698431365
transform 1 0 21056 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_192
timestamp 1698431365
transform 1 0 22848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_225
timestamp 1698431365
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_342
timestamp 1698431365
transform 1 0 39648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_364
timestamp 1698431365
transform 1 0 42112 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_57
timestamp 1698431365
transform 1 0 7728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_100
timestamp 1698431365
transform 1 0 12544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_211
timestamp 1698431365
transform 1 0 24976 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_215
timestamp 1698431365
transform 1 0 25424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_217
timestamp 1698431365
transform 1 0 25648 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_236
timestamp 1698431365
transform 1 0 27776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_281
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_285
timestamp 1698431365
transform 1 0 33264 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_289
timestamp 1698431365
transform 1 0 33712 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_306
timestamp 1698431365
transform 1 0 35616 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_342
timestamp 1698431365
transform 1 0 39648 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_358
timestamp 1698431365
transform 1 0 41440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_10
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_76
timestamp 1698431365
transform 1 0 9856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_122
timestamp 1698431365
transform 1 0 15008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_126
timestamp 1698431365
transform 1 0 15456 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_180
timestamp 1698431365
transform 1 0 21504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_184
timestamp 1698431365
transform 1 0 21952 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_200
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_222
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_272
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_292
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_300
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_335
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_339
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_360
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_364
timestamp 1698431365
transform 1 0 42112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_88
timestamp 1698431365
transform 1 0 11200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_92
timestamp 1698431365
transform 1 0 11648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_102
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_141
timestamp 1698431365
transform 1 0 17136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_145
timestamp 1698431365
transform 1 0 17584 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_162
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_166
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_170
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698431365
transform 1 0 28000 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_259
timestamp 1698431365
transform 1 0 30352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_261
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_296
timestamp 1698431365
transform 1 0 34496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_300
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_304
timestamp 1698431365
transform 1 0 35392 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_319
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_322
timestamp 1698431365
transform 1 0 37408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_342
timestamp 1698431365
transform 1 0 39648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_346
timestamp 1698431365
transform 1 0 40096 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_362
timestamp 1698431365
transform 1 0 41888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_44
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_61
timestamp 1698431365
transform 1 0 8176 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_170
timestamp 1698431365
transform 1 0 20384 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_292
timestamp 1698431365
transform 1 0 34048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_294
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_364
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_8
timestamp 1698431365
transform 1 0 2240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_12
timestamp 1698431365
transform 1 0 2688 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_62
timestamp 1698431365
transform 1 0 8288 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_162
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_164
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_352
timestamp 1698431365
transform 1 0 40768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_356
timestamp 1698431365
transform 1 0 41216 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_364
timestamp 1698431365
transform 1 0 42112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_36
timestamp 1698431365
transform 1 0 5376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_40
timestamp 1698431365
transform 1 0 5824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_61
timestamp 1698431365
transform 1 0 8176 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_90
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_92
timestamp 1698431365
transform 1 0 11648 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_127
timestamp 1698431365
transform 1 0 15568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_135
timestamp 1698431365
transform 1 0 16464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_180
timestamp 1698431365
transform 1 0 21504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_184
timestamp 1698431365
transform 1 0 21952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_201
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698431365
transform 1 0 31360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_307
timestamp 1698431365
transform 1 0 35728 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_309
timestamp 1698431365
transform 1 0 35952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_344
timestamp 1698431365
transform 1 0 39872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_364
timestamp 1698431365
transform 1 0 42112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_88
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_96
timestamp 1698431365
transform 1 0 12096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_109
timestamp 1698431365
transform 1 0 13552 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_126
timestamp 1698431365
transform 1 0 15456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_130
timestamp 1698431365
transform 1 0 15904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_134
timestamp 1698431365
transform 1 0 16352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_202
timestamp 1698431365
transform 1 0 23968 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_210
timestamp 1698431365
transform 1 0 24864 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_227
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_257
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_260
timestamp 1698431365
transform 1 0 30464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_305
timestamp 1698431365
transform 1 0 35504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_352
timestamp 1698431365
transform 1 0 40768 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_360
timestamp 1698431365
transform 1 0 41664 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_364
timestamp 1698431365
transform 1 0 42112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_16
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_40
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_58
timestamp 1698431365
transform 1 0 7840 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_134
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_154
timestamp 1698431365
transform 1 0 18592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_195
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_222
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_238
timestamp 1698431365
transform 1 0 28000 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_242
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_307
timestamp 1698431365
transform 1 0 35728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_309
timestamp 1698431365
transform 1 0 35952 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_312
timestamp 1698431365
transform 1 0 36288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_342
timestamp 1698431365
transform 1 0 39648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_364
timestamp 1698431365
transform 1 0 42112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_16
timestamp 1698431365
transform 1 0 3136 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_71
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_75
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_83
timestamp 1698431365
transform 1 0 10640 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_169
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_225
timestamp 1698431365
transform 1 0 26544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_229
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698431365
transform 1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_353
timestamp 1698431365
transform 1 0 40880 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_361
timestamp 1698431365
transform 1 0 41776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_365
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_22
timestamp 1698431365
transform 1 0 3808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_30
timestamp 1698431365
transform 1 0 4704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_34
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_96
timestamp 1698431365
transform 1 0 12096 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_173
timestamp 1698431365
transform 1 0 20720 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698431365
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_342
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_364
timestamp 1698431365
transform 1 0 42112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_16
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_47
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_161
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_187
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_203
timestamp 1698431365
transform 1 0 24080 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_281
timestamp 1698431365
transform 1 0 32816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_285
timestamp 1698431365
transform 1 0 33264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_289
timestamp 1698431365
transform 1 0 33712 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_297
timestamp 1698431365
transform 1 0 34608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_352
timestamp 1698431365
transform 1 0 40768 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_360
timestamp 1698431365
transform 1 0 41664 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_364
timestamp 1698431365
transform 1 0 42112 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_8
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_28
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_90
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_94
timestamp 1698431365
transform 1 0 11872 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_96
timestamp 1698431365
transform 1 0 12096 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_181
timestamp 1698431365
transform 1 0 21616 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_197
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698431365
transform 1 0 24304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_218
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_260
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_341
timestamp 1698431365
transform 1 0 39536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_345
timestamp 1698431365
transform 1 0 39984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_360
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_364
timestamp 1698431365
transform 1 0 42112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_113
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_202
timestamp 1698431365
transform 1 0 23968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_251
timestamp 1698431365
transform 1 0 29456 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_275
timestamp 1698431365
transform 1 0 32144 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_310
timestamp 1698431365
transform 1 0 36064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_351
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_359
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_363
timestamp 1698431365
transform 1 0 42000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_365
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_117
timestamp 1698431365
transform 1 0 14448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_119
timestamp 1698431365
transform 1 0 14672 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_169
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_237
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_241
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_245
timestamp 1698431365
transform 1 0 28784 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_262
timestamp 1698431365
transform 1 0 30688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_266
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_288
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_308
timestamp 1698431365
transform 1 0 35840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_312
timestamp 1698431365
transform 1 0 36288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_356
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_364
timestamp 1698431365
transform 1 0 42112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_14
timestamp 1698431365
transform 1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_18
timestamp 1698431365
transform 1 0 3360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_22
timestamp 1698431365
transform 1 0 3808 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_30
timestamp 1698431365
transform 1 0 4704 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_95
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_219
timestamp 1698431365
transform 1 0 25872 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_223
timestamp 1698431365
transform 1 0 26320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_227
timestamp 1698431365
transform 1 0 26768 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_257
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_292
timestamp 1698431365
transform 1 0 34048 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_362
timestamp 1698431365
transform 1 0 41888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_16
timestamp 1698431365
transform 1 0 3136 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_89
timestamp 1698431365
transform 1 0 11312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_125
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_129
timestamp 1698431365
transform 1 0 15792 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_216
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_251
timestamp 1698431365
transform 1 0 29456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_255
timestamp 1698431365
transform 1 0 29904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_259
timestamp 1698431365
transform 1 0 30352 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_316
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_320
timestamp 1698431365
transform 1 0 37184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_324
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_341
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_364
timestamp 1698431365
transform 1 0 42112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_16
timestamp 1698431365
transform 1 0 3136 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_80
timestamp 1698431365
transform 1 0 10304 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_84
timestamp 1698431365
transform 1 0 10752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_86
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_119
timestamp 1698431365
transform 1 0 14672 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_125
timestamp 1698431365
transform 1 0 15344 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_181
timestamp 1698431365
transform 1 0 21616 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_189
timestamp 1698431365
transform 1 0 22512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_195
timestamp 1698431365
transform 1 0 23184 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_230
timestamp 1698431365
transform 1 0 27104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_234
timestamp 1698431365
transform 1 0 27552 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_327
timestamp 1698431365
transform 1 0 37968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_331
timestamp 1698431365
transform 1 0 38416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_333
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_350
timestamp 1698431365
transform 1 0 40544 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_22
timestamp 1698431365
transform 1 0 3808 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_30
timestamp 1698431365
transform 1 0 4704 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_36
timestamp 1698431365
transform 1 0 5376 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_53
timestamp 1698431365
transform 1 0 7280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_89
timestamp 1698431365
transform 1 0 11312 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_105
timestamp 1698431365
transform 1 0 13104 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_113
timestamp 1698431365
transform 1 0 14000 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_117
timestamp 1698431365
transform 1 0 14448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_119
timestamp 1698431365
transform 1 0 14672 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_162
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_164
timestamp 1698431365
transform 1 0 19712 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_181
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_197
timestamp 1698431365
transform 1 0 23408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_201
timestamp 1698431365
transform 1 0 23856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_203
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_218
timestamp 1698431365
transform 1 0 25760 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_225
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_275
timestamp 1698431365
transform 1 0 32144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_292
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_329
timestamp 1698431365
transform 1 0 38192 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_331
timestamp 1698431365
transform 1 0 38416 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_342
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_360
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_364
timestamp 1698431365
transform 1 0 42112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_53
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_61
timestamp 1698431365
transform 1 0 8176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_81
timestamp 1698431365
transform 1 0 10416 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_97
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_119
timestamp 1698431365
transform 1 0 14672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_121
timestamp 1698431365
transform 1 0 14896 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_154
timestamp 1698431365
transform 1 0 18592 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_170
timestamp 1698431365
transform 1 0 20384 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_193
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_201
timestamp 1698431365
transform 1 0 23856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_203
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_220
timestamp 1698431365
transform 1 0 25984 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_228
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_272
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_276
timestamp 1698431365
transform 1 0 32256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_278
timestamp 1698431365
transform 1 0 32480 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_297
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_346
timestamp 1698431365
transform 1 0 40096 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_362
timestamp 1698431365
transform 1 0 41888 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_10
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_42
timestamp 1698431365
transform 1 0 6048 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_104
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_170
timestamp 1698431365
transform 1 0 20384 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_202
timestamp 1698431365
transform 1 0 23968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_237
timestamp 1698431365
transform 1 0 27888 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_310
timestamp 1698431365
transform 1 0 36064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_318
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_335
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_343
timestamp 1698431365
transform 1 0 39760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_347
timestamp 1698431365
transform 1 0 40208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_364
timestamp 1698431365
transform 1 0 42112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_20
timestamp 1698431365
transform 1 0 3584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_24
timestamp 1698431365
transform 1 0 4032 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_351
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_359
timestamp 1698431365
transform 1 0 41552 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_363
timestamp 1698431365
transform 1 0 42000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_365
timestamp 1698431365
transform 1 0 42224 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_12
timestamp 1698431365
transform 1 0 2688 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_25
timestamp 1698431365
transform 1 0 4144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_29
timestamp 1698431365
transform 1 0 4592 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_61
timestamp 1698431365
transform 1 0 8176 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_41
timestamp 1698431365
transform 1 0 5936 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_349
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_40
timestamp 1698431365
transform 1 0 5824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_42
timestamp 1698431365
transform 1 0 6048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_47
timestamp 1698431365
transform 1 0 6608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_51
timestamp 1698431365
transform 1 0 7056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_55
timestamp 1698431365
transform 1 0 7504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_65
timestamp 1698431365
transform 1 0 8624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_364
timestamp 1698431365
transform 1 0 42112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_85
timestamp 1698431365
transform 1 0 10864 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_365
timestamp 1698431365
transform 1 0 42224 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_16
timestamp 1698431365
transform 1 0 3136 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_112
timestamp 1698431365
transform 1 0 13888 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_128
timestamp 1698431365
transform 1 0 15680 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_223
timestamp 1698431365
transform 1 0 26320 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_229
timestamp 1698431365
transform 1 0 26992 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_261
timestamp 1698431365
transform 1 0 30576 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_277
timestamp 1698431365
transform 1 0 32368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_360
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_364
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_6
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_8
timestamp 1698431365
transform 1 0 2240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_19
timestamp 1698431365
transform 1 0 3472 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_33
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_77
timestamp 1698431365
transform 1 0 9968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_89
timestamp 1698431365
transform 1 0 11312 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_131
timestamp 1698431365
transform 1 0 16016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_143
timestamp 1698431365
transform 1 0 17360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_147
timestamp 1698431365
transform 1 0 17808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_163
timestamp 1698431365
transform 1 0 19600 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_167
timestamp 1698431365
transform 1 0 20048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_173
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_181
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_189
timestamp 1698431365
transform 1 0 22512 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_197
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_205
timestamp 1698431365
transform 1 0 24304 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_213
timestamp 1698431365
transform 1 0 25200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_239
timestamp 1698431365
transform 1 0 28112 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_243
timestamp 1698431365
transform 1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_349
timestamp 1698431365
transform 1 0 40432 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_365
timestamp 1698431365
transform 1 0 42224 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_36
timestamp 1698431365
transform 1 0 5376 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_51
timestamp 1698431365
transform 1 0 7056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_53
timestamp 1698431365
transform 1 0 7280 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_78
timestamp 1698431365
transform 1 0 10080 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_101
timestamp 1698431365
transform 1 0 12656 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_108
timestamp 1698431365
transform 1 0 13440 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_113
timestamp 1698431365
transform 1 0 14000 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_149
timestamp 1698431365
transform 1 0 18032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_161
timestamp 1698431365
transform 1 0 19376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_163
timestamp 1698431365
transform 1 0 19600 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_178
timestamp 1698431365
transform 1 0 21280 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_180
timestamp 1698431365
transform 1 0 21504 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_201
timestamp 1698431365
transform 1 0 23856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_203
timestamp 1698431365
transform 1 0 24080 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_230
timestamp 1698431365
transform 1 0 27104 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_240
timestamp 1698431365
transform 1 0 28224 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_274
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_308
timestamp 1698431365
transform 1 0 35840 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_342
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_358
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 35616 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 30688 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 40208 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 31584 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform -1 0 39648 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 34944 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 23968 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 14896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 23968 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 20384 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform 1 0 19264 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 27328 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 35728 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform 1 0 9744 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 26096 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 16800 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 16576 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform 1 0 10304 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform 1 0 6384 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform -1 0 39648 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform -1 0 39648 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform -1 0 42336 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 36064 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 39648 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform 1 0 7504 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform -1 0 39984 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 42336 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 35616 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 17920 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform -1 0 18144 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform 1 0 37072 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform 1 0 9520 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform -1 0 34608 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 27888 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 32704 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform -1 0 22624 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform -1 0 12992 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold50
timestamp 1698431365
transform -1 0 9296 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform -1 0 39536 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform -1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform -1 0 32144 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform -1 0 8512 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 40096 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform -1 0 39536 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform -1 0 7840 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform -1 0 20384 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform -1 0 29232 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 27888 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform 1 0 13664 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform 1 0 29792 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 35616 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform 1 0 5488 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform -1 0 10304 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold69
timestamp 1698431365
transform -1 0 20048 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold70
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold71
timestamp 1698431365
transform 1 0 6496 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold72
timestamp 1698431365
transform -1 0 28672 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold73
timestamp 1698431365
transform -1 0 36624 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold74
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold75
timestamp 1698431365
transform 1 0 38752 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold76
timestamp 1698431365
transform 1 0 17920 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold77
timestamp 1698431365
transform -1 0 35728 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold78
timestamp 1698431365
transform 1 0 38864 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold79
timestamp 1698431365
transform 1 0 17696 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold80
timestamp 1698431365
transform -1 0 13104 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold81
timestamp 1698431365
transform -1 0 38528 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold82
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold83
timestamp 1698431365
transform -1 0 35728 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold84
timestamp 1698431365
transform -1 0 13664 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold85
timestamp 1698431365
transform -1 0 27776 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold86
timestamp 1698431365
transform -1 0 16576 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold87
timestamp 1698431365
transform -1 0 38528 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold88
timestamp 1698431365
transform -1 0 31808 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold89
timestamp 1698431365
transform -1 0 23968 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold90
timestamp 1698431365
transform -1 0 10416 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold91
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold92
timestamp 1698431365
transform 1 0 6384 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold93
timestamp 1698431365
transform -1 0 20048 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold94
timestamp 1698431365
transform -1 0 31696 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold95
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold96
timestamp 1698431365
transform -1 0 12208 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold97
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold98
timestamp 1698431365
transform 1 0 37520 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold99
timestamp 1698431365
transform 1 0 38864 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold100
timestamp 1698431365
transform -1 0 16688 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold101
timestamp 1698431365
transform -1 0 39648 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold102
timestamp 1698431365
transform -1 0 24864 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold103
timestamp 1698431365
transform -1 0 20048 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold104
timestamp 1698431365
transform -1 0 20384 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold105
timestamp 1698431365
transform 1 0 1680 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold106
timestamp 1698431365
transform -1 0 30464 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold107
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold108
timestamp 1698431365
transform -1 0 32368 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold109
timestamp 1698431365
transform -1 0 32256 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold110
timestamp 1698431365
transform -1 0 20048 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold111
timestamp 1698431365
transform -1 0 25984 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 22288 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 9856 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 17584 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 21280 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 4144 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 8176 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 6832 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 8176 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 24304 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 4256 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 5824 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 26992 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 10192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 26320 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 6160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 19600 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 4256 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 3472 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3136 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output39
timestamp 1698431365
transform -1 0 3136 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output40
timestamp 1698431365
transform -1 0 3472 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41
timestamp 1698431365
transform 1 0 10864 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output42 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3584 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output43
timestamp 1698431365
transform -1 0 3136 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 8848 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output45
timestamp 1698431365
transform -1 0 5152 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output46
timestamp 1698431365
transform -1 0 7056 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output47
timestamp 1698431365
transform -1 0 3136 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output49
timestamp 1698431365
transform 1 0 15008 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output50
timestamp 1698431365
transform -1 0 3136 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output51
timestamp 1698431365
transform -1 0 3136 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output52
timestamp 1698431365
transform -1 0 3136 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output53
timestamp 1698431365
transform -1 0 3136 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform -1 0 3136 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output55
timestamp 1698431365
transform -1 0 3136 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output56
timestamp 1698431365
transform 1 0 10192 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output57
timestamp 1698431365
transform -1 0 3136 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output58
timestamp 1698431365
transform -1 0 8960 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform -1 0 3136 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output60
timestamp 1698431365
transform 1 0 16240 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output61
timestamp 1698431365
transform -1 0 3136 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output62
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output63
timestamp 1698431365
transform -1 0 4704 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output64
timestamp 1698431365
transform 1 0 22288 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform -1 0 5040 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform -1 0 3136 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform -1 0 3136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 18256 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output69
timestamp 1698431365
transform -1 0 3136 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_48 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 42560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_49
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_50
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 42560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 42560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 42560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 42560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 42560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 42560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 42560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 42560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 42560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 42560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 42560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 42560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 42560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 42560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 42560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 42560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 42560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 42560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 42560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 42560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 42560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 42560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 42560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 42560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 42560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 42560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 42560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 42560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 42560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 42560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 42560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 42560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 42560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 42560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 42560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__71
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__72
timestamp 1698431365
transform -1 0 3584 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__73
timestamp 1698431365
transform -1 0 13440 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__74
timestamp 1698431365
transform -1 0 2688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__75
timestamp 1698431365
transform 1 0 14560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__76
timestamp 1698431365
transform -1 0 2464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__77
timestamp 1698431365
transform -1 0 13440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__78
timestamp 1698431365
transform -1 0 23408 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__79
timestamp 1698431365
transform -1 0 18032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__80
timestamp 1698431365
transform -1 0 11312 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__81
timestamp 1698431365
transform -1 0 12208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__82
timestamp 1698431365
transform -1 0 9632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__83
timestamp 1698431365
transform -1 0 12656 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__84
timestamp 1698431365
transform -1 0 14560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__85
timestamp 1698431365
transform -1 0 6608 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__86
timestamp 1698431365
transform -1 0 2688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__87
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__88
timestamp 1698431365
transform -1 0 4256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__89
timestamp 1698431365
transform -1 0 20720 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__90
timestamp 1698431365
transform -1 0 3584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__91
timestamp 1698431365
transform -1 0 14000 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__92
timestamp 1698431365
transform -1 0 10864 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__93
timestamp 1698431365
transform -1 0 2016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__94
timestamp 1698431365
transform -1 0 2016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__95
timestamp 1698431365
transform 1 0 19936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_1__0__96
timestamp 1698431365
transform -1 0 7840 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_106
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_107
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_108
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_109
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_110
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_111
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_112
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_113
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_114
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_115
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_116
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_117
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_118
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_119
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_120
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_121
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_122
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_123
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_124
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_125
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_126
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_127
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_128
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_129
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_130
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_131
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_132
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_133
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_134
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_135
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_136
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_137
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_138
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_139
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_140
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_141
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_142
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_143
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_144
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_145
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_146
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_147
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_148
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_149
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_150
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_151
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_152
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_153
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_154
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_155
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_156
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_157
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_158
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_159
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_160
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_161
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_162
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_163
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_164
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_165
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_166
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_167
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_168
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_169
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_170
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_171
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_172
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_173
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_174
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_175
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_176
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_177
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_178
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_179
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_180
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_181
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_182
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_183
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_184
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_185
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_186
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_187
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_188
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_189
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_190
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_191
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_192
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_193
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_194
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_195
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_196
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_197
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_198
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_199
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_200
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_201
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_202
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_203
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_204
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_205
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_206
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_207
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_208
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_211
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_212
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_215
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_216
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_217
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_218
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_219
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_220
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_221
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_222
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_223
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_224
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_225
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_226
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_227
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_228
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_229
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_230
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_231
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_232
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_233
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_234
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_235
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_236
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_237
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_238
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_239
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_240
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_241
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_242
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_243
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_244
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_245
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_246
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_247
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_248
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_249
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_250
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_251
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_252
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_253
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_254
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_255
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_256
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_257
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_258
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_259
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_260
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_261
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_262
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_263
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_264
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_265
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_266
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_267
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_268
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_269
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_270
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_271
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_272
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_273
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_274
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_275
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_276
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_277
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_278
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_279
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_280
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_281
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_282
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_283
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_284
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_285
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_286
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_287
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_288
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_289
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_290
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_291
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_292
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_293
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_294
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_295
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_296
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_297
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_298
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_299
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_300
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_301
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_302
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_303
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_304
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_305
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_306
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_307
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_308
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_309
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_310
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_311
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_312
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_313
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_314
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_315
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_316
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_317
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_318
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_319
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_320
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_321
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_322
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_323
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_324
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_325
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_326
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_327
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_328
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_329
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_330
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_331
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_332
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_333
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_334
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_335
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_336
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_337
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_338
timestamp 1698431365
transform 1 0 12768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_339
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_340
timestamp 1698431365
transform 1 0 20384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 28000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_343
timestamp 1698431365
transform 1 0 31808 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_344
timestamp 1698431365
transform 1 0 35616 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_345
timestamp 1698431365
transform 1 0 39424 0 -1 40768
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 ccff_head
port 0 nsew signal input
flabel metal2 s 26880 43200 26992 44000 0 FreeSans 448 90 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 21504 43200 21616 44000 0 FreeSans 448 90 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal3 s 0 0 800 112 0 FreeSans 448 0 0 0 chanx_left_in[10]
port 3 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 chanx_left_in[11]
port 4 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 chanx_left_in[12]
port 5 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 chanx_left_in[13]
port 6 nsew signal input
flabel metal2 s 16800 43200 16912 44000 0 FreeSans 448 90 0 0 chanx_left_in[14]
port 7 nsew signal input
flabel metal2 s 19488 43200 19600 44000 0 FreeSans 448 90 0 0 chanx_left_in[15]
port 8 nsew signal input
flabel metal3 s 0 2016 800 2128 0 FreeSans 448 0 0 0 chanx_left_in[16]
port 9 nsew signal input
flabel metal2 s 0 43200 112 44000 0 FreeSans 448 90 0 0 chanx_left_in[17]
port 10 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 chanx_left_in[18]
port 11 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 chanx_left_in[19]
port 12 nsew signal input
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 chanx_left_in[1]
port 13 nsew signal input
flabel metal2 s 6720 43200 6832 44000 0 FreeSans 448 90 0 0 chanx_left_in[2]
port 14 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 chanx_left_in[3]
port 15 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 chanx_left_in[4]
port 16 nsew signal input
flabel metal2 s 23520 43200 23632 44000 0 FreeSans 448 90 0 0 chanx_left_in[5]
port 17 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 chanx_left_in[6]
port 18 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 chanx_left_in[7]
port 19 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 chanx_left_in[8]
port 20 nsew signal input
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 chanx_left_in[9]
port 21 nsew signal input
flabel metal2 s 7392 43200 7504 44000 0 FreeSans 448 90 0 0 chanx_left_out[0]
port 22 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 chanx_left_out[10]
port 23 nsew signal tristate
flabel metal2 s 24192 43200 24304 44000 0 FreeSans 448 90 0 0 chanx_left_out[11]
port 24 nsew signal tristate
flabel metal3 s 0 1344 800 1456 0 FreeSans 448 0 0 0 chanx_left_out[12]
port 25 nsew signal tristate
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 chanx_left_out[13]
port 26 nsew signal tristate
flabel metal2 s 2016 43200 2128 44000 0 FreeSans 448 90 0 0 chanx_left_out[14]
port 27 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chanx_left_out[15]
port 28 nsew signal tristate
flabel metal2 s 9408 43200 9520 44000 0 FreeSans 448 90 0 0 chanx_left_out[16]
port 29 nsew signal tristate
flabel metal2 s 2688 43200 2800 44000 0 FreeSans 448 90 0 0 chanx_left_out[17]
port 30 nsew signal tristate
flabel metal3 s 0 9408 800 9520 0 FreeSans 448 0 0 0 chanx_left_out[18]
port 31 nsew signal tristate
flabel metal2 s 8736 43200 8848 44000 0 FreeSans 448 90 0 0 chanx_left_out[19]
port 32 nsew signal tristate
flabel metal2 s 4032 43200 4144 44000 0 FreeSans 448 90 0 0 chanx_left_out[1]
port 33 nsew signal tristate
flabel metal2 s 5376 43200 5488 44000 0 FreeSans 448 90 0 0 chanx_left_out[2]
port 34 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 chanx_left_out[3]
port 35 nsew signal tristate
flabel metal2 s 20832 43200 20944 44000 0 FreeSans 448 90 0 0 chanx_left_out[4]
port 36 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 chanx_left_out[5]
port 37 nsew signal tristate
flabel metal2 s 15456 43200 15568 44000 0 FreeSans 448 90 0 0 chanx_left_out[6]
port 38 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 chanx_left_out[7]
port 39 nsew signal tristate
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 chanx_left_out[8]
port 40 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 chanx_left_out[9]
port 41 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 chanx_right_in[0]
port 42 nsew signal input
flabel metal2 s 26208 43200 26320 44000 0 FreeSans 448 90 0 0 chanx_right_in[10]
port 43 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 chanx_right_in[11]
port 44 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 chanx_right_in[12]
port 45 nsew signal input
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 chanx_right_in[13]
port 46 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chanx_right_in[14]
port 47 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 chanx_right_in[15]
port 48 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 chanx_right_in[16]
port 49 nsew signal input
flabel metal3 s 0 672 800 784 0 FreeSans 448 0 0 0 chanx_right_in[17]
port 50 nsew signal input
flabel metal2 s 25536 43200 25648 44000 0 FreeSans 448 90 0 0 chanx_right_in[18]
port 51 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 chanx_right_in[19]
port 52 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 chanx_right_in[1]
port 53 nsew signal input
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 chanx_right_in[2]
port 54 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 chanx_right_in[3]
port 55 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 chanx_right_in[4]
port 56 nsew signal input
flabel metal2 s 18816 43200 18928 44000 0 FreeSans 448 90 0 0 chanx_right_in[5]
port 57 nsew signal input
flabel metal3 s 0 2688 800 2800 0 FreeSans 448 0 0 0 chanx_right_in[6]
port 58 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 chanx_right_in[7]
port 59 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 chanx_right_in[8]
port 60 nsew signal input
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 chanx_right_in[9]
port 61 nsew signal input
flabel metal2 s 13440 43200 13552 44000 0 FreeSans 448 90 0 0 chanx_right_out[0]
port 62 nsew signal tristate
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 chanx_right_out[10]
port 63 nsew signal tristate
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 chanx_right_out[11]
port 64 nsew signal tristate
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 chanx_right_out[12]
port 65 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 chanx_right_out[13]
port 66 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 chanx_right_out[14]
port 67 nsew signal tristate
flabel metal2 s 10080 43200 10192 44000 0 FreeSans 448 90 0 0 chanx_right_out[15]
port 68 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 chanx_right_out[16]
port 69 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 chanx_right_out[17]
port 70 nsew signal tristate
flabel metal2 s 8064 43200 8176 44000 0 FreeSans 448 90 0 0 chanx_right_out[18]
port 71 nsew signal tristate
flabel metal2 s 1344 43200 1456 44000 0 FreeSans 448 90 0 0 chanx_right_out[19]
port 72 nsew signal tristate
flabel metal2 s 16128 43200 16240 44000 0 FreeSans 448 90 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal2 s 24864 43200 24976 44000 0 FreeSans 448 90 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal2 s 22176 43200 22288 44000 0 FreeSans 448 90 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 3360 43200 3472 44000 0 FreeSans 448 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal2 s 20160 43200 20272 44000 0 FreeSans 448 90 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 chany_top_in[0]
port 82 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chany_top_in[10]
port 83 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 chany_top_in[11]
port 84 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chany_top_in[12]
port 85 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chany_top_in[13]
port 86 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 chany_top_in[14]
port 87 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 chany_top_in[15]
port 88 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 chany_top_in[16]
port 89 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 chany_top_in[17]
port 90 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chany_top_in[18]
port 91 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chany_top_in[19]
port 92 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chany_top_in[1]
port 93 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 chany_top_in[2]
port 94 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chany_top_in[3]
port 95 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 chany_top_in[4]
port 96 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chany_top_in[5]
port 97 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 chany_top_in[6]
port 98 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chany_top_in[7]
port 99 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 chany_top_in[8]
port 100 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chany_top_in[9]
port 101 nsew signal input
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 chany_top_out[0]
port 102 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 chany_top_out[10]
port 103 nsew signal tristate
flabel metal2 s 14784 43200 14896 44000 0 FreeSans 448 90 0 0 chany_top_out[11]
port 104 nsew signal tristate
flabel metal2 s 672 43200 784 44000 0 FreeSans 448 90 0 0 chany_top_out[12]
port 105 nsew signal tristate
flabel metal2 s 12768 43200 12880 44000 0 FreeSans 448 90 0 0 chany_top_out[13]
port 106 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 chany_top_out[14]
port 107 nsew signal tristate
flabel metal2 s 4704 43200 4816 44000 0 FreeSans 448 90 0 0 chany_top_out[15]
port 108 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 chany_top_out[16]
port 109 nsew signal tristate
flabel metal2 s 18144 43200 18256 44000 0 FreeSans 448 90 0 0 chany_top_out[17]
port 110 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 chany_top_out[18]
port 111 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 chany_top_out[19]
port 112 nsew signal tristate
flabel metal2 s 6048 43200 6160 44000 0 FreeSans 448 90 0 0 chany_top_out[1]
port 113 nsew signal tristate
flabel metal2 s 14112 43200 14224 44000 0 FreeSans 448 90 0 0 chany_top_out[2]
port 114 nsew signal tristate
flabel metal2 s 12096 43200 12208 44000 0 FreeSans 448 90 0 0 chany_top_out[3]
port 115 nsew signal tristate
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chany_top_out[4]
port 116 nsew signal tristate
flabel metal2 s 11424 43200 11536 44000 0 FreeSans 448 90 0 0 chany_top_out[5]
port 117 nsew signal tristate
flabel metal2 s 10752 43200 10864 44000 0 FreeSans 448 90 0 0 chany_top_out[6]
port 118 nsew signal tristate
flabel metal2 s 17472 43200 17584 44000 0 FreeSans 448 90 0 0 chany_top_out[7]
port 119 nsew signal tristate
flabel metal2 s 22848 43200 22960 44000 0 FreeSans 448 90 0 0 chany_top_out[8]
port 120 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chany_top_out[9]
port 121 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 122 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 123 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 124 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 125 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 126 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 127 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 pReset
port 128 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 prog_clk
port 129 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 131 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 132 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 133 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 134 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 135 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 136 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 137 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 138 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 139 nsew signal input
flabel metal4 s 4448 3076 4768 40828 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 35168 3076 35488 40828 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 19808 3076 20128 40828 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
rlabel metal1 21952 39984 21952 39984 0 vdd
rlabel metal1 21952 40768 21952 40768 0 vss
rlabel metal2 7784 19208 7784 19208 0 _000_
rlabel metal2 8904 18816 8904 18816 0 _001_
rlabel metal2 3920 18648 3920 18648 0 _002_
rlabel metal2 5936 20216 5936 20216 0 _003_
rlabel metal3 2968 21672 2968 21672 0 _004_
rlabel metal2 3640 20944 3640 20944 0 _005_
rlabel metal2 7448 15960 7448 15960 0 _006_
rlabel metal2 4200 13328 4200 13328 0 _007_
rlabel metal2 2296 16128 2296 16128 0 _008_
rlabel metal2 2184 17248 2184 17248 0 _009_
rlabel metal2 13272 18256 13272 18256 0 _010_
rlabel metal2 12488 16856 12488 16856 0 _011_
rlabel metal2 14392 10360 14392 10360 0 _012_
rlabel metal2 12264 10248 12264 10248 0 _013_
rlabel metal2 10920 8260 10920 8260 0 _014_
rlabel metal2 8344 11536 8344 11536 0 _015_
rlabel metal3 7336 12712 7336 12712 0 _016_
rlabel metal2 9576 13328 9576 13328 0 _017_
rlabel metal2 14952 12544 14952 12544 0 _018_
rlabel metal2 10136 11816 10136 11816 0 _019_
rlabel metal2 21224 11536 21224 11536 0 _020_
rlabel metal2 21560 11816 21560 11816 0 _021_
rlabel metal2 17192 11368 17192 11368 0 _022_
rlabel metal2 17752 9352 17752 9352 0 _023_
rlabel metal2 18536 14728 18536 14728 0 _024_
rlabel metal2 16520 13944 16520 13944 0 _025_
rlabel metal2 22008 16632 22008 16632 0 _026_
rlabel metal2 20216 14112 20216 14112 0 _027_
rlabel metal2 23240 13496 23240 13496 0 _028_
rlabel metal2 21336 15120 21336 15120 0 _029_
rlabel metal2 25928 11928 25928 11928 0 _030_
rlabel metal3 27272 12712 27272 12712 0 _031_
rlabel metal2 30072 9968 30072 9968 0 _032_
rlabel metal2 28504 10864 28504 10864 0 _033_
rlabel metal2 33208 10976 33208 10976 0 _034_
rlabel metal2 29512 13328 29512 13328 0 _035_
rlabel metal2 27720 20356 27720 20356 0 _036_
rlabel metal2 26264 17080 26264 17080 0 _037_
rlabel metal2 29848 18144 29848 18144 0 _038_
rlabel metal2 29736 18144 29736 18144 0 _039_
rlabel metal2 37128 11984 37128 11984 0 _040_
rlabel metal2 33320 13104 33320 13104 0 _041_
rlabel metal2 39424 12376 39424 12376 0 _042_
rlabel metal2 37688 14224 37688 14224 0 _043_
rlabel metal3 34888 15848 34888 15848 0 _044_
rlabel metal2 37912 16688 37912 16688 0 _045_
rlabel metal2 35896 19264 35896 19264 0 _046_
rlabel metal2 36120 17136 36120 17136 0 _047_
rlabel metal2 33768 20384 33768 20384 0 _048_
rlabel metal3 32648 21784 32648 21784 0 _049_
rlabel metal3 28952 22120 28952 22120 0 _050_
rlabel metal2 28056 21952 28056 21952 0 _051_
rlabel metal2 25592 21112 25592 21112 0 _052_
rlabel metal2 21784 21952 21784 21952 0 _053_
rlabel metal3 22400 21112 22400 21112 0 _054_
rlabel metal2 17864 18704 17864 18704 0 _055_
rlabel metal2 25816 26656 25816 26656 0 _056_
rlabel metal2 25928 25088 25928 25088 0 _057_
rlabel metal2 22456 26040 22456 26040 0 _058_
rlabel metal2 22344 25872 22344 25872 0 _059_
rlabel metal3 34104 25368 34104 25368 0 _060_
rlabel metal2 33544 24920 33544 24920 0 _061_
rlabel metal2 32200 25032 32200 25032 0 _062_
rlabel metal2 29848 26880 29848 26880 0 _063_
rlabel metal2 36904 27216 36904 27216 0 _064_
rlabel metal2 39368 25032 39368 25032 0 _065_
rlabel metal2 37800 23128 37800 23128 0 _066_
rlabel metal2 39256 22568 39256 22568 0 _067_
rlabel metal3 37968 21784 37968 21784 0 _068_
rlabel metal2 35784 22624 35784 22624 0 _069_
rlabel metal3 36120 31864 36120 31864 0 _070_
rlabel metal2 35784 30912 35784 30912 0 _071_
rlabel metal2 33656 31556 33656 31556 0 _072_
rlabel metal2 37576 29792 37576 29792 0 _073_
rlabel metal2 39872 30072 39872 30072 0 _074_
rlabel metal3 38808 28392 38808 28392 0 _075_
rlabel metal2 31864 29792 31864 29792 0 _076_
rlabel metal2 31416 31920 31416 31920 0 _077_
rlabel metal2 29848 31164 29848 31164 0 _078_
rlabel metal2 28560 31192 28560 31192 0 _079_
rlabel metal2 26264 32032 26264 32032 0 _080_
rlabel metal2 24248 31556 24248 31556 0 _081_
rlabel metal2 27272 28280 27272 28280 0 _082_
rlabel metal2 25200 27944 25200 27944 0 _083_
rlabel metal2 23576 29568 23576 29568 0 _084_
rlabel metal2 20328 30016 20328 30016 0 _085_
rlabel metal3 18984 28728 18984 28728 0 _086_
rlabel metal3 19376 31528 19376 31528 0 _087_
rlabel metal2 19432 30800 19432 30800 0 _088_
rlabel metal2 16520 28952 16520 28952 0 _089_
rlabel metal2 15064 29736 15064 29736 0 _090_
rlabel metal2 12376 29232 12376 29232 0 _091_
rlabel metal3 8372 26488 8372 26488 0 _092_
rlabel metal3 7448 27048 7448 27048 0 _093_
rlabel metal2 13720 29176 13720 29176 0 _094_
rlabel metal2 10024 28112 10024 28112 0 _095_
rlabel metal2 10696 30408 10696 30408 0 _096_
rlabel metal2 8736 28392 8736 28392 0 _097_
rlabel metal2 8344 30240 8344 30240 0 _098_
rlabel metal3 6440 28952 6440 28952 0 _099_
rlabel metal2 16632 21168 16632 21168 0 _100_
rlabel metal2 16296 21840 16296 21840 0 _101_
rlabel metal2 14616 22848 14616 22848 0 _102_
rlabel metal2 19432 24192 19432 24192 0 _103_
rlabel metal2 17416 24864 17416 24864 0 _104_
rlabel metal3 20188 26376 20188 26376 0 _105_
rlabel metal2 20776 23576 20776 23576 0 _106_
rlabel metal2 16184 22512 16184 22512 0 _107_
rlabel metal2 16296 24584 16296 24584 0 _108_
rlabel metal2 12488 22176 12488 22176 0 _109_
rlabel metal2 10248 22232 10248 22232 0 _110_
rlabel metal2 8232 22904 8232 22904 0 _111_
rlabel metal2 16184 27440 16184 27440 0 _112_
rlabel metal2 26152 27328 26152 27328 0 _113_
rlabel metal3 5152 20328 5152 20328 0 _114_
rlabel metal2 13888 16072 13888 16072 0 _115_
rlabel metal2 22624 12936 22624 12936 0 _116_
rlabel metal3 30016 9800 30016 9800 0 _117_
rlabel metal2 33600 21560 33600 21560 0 _118_
rlabel metal3 21056 22344 21056 22344 0 _119_
rlabel metal2 30240 23688 30240 23688 0 _120_
rlabel metal2 29624 29120 29624 29120 0 _121_
rlabel metal2 25592 28280 25592 28280 0 _122_
rlabel metal2 7336 26208 7336 26208 0 _123_
rlabel metal2 20440 25144 20440 25144 0 _124_
rlabel metal2 1736 20832 1736 20832 0 ccff_head
rlabel metal2 27608 41496 27608 41496 0 ccff_tail
rlabel metal2 22008 40712 22008 40712 0 chanx_left_in[0]
rlabel metal2 3024 3416 3024 3416 0 chanx_left_in[10]
rlabel metal2 1736 22624 1736 22624 0 chanx_left_in[11]
rlabel metal2 1736 35336 1736 35336 0 chanx_left_in[12]
rlabel metal3 2534 43736 2534 43736 0 chanx_left_in[13]
rlabel metal2 17304 40712 17304 40712 0 chanx_left_in[14]
rlabel metal2 21000 40488 21000 40488 0 chanx_left_in[15]
rlabel metal2 3864 3192 3864 3192 0 chanx_left_in[16]
rlabel metal2 56 41706 56 41706 0 chanx_left_in[17]
rlabel metal2 1736 37576 1736 37576 0 chanx_left_in[18]
rlabel metal2 2408 30240 2408 30240 0 chanx_left_in[19]
rlabel metal2 1848 25872 1848 25872 0 chanx_left_in[1]
rlabel metal2 6888 39592 6888 39592 0 chanx_left_in[2]
rlabel metal2 7896 39368 7896 39368 0 chanx_left_in[4]
rlabel metal2 24024 40152 24024 40152 0 chanx_left_in[5]
rlabel metal3 3024 36456 3024 36456 0 chanx_left_in[6]
rlabel metal3 2058 38360 2058 38360 0 chanx_left_in[8]
rlabel metal3 3304 4424 3304 4424 0 chanx_left_in[9]
rlabel metal3 1358 24248 1358 24248 0 chanx_left_out[10]
rlabel metal2 24920 40264 24920 40264 0 chanx_left_out[11]
rlabel metal3 1414 34328 1414 34328 0 chanx_left_out[13]
rlabel metal2 2520 40600 2520 40600 0 chanx_left_out[14]
rlabel metal2 10808 854 10808 854 0 chanx_left_out[15]
rlabel metal2 2744 41762 2744 41762 0 chanx_left_out[17]
rlabel metal3 1414 9464 1414 9464 0 chanx_left_out[18]
rlabel metal2 9352 39704 9352 39704 0 chanx_left_out[19]
rlabel metal2 4088 41874 4088 41874 0 chanx_left_out[1]
rlabel metal2 5992 40768 5992 40768 0 chanx_left_out[2]
rlabel metal3 1358 5432 1358 5432 0 chanx_left_out[3]
rlabel metal2 7448 854 7448 854 0 chanx_left_out[5]
rlabel metal2 16072 40880 16072 40880 0 chanx_left_out[6]
rlabel metal3 1358 6776 1358 6776 0 chanx_left_out[7]
rlabel metal3 1358 31640 1358 31640 0 chanx_left_out[9]
rlabel metal2 1736 29176 1736 29176 0 chanx_right_in[0]
rlabel metal2 26712 40040 26712 40040 0 chanx_right_in[10]
rlabel metal2 1736 23688 1736 23688 0 chanx_right_in[12]
rlabel metal2 1736 33096 1736 33096 0 chanx_right_in[13]
rlabel metal2 10136 2086 10136 2086 0 chanx_right_in[14]
rlabel metal2 1736 28448 1736 28448 0 chanx_right_in[16]
rlabel metal2 2408 2072 2408 2072 0 chanx_right_in[17]
rlabel metal2 25592 41482 25592 41482 0 chanx_right_in[18]
rlabel metal3 1582 36344 1582 36344 0 chanx_right_in[1]
rlabel metal2 1736 3864 1736 3864 0 chanx_right_in[2]
rlabel metal2 6104 2086 6104 2086 0 chanx_right_in[4]
rlabel metal2 18872 41482 18872 41482 0 chanx_right_in[5]
rlabel metal2 3976 3136 3976 3136 0 chanx_right_in[6]
rlabel metal2 3640 36400 3640 36400 0 chanx_right_in[8]
rlabel metal2 1736 29848 1736 29848 0 chanx_right_in[9]
rlabel metal3 1414 8120 1414 8120 0 chanx_right_out[10]
rlabel metal3 1358 8792 1358 8792 0 chanx_right_out[11]
rlabel metal3 1526 26936 1526 26936 0 chanx_right_out[13]
rlabel metal2 2128 38248 2128 38248 0 chanx_right_out[14]
rlabel metal2 11256 41160 11256 41160 0 chanx_right_out[15]
rlabel metal3 1414 6104 1414 6104 0 chanx_right_out[17]
rlabel metal2 7896 41104 7896 41104 0 chanx_right_out[18]
rlabel metal3 1792 39032 1792 39032 0 chanx_right_out[19]
rlabel metal2 16856 39760 16856 39760 0 chanx_right_out[1]
rlabel metal3 1414 30968 1414 30968 0 chanx_right_out[2]
rlabel metal3 25872 40264 25872 40264 0 chanx_right_out[3]
rlabel metal3 2254 41720 2254 41720 0 chanx_right_out[5]
rlabel metal2 23352 40768 23352 40768 0 chanx_right_out[6]
rlabel metal2 4088 40040 4088 40040 0 chanx_right_out[7]
rlabel metal3 1358 43064 1358 43064 0 chanx_right_out[9]
rlabel metal3 1470 24920 1470 24920 0 chany_top_out[16]
rlabel metal3 18704 40600 18704 40600 0 chany_top_out[17]
rlabel metal3 1470 26264 1470 26264 0 chany_top_out[18]
rlabel metal2 27272 25928 27272 25928 0 clknet_0_prog_clk
rlabel metal2 6328 18088 6328 18088 0 clknet_3_0__leaf_prog_clk
rlabel metal2 20888 18032 20888 18032 0 clknet_3_1__leaf_prog_clk
rlabel metal3 3752 21560 3752 21560 0 clknet_3_2__leaf_prog_clk
rlabel metal3 18760 29288 18760 29288 0 clknet_3_3__leaf_prog_clk
rlabel metal2 24472 21056 24472 21056 0 clknet_3_4__leaf_prog_clk
rlabel via2 30072 12152 30072 12152 0 clknet_3_5__leaf_prog_clk
rlabel metal2 26824 25872 26824 25872 0 clknet_3_6__leaf_prog_clk
rlabel metal2 30912 23912 30912 23912 0 clknet_3_7__leaf_prog_clk
rlabel metal3 29876 28392 29876 28392 0 mem_left_track_1.DFFR_0_.D
rlabel metal2 29064 27888 29064 27888 0 mem_left_track_1.DFFR_0_.Q
rlabel metal3 34048 24808 34048 24808 0 mem_left_track_1.DFFR_1_.Q
rlabel metal3 36120 24136 36120 24136 0 mem_left_track_1.DFFR_2_.Q
rlabel metal2 30184 25032 30184 25032 0 mem_left_track_1.DFFR_3_.Q
rlabel metal2 23240 23800 23240 23800 0 mem_left_track_1.DFFR_4_.Q
rlabel metal3 25368 23800 25368 23800 0 mem_left_track_1.DFFR_5_.Q
rlabel metal2 26488 26544 26488 26544 0 mem_left_track_1.DFFR_6_.Q
rlabel metal2 25032 27608 25032 27608 0 mem_left_track_1.DFFR_7_.Q
rlabel metal2 16016 28840 16016 28840 0 mem_left_track_17.DFFR_0_.D
rlabel metal2 4984 31920 4984 31920 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 9128 31416 9128 31416 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 9240 29792 9240 29792 0 mem_left_track_17.DFFR_2_.Q
rlabel metal2 9912 28168 9912 28168 0 mem_left_track_17.DFFR_3_.Q
rlabel metal2 10584 26600 10584 26600 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 15960 31584 15960 31584 0 mem_left_track_17.DFFR_5_.Q
rlabel metal2 16184 28784 16184 28784 0 mem_left_track_25.DFFR_0_.Q
rlabel metal3 18200 26376 18200 26376 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 20216 21840 20216 21840 0 mem_left_track_25.DFFR_2_.Q
rlabel metal2 11816 22568 11816 22568 0 mem_left_track_25.DFFR_3_.Q
rlabel metal2 16968 21000 16968 21000 0 mem_left_track_25.DFFR_4_.Q
rlabel metal2 15736 22736 15736 22736 0 mem_left_track_25.DFFR_5_.Q
rlabel metal2 7000 23464 7000 23464 0 mem_left_track_33.DFFR_0_.Q
rlabel metal2 8120 24528 8120 24528 0 mem_left_track_33.DFFR_1_.Q
rlabel metal2 7000 21840 7000 21840 0 mem_left_track_33.DFFR_2_.Q
rlabel metal2 19376 15400 19376 15400 0 mem_left_track_33.DFFR_3_.Q
rlabel metal2 17976 21000 17976 21000 0 mem_left_track_33.DFFR_4_.Q
rlabel metal3 6664 26936 6664 26936 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 9128 28728 9128 28728 0 mem_left_track_9.DFFR_1_.Q
rlabel metal2 13048 30240 13048 30240 0 mem_left_track_9.DFFR_2_.Q
rlabel metal2 15736 33208 15736 33208 0 mem_left_track_9.DFFR_3_.Q
rlabel metal2 17080 31696 17080 31696 0 mem_left_track_9.DFFR_4_.Q
rlabel metal3 26824 18536 26824 18536 0 mem_right_track_0.DFFR_0_.D
rlabel metal2 19544 18760 19544 18760 0 mem_right_track_0.DFFR_0_.Q
rlabel metal3 26040 19096 26040 19096 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 21000 22512 21000 22512 0 mem_right_track_0.DFFR_2_.Q
rlabel metal3 35112 22400 35112 22400 0 mem_right_track_0.DFFR_3_.Q
rlabel metal2 28840 20216 28840 20216 0 mem_right_track_0.DFFR_4_.Q
rlabel metal2 29064 22064 29064 22064 0 mem_right_track_0.DFFR_5_.Q
rlabel metal2 39032 21000 39032 21000 0 mem_right_track_0.DFFR_6_.Q
rlabel metal2 34440 23968 34440 23968 0 mem_right_track_0.DFFR_7_.Q
rlabel metal2 37744 28056 37744 28056 0 mem_right_track_16.DFFR_0_.D
rlabel metal2 36904 29624 36904 29624 0 mem_right_track_16.DFFR_0_.Q
rlabel metal2 41216 36344 41216 36344 0 mem_right_track_16.DFFR_1_.Q
rlabel metal2 36792 29960 36792 29960 0 mem_right_track_16.DFFR_2_.Q
rlabel metal3 34328 33096 34328 33096 0 mem_right_track_16.DFFR_3_.Q
rlabel metal3 36960 33096 36960 33096 0 mem_right_track_16.DFFR_4_.Q
rlabel metal2 31864 31696 31864 31696 0 mem_right_track_16.DFFR_5_.Q
rlabel metal3 26040 33544 26040 33544 0 mem_right_track_24.DFFR_0_.Q
rlabel metal2 27048 32592 27048 32592 0 mem_right_track_24.DFFR_1_.Q
rlabel metal3 30296 32872 30296 32872 0 mem_right_track_24.DFFR_2_.Q
rlabel metal2 30520 32984 30520 32984 0 mem_right_track_24.DFFR_3_.Q
rlabel metal2 32760 30520 32760 30520 0 mem_right_track_24.DFFR_4_.Q
rlabel metal2 30296 30688 30296 30688 0 mem_right_track_24.DFFR_5_.Q
rlabel metal3 19656 32648 19656 32648 0 mem_right_track_32.DFFR_0_.Q
rlabel metal3 18536 33096 18536 33096 0 mem_right_track_32.DFFR_1_.Q
rlabel metal3 22232 28504 22232 28504 0 mem_right_track_32.DFFR_2_.Q
rlabel metal3 25704 29400 25704 29400 0 mem_right_track_32.DFFR_3_.Q
rlabel metal3 26936 30072 26936 30072 0 mem_right_track_32.DFFR_4_.Q
rlabel metal3 37800 17528 37800 17528 0 mem_right_track_8.DFFR_0_.Q
rlabel metal2 38136 20748 38136 20748 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 39816 24024 39816 24024 0 mem_right_track_8.DFFR_2_.Q
rlabel metal2 37016 24976 37016 24976 0 mem_right_track_8.DFFR_3_.Q
rlabel metal3 40096 25704 40096 25704 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 5320 22288 5320 22288 0 mem_top_track_0.DFFR_0_.Q
rlabel metal3 2184 20664 2184 20664 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 3080 18872 3080 18872 0 mem_top_track_0.DFFR_2_.Q
rlabel metal2 5096 19432 5096 19432 0 mem_top_track_0.DFFR_3_.Q
rlabel metal2 10528 15960 10528 15960 0 mem_top_track_0.DFFR_4_.Q
rlabel metal2 7112 18256 7112 18256 0 mem_top_track_0.DFFR_5_.Q
rlabel metal2 19712 12264 19712 12264 0 mem_top_track_10.DFFR_0_.D
rlabel metal2 20664 13160 20664 13160 0 mem_top_track_10.DFFR_0_.Q
rlabel metal2 25480 15512 25480 15512 0 mem_top_track_10.DFFR_1_.Q
rlabel metal2 23576 13216 23576 13216 0 mem_top_track_12.DFFR_0_.Q
rlabel metal2 27048 12208 27048 12208 0 mem_top_track_12.DFFR_1_.Q
rlabel metal2 27384 13496 27384 13496 0 mem_top_track_14.DFFR_0_.Q
rlabel metal3 25704 10696 25704 10696 0 mem_top_track_14.DFFR_1_.Q
rlabel metal2 29848 14168 29848 14168 0 mem_top_track_16.DFFR_0_.Q
rlabel metal3 33880 12824 33880 12824 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 29512 10696 29512 10696 0 mem_top_track_18.DFFR_0_.Q
rlabel metal3 34384 11144 34384 11144 0 mem_top_track_18.DFFR_1_.Q
rlabel metal3 11704 17864 11704 17864 0 mem_top_track_2.DFFR_0_.Q
rlabel metal2 8904 17584 8904 17584 0 mem_top_track_2.DFFR_1_.Q
rlabel metal2 1960 16016 1960 16016 0 mem_top_track_2.DFFR_2_.Q
rlabel metal2 1624 14168 1624 14168 0 mem_top_track_2.DFFR_3_.Q
rlabel metal3 4312 15960 4312 15960 0 mem_top_track_2.DFFR_4_.Q
rlabel metal2 8456 14448 8456 14448 0 mem_top_track_2.DFFR_5_.Q
rlabel metal2 37912 11368 37912 11368 0 mem_top_track_20.DFFR_0_.Q
rlabel metal2 39144 10248 39144 10248 0 mem_top_track_20.DFFR_1_.Q
rlabel metal2 39368 13104 39368 13104 0 mem_top_track_22.DFFR_0_.Q
rlabel metal2 41720 13160 41720 13160 0 mem_top_track_22.DFFR_1_.Q
rlabel metal2 36344 14784 36344 14784 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 35056 15400 35056 15400 0 mem_top_track_24.DFFR_1_.Q
rlabel metal2 37800 13888 37800 13888 0 mem_top_track_26.DFFR_0_.Q
rlabel metal2 32088 15456 32088 15456 0 mem_top_track_26.DFFR_1_.Q
rlabel metal2 28728 15624 28728 15624 0 mem_top_track_28.DFFR_0_.Q
rlabel metal3 29960 16968 29960 16968 0 mem_top_track_28.DFFR_1_.Q
rlabel metal2 39032 19432 39032 19432 0 mem_top_track_38.DFFR_0_.Q
rlabel metal3 11256 14392 11256 14392 0 mem_top_track_4.DFFR_0_.Q
rlabel metal2 7224 11984 7224 11984 0 mem_top_track_4.DFFR_1_.Q
rlabel metal3 10360 10696 10360 10696 0 mem_top_track_4.DFFR_2_.Q
rlabel metal3 12376 9128 12376 9128 0 mem_top_track_4.DFFR_3_.Q
rlabel metal3 13720 7560 13720 7560 0 mem_top_track_4.DFFR_4_.Q
rlabel metal3 16744 9352 16744 9352 0 mem_top_track_4.DFFR_5_.Q
rlabel metal2 18424 8260 18424 8260 0 mem_top_track_6.DFFR_0_.Q
rlabel metal2 22008 10136 22008 10136 0 mem_top_track_6.DFFR_1_.Q
rlabel metal2 23240 9856 23240 9856 0 mem_top_track_6.DFFR_2_.Q
rlabel metal2 20440 10528 20440 10528 0 mem_top_track_6.DFFR_3_.Q
rlabel metal2 9352 12376 9352 12376 0 mem_top_track_6.DFFR_4_.Q
rlabel metal2 15960 11592 15960 11592 0 mem_top_track_6.DFFR_5_.Q
rlabel metal2 17528 13160 17528 13160 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 2072 21112 2072 21112 0 net1
rlabel metal2 8736 38808 8736 38808 0 net10
rlabel metal2 33544 22960 33544 22960 0 net100
rlabel metal3 37520 21896 37520 21896 0 net101
rlabel metal2 29736 13776 29736 13776 0 net102
rlabel metal2 32200 19264 32200 19264 0 net103
rlabel metal2 32200 27888 32200 27888 0 net104
rlabel metal2 7336 20048 7336 20048 0 net105
rlabel metal2 21112 29232 21112 29232 0 net106
rlabel metal2 13216 10584 13216 10584 0 net107
rlabel metal2 21784 13160 21784 13160 0 net108
rlabel metal2 23352 22680 23352 22680 0 net109
rlabel metal2 2072 37184 2072 37184 0 net11
rlabel metal3 18312 31080 18312 31080 0 net110
rlabel metal2 20496 30968 20496 30968 0 net111
rlabel metal2 11816 26516 11816 26516 0 net112
rlabel metal2 20776 18760 20776 18760 0 net113
rlabel metal2 24360 12208 24360 12208 0 net114
rlabel metal3 25816 21616 25816 21616 0 net115
rlabel metal2 11368 18368 11368 18368 0 net116
rlabel metal2 23688 14952 23688 14952 0 net117
rlabel metal2 14056 31808 14056 31808 0 net118
rlabel metal2 23464 11592 23464 11592 0 net119
rlabel metal2 2744 30408 2744 30408 0 net12
rlabel metal2 13160 28952 13160 28952 0 net120
rlabel metal2 11816 17696 11816 17696 0 net121
rlabel metal3 8204 21448 8204 21448 0 net122
rlabel metal2 11256 27384 11256 27384 0 net123
rlabel metal3 38024 20832 38024 20832 0 net124
rlabel metal3 36512 19992 36512 19992 0 net125
rlabel metal2 40040 16072 40040 16072 0 net126
rlabel metal2 4088 15736 4088 15736 0 net127
rlabel metal2 33376 31752 33376 31752 0 net128
rlabel metal2 38024 22008 38024 22008 0 net129
rlabel metal2 3584 37912 3584 37912 0 net13
rlabel metal2 9240 25592 9240 25592 0 net130
rlabel metal2 12040 13384 12040 13384 0 net131
rlabel metal2 37464 14672 37464 14672 0 net132
rlabel metal3 4984 18872 4984 18872 0 net133
rlabel metal3 40264 29400 40264 29400 0 net134
rlabel metal2 32088 12600 32088 12600 0 net135
rlabel metal3 26768 33432 26768 33432 0 net136
rlabel metal2 16296 8372 16296 8372 0 net137
rlabel metal2 16296 13776 16296 13776 0 net138
rlabel metal2 37576 33264 37576 33264 0 net139
rlabel metal2 7224 39368 7224 39368 0 net14
rlabel metal2 9856 28616 9856 28616 0 net140
rlabel metal2 29624 32592 29624 32592 0 net141
rlabel metal3 25144 32984 25144 32984 0 net142
rlabel metal2 28280 12880 28280 12880 0 net143
rlabel metal2 21000 9464 21000 9464 0 net144
rlabel metal2 10360 13888 10360 13888 0 net145
rlabel metal2 6104 11816 6104 11816 0 net146
rlabel metal2 37800 26600 37800 26600 0 net147
rlabel metal2 23352 24752 23352 24752 0 net148
rlabel metal2 7112 14056 7112 14056 0 net149
rlabel metal3 6328 38696 6328 38696 0 net15
rlabel metal2 29736 26264 29736 26264 0 net150
rlabel metal2 4760 16800 4760 16800 0 net151
rlabel metal2 6104 27496 6104 27496 0 net152
rlabel metal2 37744 30184 37744 30184 0 net153
rlabel metal2 36120 30912 36120 30912 0 net154
rlabel metal2 18760 28616 18760 28616 0 net155
rlabel metal2 4760 23464 4760 23464 0 net156
rlabel metal2 17976 13328 17976 13328 0 net157
rlabel metal2 25816 16016 25816 16016 0 net158
rlabel metal2 22792 29960 22792 29960 0 net159
rlabel metal2 23800 38640 23800 38640 0 net16
rlabel metal2 15288 23184 15288 23184 0 net160
rlabel metal2 30744 10920 30744 10920 0 net161
rlabel metal2 33656 12600 33656 12600 0 net162
rlabel metal2 6104 30128 6104 30128 0 net163
rlabel metal2 8232 31024 8232 31024 0 net164
rlabel metal2 17248 23912 17248 23912 0 net165
rlabel metal3 6104 19320 6104 19320 0 net166
rlabel metal3 8260 17752 8260 17752 0 net167
rlabel metal2 24808 29456 24808 29456 0 net168
rlabel metal2 31976 15344 31976 15344 0 net169
rlabel metal2 4816 36344 4816 36344 0 net17
rlabel metal2 12376 10696 12376 10696 0 net170
rlabel metal2 40264 23912 40264 23912 0 net171
rlabel metal2 19544 8372 19544 8372 0 net172
rlabel metal2 31304 24080 31304 24080 0 net173
rlabel metal2 40040 30268 40040 30268 0 net174
rlabel metal2 18312 22008 18312 22008 0 net175
rlabel metal2 11928 31864 11928 31864 0 net176
rlabel metal2 36008 24976 36008 24976 0 net177
rlabel metal2 26824 13328 26824 13328 0 net178
rlabel metal2 33880 16016 33880 16016 0 net179
rlabel metal2 5320 37688 5320 37688 0 net18
rlabel metal2 10024 9576 10024 9576 0 net180
rlabel metal3 25088 19320 25088 19320 0 net181
rlabel metal2 13944 12600 13944 12600 0 net182
rlabel metal2 34776 11312 34776 11312 0 net183
rlabel metal2 27496 32760 27496 32760 0 net184
rlabel metal2 21560 25144 21560 25144 0 net185
rlabel metal2 6216 30016 6216 30016 0 net186
rlabel metal2 10584 24752 10584 24752 0 net187
rlabel metal2 8008 22344 8008 22344 0 net188
rlabel metal2 18424 28672 18424 28672 0 net189
rlabel metal2 2072 4816 2072 4816 0 net19
rlabel metal2 27832 18536 27832 18536 0 net190
rlabel metal2 19544 14952 19544 14952 0 net191
rlabel metal3 9632 9464 9632 9464 0 net192
rlabel metal2 13832 22232 13832 22232 0 net193
rlabel metal2 38136 18424 38136 18424 0 net194
rlabel metal2 40040 12208 40040 12208 0 net195
rlabel metal2 15064 32928 15064 32928 0 net196
rlabel metal2 34664 27496 34664 27496 0 net197
rlabel metal2 20328 18760 20328 18760 0 net198
rlabel metal2 13776 21560 13776 21560 0 net199
rlabel metal2 21784 39312 21784 39312 0 net2
rlabel metal2 2072 29736 2072 29736 0 net20
rlabel metal2 15008 23128 15008 23128 0 net200
rlabel metal2 3360 15176 3360 15176 0 net201
rlabel metal3 28840 24640 28840 24640 0 net202
rlabel metal2 3976 15344 3976 15344 0 net203
rlabel metal2 24024 15848 24024 15848 0 net204
rlabel metal2 21784 30912 21784 30912 0 net205
rlabel metal2 8568 26488 8568 26488 0 net206
rlabel metal2 24584 32592 24584 32592 0 net207
rlabel metal2 26488 39032 26488 39032 0 net21
rlabel metal3 3192 23800 3192 23800 0 net22
rlabel metal3 4648 33208 4648 33208 0 net23
rlabel metal2 10640 3416 10640 3416 0 net24
rlabel metal2 2072 28896 2072 28896 0 net25
rlabel metal2 2744 4312 2744 4312 0 net26
rlabel metal2 25816 38248 25816 38248 0 net27
rlabel metal2 2744 36736 2744 36736 0 net28
rlabel metal2 2128 3416 2128 3416 0 net29
rlabel metal2 3416 4648 3416 4648 0 net3
rlabel metal2 6664 4256 6664 4256 0 net30
rlabel metal2 19096 38864 19096 38864 0 net31
rlabel metal2 3752 4200 3752 4200 0 net32
rlabel metal2 3976 36232 3976 36232 0 net33
rlabel metal2 2072 30464 2072 30464 0 net34
rlabel metal2 14504 28224 14504 28224 0 net35
rlabel metal3 23912 23352 23912 23352 0 net36
rlabel metal3 4312 24696 4312 24696 0 net37
rlabel metal2 24584 39648 24584 39648 0 net38
rlabel metal2 2800 34888 2800 34888 0 net39
rlabel metal2 2072 22848 2072 22848 0 net4
rlabel metal2 6888 39200 6888 39200 0 net40
rlabel metal2 11032 4200 11032 4200 0 net41
rlabel metal2 5656 39928 5656 39928 0 net42
rlabel metal2 3640 6692 3640 6692 0 net43
rlabel metal2 9016 39004 9016 39004 0 net44
rlabel metal3 5992 38920 5992 38920 0 net45
rlabel metal2 6272 39144 6272 39144 0 net46
rlabel metal2 2632 5432 2632 5432 0 net47
rlabel metal2 7560 4200 7560 4200 0 net48
rlabel metal2 15176 39424 15176 39424 0 net49
rlabel metal2 2072 35952 2072 35952 0 net5
rlabel metal2 2968 6216 2968 6216 0 net50
rlabel metal2 6384 39368 6384 39368 0 net51
rlabel metal2 4312 5768 4312 5768 0 net52
rlabel metal2 3248 6104 3248 6104 0 net53
rlabel metal2 3024 26488 3024 26488 0 net54
rlabel metal2 2968 36344 2968 36344 0 net55
rlabel metal2 10360 39144 10360 39144 0 net56
rlabel metal2 2912 4536 2912 4536 0 net57
rlabel metal2 8736 39032 8736 39032 0 net58
rlabel metal3 3920 38920 3920 38920 0 net59
rlabel metal2 9464 39928 9464 39928 0 net6
rlabel metal3 13216 39368 13216 39368 0 net60
rlabel metal2 2744 31836 2744 31836 0 net61
rlabel metal2 26152 39480 26152 39480 0 net62
rlabel metal2 4368 38808 4368 38808 0 net63
rlabel metal2 22456 39200 22456 39200 0 net64
rlabel metal2 5544 39200 5544 39200 0 net65
rlabel metal2 4424 37632 4424 37632 0 net66
rlabel metal2 3080 25480 3080 25480 0 net67
rlabel metal2 18536 39088 18536 39088 0 net68
rlabel metal3 2856 34776 2856 34776 0 net69
rlabel metal3 13888 39144 13888 39144 0 net7
rlabel metal3 1246 33656 1246 33656 0 net70
rlabel metal3 3304 40600 3304 40600 0 net71
rlabel metal3 2030 7448 2030 7448 0 net72
rlabel metal2 13160 41272 13160 41272 0 net73
rlabel metal2 2464 35784 2464 35784 0 net74
rlabel metal2 14840 41930 14840 41930 0 net75
rlabel metal2 2184 34776 2184 34776 0 net76
rlabel metal2 12152 1246 12152 1246 0 net77
rlabel metal2 23128 40208 23128 40208 0 net78
rlabel metal2 17640 40600 17640 40600 0 net79
rlabel metal2 20776 39368 20776 39368 0 net8
rlabel metal2 10920 39480 10920 39480 0 net80
rlabel metal2 11928 41272 11928 41272 0 net81
rlabel metal2 8120 2030 8120 2030 0 net82
rlabel metal2 12264 40600 12264 40600 0 net83
rlabel metal2 14224 40600 14224 40600 0 net84
rlabel metal2 6104 40950 6104 40950 0 net85
rlabel metal3 1582 4088 1582 4088 0 net86
rlabel metal2 6776 2030 6776 2030 0 net87
rlabel metal3 2366 39704 2366 39704 0 net88
rlabel metal2 20440 40376 20440 40376 0 net89
rlabel metal2 3304 4480 3304 4480 0 net9
rlabel metal2 3304 34944 3304 34944 0 net90
rlabel metal2 13608 40600 13608 40600 0 net91
rlabel metal2 10584 39872 10584 39872 0 net92
rlabel metal3 1302 1400 1302 1400 0 net93
rlabel metal3 1246 32312 1246 32312 0 net94
rlabel metal2 20216 40768 20216 40768 0 net95
rlabel metal2 7504 39032 7504 39032 0 net96
rlabel metal2 33432 29960 33432 29960 0 net97
rlabel metal3 33096 21224 33096 21224 0 net98
rlabel metal2 28224 27048 28224 27048 0 net99
rlabel metal2 1736 27720 1736 27720 0 pReset
rlabel metal3 2814 22232 2814 22232 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 44000 44000
<< end >>
