magic
tech gf180mcuD
magscale 1 5
timestamp 1702149120
<< obsm1 >>
rect 672 1538 7360 6302
<< metal2 >>
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
<< obsm2 >>
rect 854 430 7346 6291
rect 854 350 2658 430
rect 2774 350 2994 430
rect 3110 350 3330 430
rect 3446 350 3666 430
rect 3782 350 4002 430
rect 4118 350 4338 430
rect 4454 350 7346 430
<< metal3 >>
rect 0 4704 400 4760
rect 7600 4704 8000 4760
rect 0 4368 400 4424
rect 7600 4368 8000 4424
rect 0 3696 400 3752
rect 7600 3696 8000 3752
rect 0 3360 400 3416
rect 7600 3360 8000 3416
rect 0 3024 400 3080
rect 7600 3024 8000 3080
<< obsm3 >>
rect 400 4790 7658 6286
rect 430 4674 7570 4790
rect 400 4454 7658 4674
rect 430 4338 7570 4454
rect 400 3782 7658 4338
rect 430 3666 7570 3782
rect 400 3446 7658 3666
rect 430 3330 7570 3446
rect 400 3110 7658 3330
rect 430 2994 7570 3110
rect 400 462 7658 2994
<< metal4 >>
rect 1418 1538 1578 6302
rect 2244 1538 2404 6302
rect 3070 1538 3230 6302
rect 3896 1538 4056 6302
rect 4722 1538 4882 6302
rect 5548 1538 5708 6302
rect 6374 1538 6534 6302
rect 7200 1538 7360 6302
<< labels >>
rlabel metal2 s 2688 0 2744 400 6 bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 1 nsew signal output
rlabel metal2 s 3024 0 3080 400 6 bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 2 nsew signal input
rlabel metal3 s 0 3696 400 3752 6 bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 3 nsew signal output
rlabel metal3 s 0 3024 400 3080 6 bottom_width_0_height_0_subtile_1__pin_outpad_0_
port 4 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 5 nsew signal output
rlabel metal2 s 3696 0 3752 400 6 bottom_width_0_height_0_subtile_2__pin_outpad_0_
port 6 nsew signal input
rlabel metal3 s 7600 3696 8000 3752 6 bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 7 nsew signal output
rlabel metal3 s 7600 3024 8000 3080 6 bottom_width_0_height_0_subtile_3__pin_outpad_0_
port 8 nsew signal input
rlabel metal3 s 0 4368 400 4424 6 ccff_head
port 9 nsew signal input
rlabel metal3 s 7600 4704 8000 4760 6 ccff_tail
port 10 nsew signal output
rlabel metal2 s 3360 0 3416 400 6 gfpga_pad_GPIO_PAD[0]
port 11 nsew signal bidirectional
rlabel metal3 s 0 3360 400 3416 6 gfpga_pad_GPIO_PAD[1]
port 12 nsew signal bidirectional
rlabel metal2 s 4032 0 4088 400 6 gfpga_pad_GPIO_PAD[2]
port 13 nsew signal bidirectional
rlabel metal3 s 7600 3360 8000 3416 6 gfpga_pad_GPIO_PAD[3]
port 14 nsew signal bidirectional
rlabel metal3 s 7600 4368 8000 4424 6 pReset
port 15 nsew signal input
rlabel metal3 s 0 4704 400 4760 6 prog_clk
port 16 nsew signal input
rlabel metal4 s 1418 1538 1578 6302 6 vdd
port 17 nsew power bidirectional
rlabel metal4 s 3070 1538 3230 6302 6 vdd
port 17 nsew power bidirectional
rlabel metal4 s 4722 1538 4882 6302 6 vdd
port 17 nsew power bidirectional
rlabel metal4 s 6374 1538 6534 6302 6 vdd
port 17 nsew power bidirectional
rlabel metal4 s 2244 1538 2404 6302 6 vss
port 18 nsew ground bidirectional
rlabel metal4 s 3896 1538 4056 6302 6 vss
port 18 nsew ground bidirectional
rlabel metal4 s 5548 1538 5708 6302 6 vss
port 18 nsew ground bidirectional
rlabel metal4 s 7200 1538 7360 6302 6 vss
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 8000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 163632
string GDS_FILE /home/baungarten/Desktop/2x2_FPGA_180nmD/openlane/grid_io_top/runs/23_12_09_13_11/results/signoff/grid_io_top.magic.gds
string GDS_START 74482
<< end >>

