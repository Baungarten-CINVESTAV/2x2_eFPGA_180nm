* NGSPICE file created from cby_1__1_.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

.subckt cby_1__1_ ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] left_grid_right_width_0_height_0_subtile_0__pin_I_1_
+ left_grid_right_width_0_height_0_subtile_0__pin_I_5_ pReset prog_clk right_grid_left_width_0_height_0_subtile_0__pin_I_3_
+ right_grid_left_width_0_height_0_subtile_0__pin_I_7_ vdd vss right_grid_left_width_0_height_0_subtile_0__pin_I_11_
+ left_grid_right_width_0_height_0_subtile_0__pin_I_9_
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__069__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_131_ net23 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_062_ _038_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input36_I chany_top_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_114_ net113 _034_ clknet_2_0__leaf_prog_clk mem_right_ipin_2.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_045_ _037_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold30 mem_right_ipin_0.DFFR_1_.Q net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput75 net75 chany_top_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput53 net53 chany_bottom_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput64 net64 chany_top_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input29_I chany_top_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_130_ net24 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_061_ _038_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_3_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_113_ net96 _033_ clknet_2_0__leaf_prog_clk mem_right_ipin_2.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_044_ _037_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_16_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold31 mem_right_ipin_0.DFFR_0_.Q net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold20 mem_right_ipin_0.DFFR_5_.Q net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_16_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I chany_bottom_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput76 net76 chany_top_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput65 net65 chany_top_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput54 net54 chany_bottom_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput43 net43 ccff_tail vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input3_I chany_bottom_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_060_ _038_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_10_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_043_ _037_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input41_I chany_top_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_112_ net115 _032_ clknet_2_0__leaf_prog_clk mem_right_ipin_2.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_8_Left_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold21 mem_left_ipin_2.DFFR_3_.Q net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 mem_left_ipin_1.DFFR_4_.Q net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold32 mem_right_ipin_1.DFFR_1_.Q net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput66 net66 chany_top_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput44 net44 chany_bottom_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput77 net77 chany_top_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput55 net55 chany_bottom_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I chany_top_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_111_ net92 _031_ clknet_2_2__leaf_prog_clk mem_right_ipin_2.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_042_ _037_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_21_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold11 mem_left_ipin_1.DFFR_5_.Q net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold22 mem_left_ipin_1.DFFR_2_.Q net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_15_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold33 mem_right_ipin_1.DFFR_4_.Q net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput78 net78 chany_top_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput56 net56 chany_bottom_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput45 net45 chany_bottom_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput67 net67 chany_top_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_11_Left_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__110__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input27_I chany_top_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_110_ net101 _030_ clknet_2_2__leaf_prog_clk net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_041_ _036_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_21_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold34 mem_left_ipin_0.DFFR_0_.Q net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold23 mem_left_ipin_0.DFFR_2_.Q net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold12 mem_right_ipin_2.DFFR_4_.Q net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xcby_1__1__84 left_grid_right_width_0_height_0_subtile_0__pin_I_9_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_2_3__f_prog_clk clknet_0_prog_clk clknet_2_3__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput57 net57 chany_bottom_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput46 net46 chany_bottom_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput79 net79 chany_top_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput68 net68 chany_top_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I ccff_head vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2__f_prog_clk clknet_0_prog_clk clknet_2_2__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_040_ net42 _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold35 mem_right_ipin_1.DFFR_5_.Q net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold13 mem_right_ipin_1.DFFR_2_.Q net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold24 mem_right_ipin_2.DFFR_0_.Q net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcby_1__1__85 left_grid_right_width_0_height_0_subtile_0__pin_I_5_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput58 net58 chany_bottom_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput69 net69 chany_top_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput47 net47 chany_bottom_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_1__f_prog_clk clknet_0_prog_clk clknet_2_1__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__098__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_28_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_099_ net104 _019_ clknet_2_3__leaf_prog_clk mem_right_ipin_0.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold14 mem_left_ipin_2.DFFR_4_.Q net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 mem_right_ipin_1.DFFR_0_.Q net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input32_I chany_top_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcby_1__1__86 left_grid_right_width_0_height_0_subtile_0__pin_I_1_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_6_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput59 net59 chany_bottom_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput48 net48 chany_bottom_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_0__f_prog_clk clknet_0_prog_clk clknet_2_0__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_098_ net94 _018_ clknet_2_2__leaf_prog_clk mem_right_ipin_0.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_3_Left_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold15 mem_right_ipin_0.DFFR_3_.Q net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input25_I chany_top_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold26 mem_right_ipin_2.DFFR_2_.Q net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcby_1__1__87 right_grid_left_width_0_height_0_subtile_0__pin_I_11_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_20_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput49 net49 chany_bottom_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_26_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_097_ net100 _017_ clknet_2_1__leaf_prog_clk mem_left_ipin_2.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold16 mem_left_ipin_2.DFFR_0_.Q net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold27 mem_right_ipin_0.DFFR_2_.Q net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input18_I chany_bottom_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcby_1__1__88 right_grid_left_width_0_height_0_subtile_0__pin_I_3_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_149_ net5 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_096_ net105 _016_ clknet_2_1__leaf_prog_clk mem_left_ipin_2.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold17 mem_left_ipin_2.DFFR_1_.Q net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 mem_left_ipin_0.DFFR_1_.Q net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_10_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_148_ net6 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcby_1__1__89 right_grid_left_width_0_height_0_subtile_0__pin_I_7_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_14_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_079_ _036_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input30_I chany_top_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_19_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__106__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_095_ net106 _015_ clknet_2_1__leaf_prog_clk mem_left_ipin_2.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold18 mem_left_ipin_1.DFFR_3_.Q net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold29 mem_right_ipin_1.DFFR_3_.Q net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_29_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Left_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_147_ net7 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_078_ _036_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input23_I chany_top_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__064__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_094_ net90 _014_ clknet_2_3__leaf_prog_clk mem_left_ipin_2.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_23_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold19 mem_left_ipin_0.DFFR_3_.Q net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__072__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_146_ net8 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__067__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_077_ _036_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input16_I chany_bottom_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I chany_bottom_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_129_ net25 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_10_Left_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_093_ net110 _013_ clknet_2_3__leaf_prog_clk mem_left_ipin_2.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_15_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_prog_clk prog_clk clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput1 ccff_head net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_29_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_145_ net9 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_076_ _036_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_059_ _038_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_128_ net26 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__109__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input39_I chany_top_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_161_ net2 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_092_ net103 _012_ clknet_2_3__leaf_prog_clk mem_left_ipin_2.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 chany_bottom_in[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_144_ net10 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_075_ _036_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_11_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_127_ net27 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_058_ _038_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input21_I chany_bottom_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_160_ net13 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_091_ net93 _011_ clknet_2_1__leaf_prog_clk mem_left_ipin_1.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 chany_bottom_in[10] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_143_ net11 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_074_ _036_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_27_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_126_ net28 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_057_ _038_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input14_I chany_bottom_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_22_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input6_I chany_bottom_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_109_ net109 _029_ clknet_2_2__leaf_prog_clk mem_right_ipin_1.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_12_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_090_ net91 _010_ clknet_2_3__leaf_prog_clk mem_left_ipin_1.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 chany_bottom_in[11] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_142_ net12 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_073_ _039_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_2_Left_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_125_ net29 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_056_ _038_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xinput40 chany_top_in[8] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_108_ net114 _028_ clknet_2_2__leaf_prog_clk mem_right_ipin_1.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_8_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 chany_bottom_in[12] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input37_I chany_top_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_141_ net22 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_072_ _039_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_055_ _038_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_124_ net30 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput41 chany_top_in[9] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput30 chany_top_in[17] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_107_ net121 _027_ clknet_2_2__leaf_prog_clk mem_right_ipin_1.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 chany_bottom_in[13] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_140_ net33 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_071_ _039_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_123_ net31 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 chany_top_in[18] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_054_ _038_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xinput20 chany_bottom_in[8] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 pReset net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_106_ net102 _026_ clknet_2_2__leaf_prog_clk mem_right_ipin_1.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input12_I chany_bottom_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I chany_bottom_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 chany_bottom_in[14] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_070_ _039_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Left_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input42_I pReset vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_053_ _038_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_122_ net32 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 chany_bottom_in[9] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 chany_top_in[19] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 chany_bottom_in[17] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_105_ net118 _025_ clknet_2_2__leaf_prog_clk mem_right_ipin_1.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 chany_bottom_in[15] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input35_I chany_top_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_22_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_052_ _036_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput11 chany_bottom_in[18] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 chany_top_in[0] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput33 chany_top_in[1] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_104_ net122 _024_ clknet_2_2__leaf_prog_clk mem_right_ipin_1.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 chany_bottom_in[16] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input28_I chany_top_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_051_ _037_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xinput34 chany_top_in[2] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 chany_top_in[10] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput12 chany_bottom_in[19] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_103_ net97 _023_ clknet_2_3__leaf_prog_clk mem_right_ipin_0.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold1 mem_left_ipin_2.DFFR_2_.Q net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input10_I chany_bottom_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I chany_bottom_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__105__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_050_ _037_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xinput13 chany_bottom_in[1] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 chany_top_in[3] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput24 chany_top_in[11] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_7_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input40_I chany_top_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_102_ net120 _022_ clknet_2_3__leaf_prog_clk mem_right_ipin_0.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_12_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold2 mem_left_ipin_1.DFFR_0_.Q net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_4_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput14 chany_bottom_in[2] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 chany_top_in[4] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 chany_top_in[12] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_7_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_101_ net119 _021_ clknet_2_3__leaf_prog_clk mem_right_ipin_0.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input33_I chany_top_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__070__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold3 mem_right_ipin_2.DFFR_3_.Q net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__065__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__073__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 chany_bottom_in[3] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput37 chany_top_in[5] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__068__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput26 chany_top_in[13] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_100_ net116 _020_ clknet_2_3__leaf_prog_clk mem_right_ipin_0.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input26_I chany_top_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__108__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold4 mem_left_ipin_0.DFFR_5_.Q net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_4_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_prog_clk_I prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput16 chany_bottom_in[4] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 chany_top_in[14] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput38 chany_top_in[6] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input19_I chany_bottom_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_159_ net14 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 mem_right_ipin_0.DFFR_4_.Q net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_28_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 chany_bottom_in[5] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 chany_top_in[15] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 chany_top_in[7] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_158_ net15 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_089_ net95 _009_ clknet_2_1__leaf_prog_clk mem_left_ipin_1.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input31_I chany_top_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold6 mem_left_ipin_1.DFFR_1_.Q net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_17_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 chany_top_in[16] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput18 chany_bottom_in[6] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Left_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_157_ net16 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_088_ net111 _008_ clknet_2_1__leaf_prog_clk mem_left_ipin_1.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_12_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input24_I chany_top_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold7 mem_right_ipin_2.DFFR_1_.Q net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 chany_bottom_in[7] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_156_ net17 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_087_ net107 _007_ clknet_2_1__leaf_prog_clk mem_left_ipin_1.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input17_I chany_bottom_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold8 mem_left_ipin_2.DFFR_5_.Q net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input9_I chany_bottom_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_139_ net34 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__111__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_086_ net99 _006_ clknet_2_1__leaf_prog_clk mem_left_ipin_1.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_12_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_155_ net18 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold9 mem_left_ipin_0.DFFR_4_.Q net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_138_ net35 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_069_ _039_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_154_ net19 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_085_ net1 _005_ clknet_2_0__leaf_prog_clk mem_left_ipin_0.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_9_Left_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_137_ net36 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_068_ _039_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input22_I chany_top_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput80 net80 chany_top_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_5_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_084_ net123 _004_ clknet_2_0__leaf_prog_clk mem_left_ipin_0.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_153_ net20 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_136_ net37 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_067_ _039_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_0_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I chany_bottom_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I chany_bottom_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 chany_top_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput81 net81 chany_top_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_152_ net21 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_0_Left_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_083_ net117 _003_ clknet_2_0__leaf_prog_clk mem_left_ipin_0.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_28_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_135_ net38 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_066_ _039_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_049_ _037_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_26_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__104__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput71 net71 chany_top_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput60 net60 chany_bottom_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_18_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput82 net82 chany_top_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_24_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input38_I chany_top_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_151_ net3 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_082_ net112 _002_ clknet_2_0__leaf_prog_clk mem_left_ipin_0.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_29_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_134_ net39 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_065_ _039_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_048_ _037_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input20_I chany_bottom_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput61 net61 chany_bottom_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_27_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput50 net50 chany_bottom_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput83 net83 chany_top_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput72 net72 chany_top_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_24_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_150_ net4 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_081_ net108 _001_ clknet_2_0__leaf_prog_clk mem_left_ipin_0.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_1_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_29_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_133_ net40 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_064_ _039_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_047_ _037_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input13_I chany_bottom_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I chany_bottom_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput51 net51 chany_bottom_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput73 net73 chany_top_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_27_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput62 net62 chany_bottom_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_24_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_080_ net98 _000_ clknet_2_0__leaf_prog_clk mem_left_ipin_0.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_29_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_132_ net41 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_4_Left_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_063_ _036_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_28_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__107__CLK clknet_2_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__071__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_046_ _037_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_115_ net124 _035_ clknet_2_0__leaf_prog_clk mem_right_ipin_2.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__066__I _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput52 net52 chany_bottom_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput74 net74 chany_top_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput63 net63 chany_bottom_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends

