* NGSPICE file created from sb_0__1_.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

.subckt sb_0__1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
+ bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
+ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
+ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[10]
+ chany_bottom_out[11] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[9] pReset prog_clk right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
+ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vdd vss chany_bottom_out[8]
+ chany_bottom_out[12] chany_bottom_out[16] chanx_right_out[10] chany_top_out[0] chanx_right_out[0]
+ chanx_right_out[11] chany_top_out[4] chany_top_out[8] chanx_right_out[1] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[2] chanx_right_out[14] chany_top_out[16] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[19] chany_bottom_out[0] chanx_right_out[5] chany_bottom_out[4]
+ chanx_right_out[6] chanx_right_out[7]
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_294_ net192 _058_ clknet_3_7__leaf_prog_clk net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__164__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__159__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_277_ net182 _041_ clknet_3_4__leaf_prog_clk mem_bottom_track_9.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input36_I pReset vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_200_ _115_ _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_10_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_131_ _107_ _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_4_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_329_ net114 _093_ clknet_3_3__leaf_prog_clk mem_right_track_6.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_10_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold52 mem_right_track_2.DFFR_3_.Q net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold63 mem_right_track_2.DFFR_2_.Q net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold30 mem_bottom_track_33.DFFR_0_.Q net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold85 mem_bottom_track_9.DFFR_3_.Q net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold74 mem_top_track_32.DFFR_1_.Q net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold41 mem_top_track_0.DFFR_2_.Q net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold96 mem_bottom_track_1.DFFR_2_.Q net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__247__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput42 net42 chany_bottom_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_3_7__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput64 net64 chany_top_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_18_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput53 net53 chany_bottom_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_15_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_293_ net115 _057_ clknet_3_7__leaf_prog_clk mem_bottom_track_25.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__180__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__308__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__175__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_276_ net102 _040_ clknet_3_5__leaf_prog_clk mem_bottom_track_17.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_130_ _108_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I chany_top_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_328_ net140 _092_ clknet_3_3__leaf_prog_clk mem_right_track_6.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__280__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_259_ net117 _023_ clknet_3_4__leaf_prog_clk mem_top_track_16.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold75 mem_right_track_10.DFFR_0_.D net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 mem_bottom_track_33.DFFR_3_.Q net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 mem_bottom_track_17.DFFR_3_.Q net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 mem_bottom_track_1.DFFR_6_.Q net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold64 mem_top_track_0.DFFR_5_.Q net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold31 mem_top_track_16.DFFR_4_.Q net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold97 mem_top_track_32.DFFR_3_.Q net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold20 mem_top_track_16.DFFR_3_.Q net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__183__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I chany_bottom_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput65 net65 chany_top_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput54 net54 chany_bottom_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__178__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput43 net43 chany_bottom_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_17_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I chany_bottom_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ net157 _056_ clknet_3_7__leaf_prog_clk mem_bottom_track_25.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_9_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__237__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_275_ net130 _039_ clknet_3_4__leaf_prog_clk mem_top_track_32.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__186__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_327_ net188 _091_ clknet_3_3__leaf_prog_clk mem_right_track_4.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_189_ _114_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_258_ net128 _022_ clknet_3_4__leaf_prog_clk mem_top_track_16.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_33_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__270__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold98 mem_bottom_track_25.DFFR_4_.Q net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold43 mem_right_track_6.DFFR_4_.Q net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold21 mem_bottom_track_33.DFFR_1_.Q net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 mem_right_track_8.DFFR_0_.Q net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold76 mem_bottom_track_17.DFFR_0_.D net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold32 mem_bottom_track_1.DFFR_0_.D net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold54 mem_bottom_track_1.DFFR_1_.Q net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 mem_top_track_16.DFFR_1_.Q net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 mem_top_track_24.DFFR_1_.Q net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__374__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput44 net44 chany_bottom_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput66 net66 chany_top_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput55 net55 chany_bottom_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_18_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_291_ net108 _055_ clknet_3_5__leaf_prog_clk mem_bottom_track_25.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_9_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__331__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_274_ net112 _038_ clknet_3_5__leaf_prog_clk mem_top_track_32.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_326_ net153 _090_ clknet_3_3__leaf_prog_clk mem_right_track_4.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_188_ _114_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_10_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_257_ net116 _021_ clknet_3_4__leaf_prog_clk mem_top_track_8.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_27_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input34_I chany_top_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__197__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_309_ net196 _073_ clknet_3_2__leaf_prog_clk mem_right_track_22.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold44 mem_right_track_2.DFFR_1_.Q net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 mem_right_track_0.DFFR_1_.Q net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 mem_right_track_6.DFFR_5_.Q net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold11 mem_bottom_track_25.DFFR_1_.Q net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold99 mem_right_track_20.DFFR_1_.Q net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 mem_top_track_24.DFFR_5_.Q net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold22 mem_top_track_0.DFFR_4_.Q net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 mem_top_track_8.DFFR_4_.Q net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 mem_top_track_16.DFFR_5_.Q net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_32_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput45 net45 chany_bottom_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput56 net56 chany_bottom_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput67 net67 chany_top_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__260__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_290_ net124 _054_ clknet_3_7__leaf_prog_clk mem_bottom_track_25.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__283__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_273_ net171 _037_ clknet_3_5__leaf_prog_clk mem_top_track_32.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_0_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_325_ net126 _089_ clknet_3_3__leaf_prog_clk mem_right_track_4.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_187_ _114_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_256_ net181 _020_ clknet_3_4__leaf_prog_clk mem_top_track_8.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input27_I chany_top_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_308_ net98 _072_ clknet_3_0__leaf_prog_clk mem_right_track_22.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_1_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_239_ net166 _003_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold56 mem_right_track_4.DFFR_0_.Q net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold78 mem_right_track_12.DFFR_1_.Q net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold12 mem_right_track_18.DFFR_0_.Q net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 mem_bottom_track_17.DFFR_4_.Q net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold89 mem_right_track_16.DFFR_1_.Q net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold45 mem_right_track_20.DFFR_0_.Q net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold67 mem_top_track_32.DFFR_4_.Q net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_7_Left_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold23 mem_top_track_16.DFFR_0_.Q net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_32_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput46 net46 chany_bottom_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput57 net57 chany_top_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput68 net68 chany_top_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I ccff_head vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ net186 _105_ clknet_3_3__leaf_prog_clk mem_right_track_18.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_20_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__250__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_272_ net187 _036_ clknet_3_5__leaf_prog_clk mem_top_track_32.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_20_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__273__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_324_ net178 _088_ clknet_3_3__leaf_prog_clk mem_right_track_4.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_186_ _106_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_255_ net189 _019_ clknet_3_1__leaf_prog_clk mem_top_track_8.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_27_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_307_ net191 _071_ clknet_3_2__leaf_prog_clk mem_right_track_20.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__311__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_169_ _112_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_238_ net119 _002_ clknet_3_1__leaf_prog_clk mem_top_track_0.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_30_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold79 mem_right_track_6.DFFR_1_.Q net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold57 mem_right_track_14.DFFR_0_.Q net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold35 mem_bottom_track_9.DFFR_2_.Q net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold13 mem_right_track_26.DFFR_0_.Q net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold24 mem_bottom_track_9.DFFR_1_.Q net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 mem_right_track_24.DFFR_0_.Q net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 mem_top_track_16.DFFR_0_.D net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__334__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput47 net47 chany_bottom_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput69 net69 chany_top_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput58 net58 chany_top_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_32_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_340_ net109 _104_ clknet_3_6__leaf_prog_clk mem_right_track_18.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_11_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_271_ net194 _035_ clknet_3_5__leaf_prog_clk mem_top_track_32.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__200__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_323_ net99 _087_ clknet_3_6__leaf_prog_clk mem_right_track_4.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_185_ _113_ _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_254_ net105 _018_ clknet_3_0__leaf_prog_clk mem_top_track_8.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__240__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_306_ net142 _070_ clknet_3_2__leaf_prog_clk mem_right_track_20.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_168_ _112_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_237_ net161 _001_ clknet_3_1__leaf_prog_clk mem_top_track_0.DFFR_6_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__263__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold14 mem_right_track_2.DFFR_4_.Q net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold36 mem_right_track_6.DFFR_2_.Q net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input32_I chany_top_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold47 mem_right_track_24.DFFR_1_.Q net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 mem_top_track_24.DFFR_4_.Q net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 mem_top_track_0.DFFR_3_.Q net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold58 mem_bottom_track_1.DFFR_0_.Q net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__286__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput48 net48 chany_bottom_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput59 net59 chany_top_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_26_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput37 net37 ccff_tail vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__203__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold100 mem_bottom_track_25.DFFR_3_.Q net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_270_ net164 _034_ clknet_3_5__leaf_prog_clk mem_right_track_0.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_399_ net13 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_322_ net113 _086_ clknet_3_7__leaf_prog_clk mem_right_track_4.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_184_ _113_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_27_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_253_ net145 _017_ clknet_3_0__leaf_prog_clk mem_top_track_8.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__241__RN _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_305_ net172 _069_ clknet_3_6__leaf_prog_clk mem_right_track_10.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_167_ _112_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_236_ net146 _000_ clknet_3_1__leaf_prog_clk mem_top_track_0.DFFR_7_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__121__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__206__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold59 mem_right_track_6.DFFR_0_.Q net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input25_I chany_top_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold37 mem_bottom_track_33.DFFR_2_.Q net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold26 mem_bottom_track_1.DFFR_5_.Q net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold15 mem_top_track_32.DFFR_0_.Q net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 mem_top_track_8.DFFR_3_.Q net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_32_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_219_ _106_ _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__253__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput38 net38 chanx_right_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput49 net49 chany_bottom_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_34_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__276__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__299__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold101 mem_top_track_0.DFFR_0_.Q net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__124__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_398_ net15 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__314__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_321_ net185 _085_ clknet_3_3__leaf_prog_clk mem_right_track_2.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_24_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__119__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_183_ _113_ _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__337__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_252_ net174 _016_ clknet_3_0__leaf_prog_clk mem_top_track_16.DFFR_0_.D vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_304_ net135 _068_ clknet_3_6__leaf_prog_clk mem_right_track_10.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_235_ _107_ _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_166_ _112_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold16 mem_right_track_4.DFFR_4_.Q net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold27 mem_bottom_track_25.DFFR_2_.Q net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold38 mem_right_track_10.DFFR_0_.Q net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__222__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I chany_bottom_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__132__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold49 mem_top_track_0.DFFR_6_.Q net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_218_ _116_ _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_27_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_149_ _110_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XTAP_TAPCELL_ROW_6_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput39 net39 chanx_right_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_11_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__127__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__230__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__243__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold102 mem_top_track_24.DFFR_3_.Q net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_24_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_397_ net16 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__140__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__266__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__225__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_320_ net100 _084_ clknet_3_6__leaf_prog_clk mem_right_track_2.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_182_ _113_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__135__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_251_ net129 _015_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__304__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_303_ net152 _067_ clknet_3_3__leaf_prog_clk mem_right_track_8.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_234_ _107_ _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_165_ _112_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold17 mem_right_track_6.DFFR_3_.Q net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_30_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold28 mem_right_track_22.DFFR_1_.Q net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold39 mem_bottom_track_1.DFFR_3_.Q net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_32_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_217_ _116_ _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_29_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_148_ _110_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XTAP_TAPCELL_ROW_6_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__233__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input30_I chany_top_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__143__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__228__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__138__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold103 mem_right_track_10.DFFR_1_.Q net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_396_ net17 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_181_ _113_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_250_ net155 _014_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__151__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_379_ net35 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_302_ net107 _066_ clknet_3_6__leaf_prog_clk mem_right_track_10.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_233_ _107_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_164_ _106_ _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__146__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold29 mem_right_track_4.DFFR_1_.Q net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_23_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold18 mem_bottom_track_17.DFFR_5_.Q net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_11_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_216_ _116_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_147_ _110_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input23_I chany_top_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__317__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__154__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold104 mem_bottom_track_25.DFFR_5_.Q net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__149__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_395_ net19 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_180_ _113_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_2_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_378_ net22 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_301_ net202 _065_ clknet_3_7__leaf_prog_clk mem_right_track_0.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_232_ _107_ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__162__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_163_ _111_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold19 mem_top_track_0.DFFR_7_.Q net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_215_ _116_ _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_146_ _110_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__157__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__246__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I chany_bottom_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_129_ _108_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XTAP_TAPCELL_ROW_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I chany_bottom_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold105 mem_right_track_0.DFFR_0_.D net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__307__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_394_ net20 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_377_ net23 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_300_ net159 _064_ clknet_3_7__leaf_prog_clk mem_right_track_0.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_231_ _107_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_24_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_162_ _111_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_3_Left_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_prog_clk prog_clk clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput1 ccff_head net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ _116_ _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_145_ _110_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_11_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__340__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_128_ _108_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_32_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__236__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__181__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_393_ net3 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__176__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_376_ net24 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_230_ _107_ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_161_ _111_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 chany_bottom_in[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_213_ _116_ _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_144_ _110_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__184__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_127_ _108_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input21_I chany_top_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__179__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__330__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_392_ net5 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_6__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output52_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_375_ net25 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__249__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_160_ _111_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_289_ net197 _053_ clknet_3_7__leaf_prog_clk mem_bottom_track_25.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 chany_bottom_in[10] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_212_ _116_ _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_143_ _110_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__380__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_126_ _108_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_33_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I chany_bottom_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__282__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I chany_bottom_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_391_ net6 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__320__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_374_ net26 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_288_ net195 _052_ clknet_3_7__leaf_prog_clk mem_bottom_track_25.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 chany_bottom_in[11] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_211_ _116_ _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_142_ _107_ _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_9_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__198__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__239__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_125_ _108_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_33_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_390_ net7 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_373_ net27 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__272__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 chany_bottom_in[12] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_287_ net173 _051_ clknet_3_5__leaf_prog_clk mem_bottom_track_17.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__310__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_210_ _116_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_141_ _109_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_9_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__333__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_339_ net103 _103_ clknet_3_3__leaf_prog_clk mem_right_track_16.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_124_ _108_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_26_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput30 chany_top_in[2] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_372_ net28 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output50_I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_286_ net167 _050_ clknet_3_5__leaf_prog_clk mem_bottom_track_17.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput6 chany_bottom_in[13] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__262__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_140_ _109_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_338_ net179 _102_ clknet_3_3__leaf_prog_clk mem_right_track_16.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_269_ net163 _033_ clknet_3_4__leaf_prog_clk mem_top_track_24.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_34_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput20 chany_bottom_in[9] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_123_ _108_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xinput31 chany_top_in[4] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__323__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_3__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I chany_bottom_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I chany_bottom_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ net8 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__201__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_285_ net190 _049_ clknet_3_3__leaf_prog_clk mem_bottom_track_17.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput7 chany_bottom_in[14] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_199_ _115_ _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_337_ net175 _101_ clknet_3_2__leaf_prog_clk mem_right_track_14.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_268_ net104 _032_ clknet_3_5__leaf_prog_clk mem_top_track_24.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_34_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_122_ _108_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__252__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput32 chany_top_in[5] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 chany_top_in[0] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 chany_bottom_in[17] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__298__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__204__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__313__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_370_ net4 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__336__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_284_ net101 _048_ clknet_3_6__leaf_prog_clk mem_bottom_track_17.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_17_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 chany_bottom_in[15] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_336_ net154 _100_ clknet_3_2__leaf_prog_clk mem_right_track_14.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_22_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_198_ _115_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__122__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_267_ net184 _031_ clknet_3_5__leaf_prog_clk mem_top_track_24.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_19_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__207__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I chany_top_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_121_ _108_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_319_ net141 _083_ clknet_3_6__leaf_prog_clk mem_right_track_2.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput33 chany_top_in[6] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 chany_bottom_in[18] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 chany_top_in[10] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_30_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__220__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__242__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__130__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__265__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__125__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_0__1__90 chanx_right_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_17_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_283_ net150 _047_ clknet_3_6__leaf_prog_clk mem_bottom_track_17.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput9 chany_bottom_in[16] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_335_ net200 _099_ clknet_3_2__leaf_prog_clk mem_right_track_12.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_197_ _106_ _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_266_ net147 _030_ clknet_3_5__leaf_prog_clk mem_top_track_24.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__223__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__133__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_120_ _107_ _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA_input28_I chany_top_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 chany_bottom_in[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_318_ net160 _082_ clknet_3_6__leaf_prog_clk mem_right_track_2.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 chany_top_in[8] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_249_ net151 _013_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 chany_top_in[12] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_30_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__128__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1 mem_right_track_22.DFFR_0_.Q net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__243__RN _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__231__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input10_I chany_bottom_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__141__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_0__1__80 chany_bottom_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__91 chanx_right_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input2_I chany_bottom_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__226__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_282_ net131 _046_ clknet_3_6__leaf_prog_clk mem_bottom_track_17.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__136__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__255__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_334_ net158 _098_ clknet_3_2__leaf_prog_clk mem_right_track_12.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_13_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_196_ _114_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_265_ net199 _029_ clknet_3_1__leaf_prog_clk mem_top_track_24.DFFR_4_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_33_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_317_ net149 _081_ clknet_3_6__leaf_prog_clk mem_right_track_2.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_179_ _113_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput24 chany_top_in[13] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 chany_top_in[9] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_248_ net193 _012_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput13 chany_bottom_in[2] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__234__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__144__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__229__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__139__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold2 mem_right_track_4.DFFR_3_.Q net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_20_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_0__1__92 chanx_right_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__81 chany_bottom_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_281_ net170 _045_ clknet_3_1__leaf_prog_clk mem_bottom_track_9.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__152__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ net180 _097_ clknet_3_2__leaf_prog_clk mem_right_track_6.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_28_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_195_ _114_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_264_ net122 _028_ clknet_3_4__leaf_prog_clk mem_top_track_24.DFFR_5_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__147__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 pReset net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_316_ net111 _080_ clknet_3_7__leaf_prog_clk mem_right_track_2.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput25 chany_top_in[14] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__245__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_247_ net136 _011_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput14 chany_bottom_in[3] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_178_ _113_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__268__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__160__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input33_I chany_top_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold3 mem_right_track_2.DFFR_0_.Q net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__155__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__306__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_0__1__82 chanx_right_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__93 chanx_right_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_280_ net177 _044_ clknet_3_1__leaf_prog_clk mem_bottom_track_9.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_332_ net156 _096_ clknet_3_2__leaf_prog_clk mem_right_track_6.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_401_ net2 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_194_ _114_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__163__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_263_ net143 _027_ clknet_3_0__leaf_prog_clk mem_top_track_16.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__158__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_177_ _113_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_315_ net168 _079_ clknet_3_3__leaf_prog_clk mem_right_track_28.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_246_ net148 _010_ clknet_3_0__leaf_prog_clk mem_bottom_track_1.DFFR_5_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput26 chany_top_in[16] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 chany_bottom_in[4] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input26_I chany_top_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_229_ _117_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk clknet_3_7__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 mem_bottom_track_17.DFFR_2_.Q net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_9_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_0__1__94 chanx_right_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__72 chany_top_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__83 chanx_right_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_clkbuf_0_prog_clk_I prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_400_ net12 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__319__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_331_ net176 _095_ clknet_3_2__leaf_prog_clk mem_right_track_6.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_193_ _114_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_22_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_262_ net120 _026_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_12_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__291__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput27 chany_top_in[17] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk clknet_3_6__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_24_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_176_ _113_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_314_ net106 _078_ clknet_3_1__leaf_prog_clk mem_bottom_track_1.DFFR_0_.D vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_245_ net123 _009_ clknet_3_1__leaf_prog_clk mem_bottom_track_1.DFFR_6_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput16 chany_bottom_in[5] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input19_I chany_bottom_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_228_ _117_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_25_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_159_ _111_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_8_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold5 mem_bottom_track_9.DFFR_4_.Q net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__182__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_0__1__95 chanx_right_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_15_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_0__1__84 chanx_right_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__73 chany_top_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__177__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__248__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_192_ _114_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_330_ net133 _094_ clknet_3_2__leaf_prog_clk mem_right_track_6.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk clknet_3_5__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_261_ net162 _025_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_175_ _106_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_313_ net144 _077_ clknet_3_2__leaf_prog_clk mem_right_track_26.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_244_ net139 _008_ clknet_3_1__leaf_prog_clk mem_bottom_track_1.DFFR_7_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput17 chany_bottom_in[6] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 chany_top_in[18] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__309__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_227_ _117_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__185__I _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_158_ _111_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__281__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input31_I chany_top_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold6 mem_right_track_14.DFFR_1_.Q net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_28_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_0__1__85 chanx_right_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_31_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_0__1__96 chanx_right_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__74 chany_top_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_output62_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk clknet_3_4__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_260_ net137 _024_ clknet_3_1__leaf_prog_clk mem_top_track_16.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_191_ _114_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_27_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_389_ net9 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__238__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_312_ net110 _076_ clknet_3_3__leaf_prog_clk mem_right_track_26.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput18 chany_bottom_in[7] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_174_ _112_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_243_ net1 _007_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_0_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput29 chany_top_in[1] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__381__I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_226_ _117_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_18_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_157_ _111_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input24_I chany_top_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold7 mem_top_track_24.DFFR_0_.Q net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_209_ _116_ _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk clknet_3_3__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_0__1__75 chany_top_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__86 chanx_right_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_3_5__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__271__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_0__1__97 chanx_right_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_190_ _114_ _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_388_ net10 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__332__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput19 chany_bottom_in[8] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_173_ _112_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_311_ net125 _075_ clknet_3_2__leaf_prog_clk mem_right_track_24.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_242_ net198 _006_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_1_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__199__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_225_ _117_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_18_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_156_ _111_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_34_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk clknet_3_2__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input17_I chany_bottom_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold8 mem_top_track_8.DFFR_2_.Q net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_208_ _106_ _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_139_ _109_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input9_I chany_bottom_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsb_0__1__76 chany_top_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsb_0__1__87 chanx_right_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_22_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__261__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_387_ net11 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__395__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__284__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_310_ net165 _074_ clknet_3_2__leaf_prog_clk mem_right_track_24.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_1_Left_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_172_ _112_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_15_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk clknet_3_1__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_241_ net169 _005_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_2_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_224_ _117_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_14_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_155_ _111_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_34_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 mem_right_track_28.DFFR_0_.Q net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_207_ _115_ _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_138_ _109_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xsb_0__1__88 chanx_right_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsb_0__1__77 chany_bottom_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_5_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_386_ net21 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk clknet_3_0__leaf_prog_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_171_ _112_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_240_ net138 _004_ clknet_3_0__leaf_prog_clk mem_top_track_0.DFFR_3_.Q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ net18 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__251__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_223_ _117_ _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_154_ _111_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__274__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_206_ _115_ _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_137_ _109_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_9_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input22_I chany_top_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsb_0__1__89 chanx_right_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_0_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsb_0__1__78 chany_bottom_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__335__CLK clknet_3_2__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold90 mem_top_track_32.DFFR_2_.Q net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__202__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_385_ net29 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_170_ _112_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_299_ net201 _063_ clknet_3_6__leaf_prog_clk mem_bottom_track_33.DFFR_0_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_368_ net14 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_222_ _117_ _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_153_ _107_ _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_11_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_205_ _115_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_136_ _109_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__241__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__120__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__205__I _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2__f_prog_clk_I clknet_0_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input15_I chany_bottom_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xsb_0__1__79 chany_bottom_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_119_ _106_ _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_15_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I chany_bottom_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__287__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold91 mem_right_track_2.DFFR_5_.Q net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold80 mem_bottom_track_9.DFFR_0_.Q net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__302__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_384_ net30 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput70 net70 chany_top_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__123__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_298_ net127 _062_ clknet_3_6__leaf_prog_clk mem_bottom_track_33.DFFR_1_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__208__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_221_ _117_ _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_12_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_152_ _110_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_11_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_204_ _115_ _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_6_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_135_ _109_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__221__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_118_ net36 _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__131__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_8_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold81 mem_right_track_4.DFFR_2_.Q net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_34_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold70 mem_bottom_track_17.DFFR_0_.Q net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__126__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold92 mem_top_track_8.DFFR_1_.Q net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__254__CLK clknet_3_0__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_383_ net31 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput71 net71 chany_top_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput60 net60 chany_top_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_297_ net118 _061_ clknet_3_7__leaf_prog_clk mem_bottom_track_33.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_21_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__224__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_220_ _117_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__134__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_151_ _110_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_34_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__219__I _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__129__I _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_203_ _115_ _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_134_ _109_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__232__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__142__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input20_I chany_bottom_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold82 mem_right_track_16.DFFR_0_.Q net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold93 mem_bottom_track_17.DFFR_1_.Q net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold71 mem_right_track_26.DFFR_1_.Q net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold60 mem_bottom_track_25.DFFR_0_.Q net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__227__I _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput50 net50 chany_bottom_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__137__I _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_382_ net32 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput61 net61 chany_top_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_24_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_296_ net134 _060_ clknet_3_7__leaf_prog_clk mem_bottom_track_33.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__244__CLK clknet_3_1__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__267__CLK clknet_3_5__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_150_ _110_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_279_ net121 _043_ clknet_3_4__leaf_prog_clk mem_bottom_track_9.DFFR_2_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__150__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__235__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_133_ _109_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_202_ _115_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__145__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__305__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I chany_bottom_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold83 mem_right_track_4.DFFR_5_.Q net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold61 mem_right_track_12.DFFR_0_.Q net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold94 mem_right_track_18.DFFR_1_.Q net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_21_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold72 mem_top_track_0.DFFR_1_.Q net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold50 mem_top_track_24.DFFR_2_.Q net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_6_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input5_I chany_bottom_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput40 net40 chanx_right_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput62 net62 chany_top_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_381_ net33 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__153__I _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput51 net51 chany_bottom_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__148__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_295_ net183 _059_ clknet_3_7__leaf_prog_clk mem_bottom_track_33.DFFR_4_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_23_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_278_ net132 _042_ clknet_3_4__leaf_prog_clk mem_bottom_track_9.DFFR_3_.Q vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_34_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_201_ _115_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_132_ _109_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__161__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__156__I _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold95 mem_bottom_track_33.DFFR_4_.Q net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 mem_right_track_0.DFFR_0_.Q net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold51 mem_bottom_track_1.DFFR_4_.Q net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold73 mem_bottom_track_1.DFFR_7_.Q net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold84 mem_top_track_8.DFFR_0_.Q net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold40 mem_top_track_16.DFFR_2_.Q net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_32_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput52 net52 chany_bottom_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_380_ net34 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput41 net41 chanx_right_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__318__CLK clknet_3_6__leaf_prog_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput63 net63 chany_top_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends

