magic
tech gf180mcuD
magscale 1 10
timestamp 1702149233
<< metal1 >>
rect 29250 30718 29262 30770
rect 29314 30767 29326 30770
rect 30146 30767 30158 30770
rect 29314 30721 30158 30767
rect 29314 30718 29326 30721
rect 30146 30718 30158 30721
rect 30210 30718 30222 30770
rect 1344 30602 32592 30636
rect 1344 30550 5120 30602
rect 5172 30550 5224 30602
rect 5276 30550 5328 30602
rect 5380 30550 12932 30602
rect 12984 30550 13036 30602
rect 13088 30550 13140 30602
rect 13192 30550 20744 30602
rect 20796 30550 20848 30602
rect 20900 30550 20952 30602
rect 21004 30550 28556 30602
rect 28608 30550 28660 30602
rect 28712 30550 28764 30602
rect 28816 30550 32592 30602
rect 1344 30516 32592 30550
rect 7410 30270 7422 30322
rect 7474 30270 7486 30322
rect 11554 30270 11566 30322
rect 11618 30270 11630 30322
rect 14914 30270 14926 30322
rect 14978 30270 14990 30322
rect 17938 30270 17950 30322
rect 18002 30270 18014 30322
rect 21746 30270 21758 30322
rect 21810 30270 21822 30322
rect 30146 30270 30158 30322
rect 30210 30270 30222 30322
rect 2158 30210 2210 30222
rect 2158 30146 2210 30158
rect 13582 30210 13634 30222
rect 13582 30146 13634 30158
rect 14030 30210 14082 30222
rect 21422 30210 21474 30222
rect 19954 30158 19966 30210
rect 20018 30158 20030 30210
rect 25218 30158 25230 30210
rect 25282 30158 25294 30210
rect 26898 30158 26910 30210
rect 26962 30158 26974 30210
rect 14030 30146 14082 30158
rect 21422 30146 21474 30158
rect 3390 30098 3442 30110
rect 3390 30034 3442 30046
rect 4958 30098 5010 30110
rect 4958 30034 5010 30046
rect 5630 30098 5682 30110
rect 9438 30098 9490 30110
rect 5954 30046 5966 30098
rect 6018 30046 6030 30098
rect 8642 30046 8654 30098
rect 8706 30046 8718 30098
rect 5630 30034 5682 30046
rect 9438 30034 9490 30046
rect 9774 30098 9826 30110
rect 12014 30098 12066 30110
rect 10546 30046 10558 30098
rect 10610 30046 10622 30098
rect 9774 30034 9826 30046
rect 12014 30034 12066 30046
rect 13246 30098 13298 30110
rect 23886 30098 23938 30110
rect 16258 30046 16270 30098
rect 16322 30046 16334 30098
rect 19170 30046 19182 30098
rect 19234 30046 19246 30098
rect 22754 30046 22766 30098
rect 22818 30046 22830 30098
rect 23538 30046 23550 30098
rect 23602 30046 23614 30098
rect 13246 30034 13298 30046
rect 23886 30034 23938 30046
rect 24782 30098 24834 30110
rect 27358 30098 27410 30110
rect 26674 30046 26686 30098
rect 26738 30046 26750 30098
rect 24782 30034 24834 30046
rect 27358 30034 27410 30046
rect 28478 30098 28530 30110
rect 28802 30046 28814 30098
rect 28866 30046 28878 30098
rect 31266 30046 31278 30098
rect 31330 30046 31342 30098
rect 28478 30034 28530 30046
rect 1934 29986 1986 29998
rect 1934 29922 1986 29934
rect 2942 29986 2994 29998
rect 2942 29922 2994 29934
rect 3838 29986 3890 29998
rect 3838 29922 3890 29934
rect 4174 29986 4226 29998
rect 4174 29922 4226 29934
rect 6414 29986 6466 29998
rect 6414 29922 6466 29934
rect 6974 29986 7026 29998
rect 6974 29922 7026 29934
rect 19742 29986 19794 29998
rect 19742 29922 19794 29934
rect 21086 29986 21138 29998
rect 21086 29922 21138 29934
rect 25902 29986 25954 29998
rect 25902 29922 25954 29934
rect 27470 29986 27522 29998
rect 27470 29922 27522 29934
rect 1344 29818 32752 29852
rect 1344 29766 9026 29818
rect 9078 29766 9130 29818
rect 9182 29766 9234 29818
rect 9286 29766 16838 29818
rect 16890 29766 16942 29818
rect 16994 29766 17046 29818
rect 17098 29766 24650 29818
rect 24702 29766 24754 29818
rect 24806 29766 24858 29818
rect 24910 29766 32462 29818
rect 32514 29766 32566 29818
rect 32618 29766 32670 29818
rect 32722 29766 32752 29818
rect 1344 29732 32752 29766
rect 1822 29650 1874 29662
rect 1822 29586 1874 29598
rect 9550 29650 9602 29662
rect 9550 29586 9602 29598
rect 10782 29650 10834 29662
rect 10782 29586 10834 29598
rect 19070 29650 19122 29662
rect 19070 29586 19122 29598
rect 19406 29650 19458 29662
rect 23998 29650 24050 29662
rect 20178 29598 20190 29650
rect 20242 29598 20254 29650
rect 19406 29586 19458 29598
rect 23998 29586 24050 29598
rect 28142 29650 28194 29662
rect 28142 29586 28194 29598
rect 5182 29538 5234 29550
rect 8978 29486 8990 29538
rect 9042 29486 9054 29538
rect 12002 29486 12014 29538
rect 12066 29486 12078 29538
rect 16594 29486 16606 29538
rect 16658 29486 16670 29538
rect 27234 29486 27246 29538
rect 27298 29486 27310 29538
rect 30258 29486 30270 29538
rect 30322 29486 30334 29538
rect 5182 29474 5234 29486
rect 2606 29426 2658 29438
rect 2606 29362 2658 29374
rect 2942 29426 2994 29438
rect 8094 29426 8146 29438
rect 23102 29426 23154 29438
rect 25342 29426 25394 29438
rect 7410 29374 7422 29426
rect 7474 29374 7486 29426
rect 8754 29374 8766 29426
rect 8818 29374 8830 29426
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 17490 29374 17502 29426
rect 17554 29374 17566 29426
rect 22530 29374 22542 29426
rect 22594 29374 22606 29426
rect 24322 29374 24334 29426
rect 24386 29374 24398 29426
rect 2942 29362 2994 29374
rect 8094 29362 8146 29374
rect 23102 29362 23154 29374
rect 25342 29362 25394 29374
rect 30942 29426 30994 29438
rect 30942 29362 30994 29374
rect 4174 29314 4226 29326
rect 3602 29262 3614 29314
rect 3666 29262 3678 29314
rect 4174 29250 4226 29262
rect 11342 29314 11394 29326
rect 32174 29314 32226 29326
rect 13010 29262 13022 29314
rect 13074 29262 13086 29314
rect 15362 29262 15374 29314
rect 15426 29262 15438 29314
rect 17826 29262 17838 29314
rect 17890 29262 17902 29314
rect 26226 29262 26238 29314
rect 26290 29262 26302 29314
rect 29026 29262 29038 29314
rect 29090 29262 29102 29314
rect 11342 29250 11394 29262
rect 32174 29250 32226 29262
rect 4398 29202 4450 29214
rect 4398 29138 4450 29150
rect 31726 29202 31778 29214
rect 31726 29138 31778 29150
rect 1344 29034 32592 29068
rect 1344 28982 5120 29034
rect 5172 28982 5224 29034
rect 5276 28982 5328 29034
rect 5380 28982 12932 29034
rect 12984 28982 13036 29034
rect 13088 28982 13140 29034
rect 13192 28982 20744 29034
rect 20796 28982 20848 29034
rect 20900 28982 20952 29034
rect 21004 28982 28556 29034
rect 28608 28982 28660 29034
rect 28712 28982 28764 29034
rect 28816 28982 32592 29034
rect 1344 28948 32592 28982
rect 17054 28866 17106 28878
rect 9314 28814 9326 28866
rect 9378 28863 9390 28866
rect 9986 28863 9998 28866
rect 9378 28817 9998 28863
rect 9378 28814 9390 28817
rect 9986 28814 9998 28817
rect 10050 28814 10062 28866
rect 17054 28802 17106 28814
rect 20862 28866 20914 28878
rect 20862 28802 20914 28814
rect 9550 28754 9602 28766
rect 4050 28702 4062 28754
rect 4114 28702 4126 28754
rect 6850 28702 6862 28754
rect 6914 28702 6926 28754
rect 9090 28702 9102 28754
rect 9154 28702 9166 28754
rect 9550 28690 9602 28702
rect 10110 28754 10162 28766
rect 11666 28702 11678 28754
rect 11730 28702 11742 28754
rect 21858 28702 21870 28754
rect 21922 28702 21934 28754
rect 27570 28702 27582 28754
rect 27634 28702 27646 28754
rect 30146 28702 30158 28754
rect 30210 28702 30222 28754
rect 10110 28690 10162 28702
rect 6190 28642 6242 28654
rect 2034 28590 2046 28642
rect 2098 28590 2110 28642
rect 6190 28578 6242 28590
rect 7310 28642 7362 28654
rect 22542 28642 22594 28654
rect 26238 28642 26290 28654
rect 13458 28590 13470 28642
rect 13522 28590 13534 28642
rect 13906 28590 13918 28642
rect 13970 28590 13982 28642
rect 17266 28590 17278 28642
rect 17330 28590 17342 28642
rect 17714 28590 17726 28642
rect 17778 28590 17790 28642
rect 25890 28590 25902 28642
rect 25954 28590 25966 28642
rect 7310 28578 7362 28590
rect 22542 28578 22594 28590
rect 26238 28578 26290 28590
rect 2270 28530 2322 28542
rect 5742 28530 5794 28542
rect 21310 28530 21362 28542
rect 3042 28478 3054 28530
rect 3106 28478 3118 28530
rect 7746 28478 7758 28530
rect 7810 28478 7822 28530
rect 12786 28478 12798 28530
rect 12850 28478 12862 28530
rect 2270 28466 2322 28478
rect 5742 28466 5794 28478
rect 21310 28466 21362 28478
rect 23550 28530 23602 28542
rect 23550 28466 23602 28478
rect 26798 28530 26850 28542
rect 31950 28530 32002 28542
rect 31154 28478 31166 28530
rect 31218 28478 31230 28530
rect 26798 28466 26850 28478
rect 31950 28466 32002 28478
rect 22766 28418 22818 28430
rect 16482 28366 16494 28418
rect 16546 28366 16558 28418
rect 20066 28366 20078 28418
rect 20130 28366 20142 28418
rect 22766 28354 22818 28366
rect 27134 28418 27186 28430
rect 27134 28354 27186 28366
rect 1344 28250 32752 28284
rect 1344 28198 9026 28250
rect 9078 28198 9130 28250
rect 9182 28198 9234 28250
rect 9286 28198 16838 28250
rect 16890 28198 16942 28250
rect 16994 28198 17046 28250
rect 17098 28198 24650 28250
rect 24702 28198 24754 28250
rect 24806 28198 24858 28250
rect 24910 28198 32462 28250
rect 32514 28198 32566 28250
rect 32618 28198 32670 28250
rect 32722 28198 32752 28250
rect 1344 28164 32752 28198
rect 8990 28082 9042 28094
rect 16942 28082 16994 28094
rect 12562 28030 12574 28082
rect 12626 28030 12638 28082
rect 16370 28030 16382 28082
rect 16434 28030 16446 28082
rect 23314 28030 23326 28082
rect 23378 28030 23390 28082
rect 31490 28030 31502 28082
rect 31554 28030 31566 28082
rect 8990 28018 9042 28030
rect 16942 28018 16994 28030
rect 5182 27970 5234 27982
rect 2146 27918 2158 27970
rect 2210 27918 2222 27970
rect 5182 27906 5234 27918
rect 8654 27970 8706 27982
rect 24110 27970 24162 27982
rect 20066 27918 20078 27970
rect 20130 27918 20142 27970
rect 24322 27918 24334 27970
rect 24386 27918 24398 27970
rect 27234 27918 27246 27970
rect 27298 27918 27310 27970
rect 8654 27906 8706 27918
rect 24110 27906 24162 27918
rect 8094 27858 8146 27870
rect 7410 27806 7422 27858
rect 7474 27806 7486 27858
rect 8094 27794 8146 27806
rect 9662 27858 9714 27870
rect 20638 27858 20690 27870
rect 28590 27858 28642 27870
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 13346 27806 13358 27858
rect 13410 27806 13422 27858
rect 13794 27806 13806 27858
rect 13858 27806 13870 27858
rect 21074 27806 21086 27858
rect 21138 27806 21150 27858
rect 24546 27806 24558 27858
rect 24610 27806 24622 27858
rect 29250 27806 29262 27858
rect 29314 27806 29326 27858
rect 9662 27794 9714 27806
rect 20638 27794 20690 27806
rect 28590 27794 28642 27806
rect 25342 27746 25394 27758
rect 28030 27746 28082 27758
rect 3154 27694 3166 27746
rect 3218 27694 3230 27746
rect 18722 27694 18734 27746
rect 18786 27694 18798 27746
rect 26226 27694 26238 27746
rect 26290 27694 26302 27746
rect 28354 27694 28366 27746
rect 28418 27694 28430 27746
rect 25342 27682 25394 27694
rect 28030 27682 28082 27694
rect 4398 27634 4450 27646
rect 4398 27570 4450 27582
rect 13134 27634 13186 27646
rect 13134 27570 13186 27582
rect 32286 27634 32338 27646
rect 32286 27570 32338 27582
rect 1344 27466 32592 27500
rect 1344 27414 5120 27466
rect 5172 27414 5224 27466
rect 5276 27414 5328 27466
rect 5380 27414 12932 27466
rect 12984 27414 13036 27466
rect 13088 27414 13140 27466
rect 13192 27414 20744 27466
rect 20796 27414 20848 27466
rect 20900 27414 20952 27466
rect 21004 27414 28556 27466
rect 28608 27414 28660 27466
rect 28712 27414 28764 27466
rect 28816 27414 32592 27466
rect 1344 27380 32592 27414
rect 8766 27298 8818 27310
rect 8766 27234 8818 27246
rect 19742 27298 19794 27310
rect 19742 27234 19794 27246
rect 22206 27298 22258 27310
rect 22206 27234 22258 27246
rect 4510 27186 4562 27198
rect 7982 27186 8034 27198
rect 20750 27186 20802 27198
rect 4050 27134 4062 27186
rect 4114 27134 4126 27186
rect 7522 27134 7534 27186
rect 7586 27134 7598 27186
rect 13682 27134 13694 27186
rect 13746 27134 13758 27186
rect 14802 27134 14814 27186
rect 14866 27134 14878 27186
rect 19954 27134 19966 27186
rect 20018 27134 20030 27186
rect 4510 27122 4562 27134
rect 7982 27122 8034 27134
rect 20750 27122 20802 27134
rect 21646 27186 21698 27198
rect 27570 27134 27582 27186
rect 27634 27134 27646 27186
rect 30706 27134 30718 27186
rect 30770 27134 30782 27186
rect 21646 27122 21698 27134
rect 12462 27074 12514 27086
rect 2034 27022 2046 27074
rect 2098 27022 2110 27074
rect 11890 27022 11902 27074
rect 11954 27022 11966 27074
rect 12462 27010 12514 27022
rect 15598 27074 15650 27086
rect 15598 27010 15650 27022
rect 16270 27074 16322 27086
rect 25678 27074 25730 27086
rect 16594 27022 16606 27074
rect 16658 27022 16670 27074
rect 25218 27022 25230 27074
rect 25282 27022 25294 27074
rect 16270 27010 16322 27022
rect 25678 27010 25730 27022
rect 2270 26962 2322 26974
rect 9550 26962 9602 26974
rect 3042 26910 3054 26962
rect 3106 26910 3118 26962
rect 6514 26910 6526 26962
rect 6578 26910 6590 26962
rect 2270 26898 2322 26910
rect 9550 26898 9602 26910
rect 14030 26962 14082 26974
rect 14030 26898 14082 26910
rect 14366 26962 14418 26974
rect 14366 26898 14418 26910
rect 20302 26962 20354 26974
rect 22990 26962 23042 26974
rect 21298 26910 21310 26962
rect 21362 26910 21374 26962
rect 26562 26910 26574 26962
rect 26626 26910 26638 26962
rect 31938 26910 31950 26962
rect 32002 26910 32014 26962
rect 20302 26898 20354 26910
rect 22990 26898 23042 26910
rect 5742 26850 5794 26862
rect 5742 26786 5794 26798
rect 8542 26850 8594 26862
rect 8542 26786 8594 26798
rect 12686 26850 12738 26862
rect 29374 26850 29426 26862
rect 18946 26798 18958 26850
rect 19010 26798 19022 26850
rect 12686 26786 12738 26798
rect 29374 26786 29426 26798
rect 1344 26682 32752 26716
rect 1344 26630 9026 26682
rect 9078 26630 9130 26682
rect 9182 26630 9234 26682
rect 9286 26630 16838 26682
rect 16890 26630 16942 26682
rect 16994 26630 17046 26682
rect 17098 26630 24650 26682
rect 24702 26630 24754 26682
rect 24806 26630 24858 26682
rect 24910 26630 32462 26682
rect 32514 26630 32566 26682
rect 32618 26630 32670 26682
rect 32722 26630 32752 26682
rect 1344 26596 32752 26630
rect 10222 26514 10274 26526
rect 16942 26514 16994 26526
rect 24110 26514 24162 26526
rect 16370 26462 16382 26514
rect 16434 26462 16446 26514
rect 21298 26462 21310 26514
rect 21362 26462 21374 26514
rect 10222 26450 10274 26462
rect 16942 26450 16994 26462
rect 24110 26450 24162 26462
rect 24558 26514 24610 26526
rect 32174 26514 32226 26526
rect 31266 26462 31278 26514
rect 31330 26462 31342 26514
rect 24558 26450 24610 26462
rect 32174 26450 32226 26462
rect 2382 26402 2434 26414
rect 8318 26402 8370 26414
rect 3154 26350 3166 26402
rect 3218 26350 3230 26402
rect 2382 26338 2434 26350
rect 8318 26338 8370 26350
rect 9102 26402 9154 26414
rect 9102 26338 9154 26350
rect 9886 26402 9938 26414
rect 21982 26402 22034 26414
rect 10994 26350 11006 26402
rect 11058 26350 11070 26402
rect 17378 26350 17390 26402
rect 17442 26350 17454 26402
rect 22306 26350 22318 26402
rect 22370 26350 22382 26402
rect 27234 26350 27246 26402
rect 27298 26350 27310 26402
rect 9886 26338 9938 26350
rect 21982 26338 22034 26350
rect 5630 26290 5682 26302
rect 13022 26290 13074 26302
rect 18286 26290 18338 26302
rect 28366 26290 28418 26302
rect 2146 26238 2158 26290
rect 2210 26238 2222 26290
rect 5954 26238 5966 26290
rect 6018 26238 6030 26290
rect 13346 26238 13358 26290
rect 13410 26238 13422 26290
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 18834 26238 18846 26290
rect 18898 26238 18910 26290
rect 28802 26238 28814 26290
rect 28866 26238 28878 26290
rect 5630 26226 5682 26238
rect 13022 26226 13074 26238
rect 18286 26226 18338 26238
rect 28366 26226 28418 26238
rect 4734 26178 4786 26190
rect 4162 26126 4174 26178
rect 4226 26126 4238 26178
rect 4734 26114 4786 26126
rect 5070 26178 5122 26190
rect 12462 26178 12514 26190
rect 11890 26126 11902 26178
rect 11954 26126 11966 26178
rect 5070 26114 5122 26126
rect 12462 26114 12514 26126
rect 17726 26178 17778 26190
rect 25454 26178 25506 26190
rect 23426 26126 23438 26178
rect 23490 26126 23502 26178
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 17726 26114 17778 26126
rect 25454 26114 25506 26126
rect 31838 26066 31890 26078
rect 31838 26002 31890 26014
rect 1344 25898 32592 25932
rect 1344 25846 5120 25898
rect 5172 25846 5224 25898
rect 5276 25846 5328 25898
rect 5380 25846 12932 25898
rect 12984 25846 13036 25898
rect 13088 25846 13140 25898
rect 13192 25846 20744 25898
rect 20796 25846 20848 25898
rect 20900 25846 20952 25898
rect 21004 25846 28556 25898
rect 28608 25846 28660 25898
rect 28712 25846 28764 25898
rect 28816 25846 32592 25898
rect 1344 25812 32592 25846
rect 6078 25730 6130 25742
rect 6078 25666 6130 25678
rect 14590 25730 14642 25742
rect 24894 25730 24946 25742
rect 22642 25727 22654 25730
rect 14590 25666 14642 25678
rect 22097 25681 22654 25727
rect 4734 25618 4786 25630
rect 1922 25566 1934 25618
rect 1986 25566 1998 25618
rect 3826 25566 3838 25618
rect 3890 25566 3902 25618
rect 4734 25554 4786 25566
rect 8094 25618 8146 25630
rect 22097 25618 22143 25681
rect 22642 25678 22654 25681
rect 22706 25678 22718 25730
rect 24894 25666 24946 25678
rect 22654 25618 22706 25630
rect 12562 25566 12574 25618
rect 12626 25566 12638 25618
rect 16482 25566 16494 25618
rect 16546 25566 16558 25618
rect 19282 25566 19294 25618
rect 19346 25566 19358 25618
rect 21746 25566 21758 25618
rect 21810 25566 21822 25618
rect 22082 25566 22094 25618
rect 22146 25566 22158 25618
rect 24322 25566 24334 25618
rect 24386 25566 24398 25618
rect 30146 25566 30158 25618
rect 30210 25566 30222 25618
rect 8094 25554 8146 25566
rect 22654 25554 22706 25566
rect 11790 25506 11842 25518
rect 15262 25506 15314 25518
rect 28366 25506 28418 25518
rect 2930 25454 2942 25506
rect 2994 25454 3006 25506
rect 3378 25454 3390 25506
rect 3442 25454 3454 25506
rect 11106 25454 11118 25506
rect 11170 25454 11182 25506
rect 13794 25454 13806 25506
rect 13858 25454 13870 25506
rect 21522 25454 21534 25506
rect 21586 25454 21598 25506
rect 27906 25454 27918 25506
rect 27970 25454 27982 25506
rect 11790 25442 11842 25454
rect 15262 25442 15314 25454
rect 28366 25442 28418 25454
rect 4958 25394 5010 25406
rect 7758 25394 7810 25406
rect 7410 25342 7422 25394
rect 7474 25342 7486 25394
rect 4958 25330 5010 25342
rect 7758 25330 7810 25342
rect 12014 25394 12066 25406
rect 12014 25330 12066 25342
rect 12798 25394 12850 25406
rect 25678 25394 25730 25406
rect 32174 25394 32226 25406
rect 17490 25342 17502 25394
rect 17554 25342 17566 25394
rect 20290 25342 20302 25394
rect 20354 25342 20366 25394
rect 23202 25342 23214 25394
rect 23266 25342 23278 25394
rect 31490 25342 31502 25394
rect 31554 25342 31566 25394
rect 12798 25330 12850 25342
rect 25678 25330 25730 25342
rect 32174 25330 32226 25342
rect 5742 25282 5794 25294
rect 5742 25218 5794 25230
rect 6862 25282 6914 25294
rect 22206 25282 22258 25294
rect 8866 25230 8878 25282
rect 8930 25230 8942 25282
rect 6862 25218 6914 25230
rect 22206 25218 22258 25230
rect 1344 25114 32752 25148
rect 1344 25062 9026 25114
rect 9078 25062 9130 25114
rect 9182 25062 9234 25114
rect 9286 25062 16838 25114
rect 16890 25062 16942 25114
rect 16994 25062 17046 25114
rect 17098 25062 24650 25114
rect 24702 25062 24754 25114
rect 24806 25062 24858 25114
rect 24910 25062 32462 25114
rect 32514 25062 32566 25114
rect 32618 25062 32670 25114
rect 32722 25062 32752 25114
rect 1344 25028 32752 25062
rect 3726 24946 3778 24958
rect 3726 24882 3778 24894
rect 8094 24946 8146 24958
rect 8094 24882 8146 24894
rect 8878 24946 8930 24958
rect 8878 24882 8930 24894
rect 10782 24946 10834 24958
rect 15486 24946 15538 24958
rect 14690 24894 14702 24946
rect 14754 24894 14766 24946
rect 10782 24882 10834 24894
rect 15486 24882 15538 24894
rect 16830 24946 16882 24958
rect 16830 24882 16882 24894
rect 18958 24946 19010 24958
rect 18958 24882 19010 24894
rect 19742 24946 19794 24958
rect 19742 24882 19794 24894
rect 24446 24946 24498 24958
rect 32286 24946 32338 24958
rect 31714 24894 31726 24946
rect 31778 24894 31790 24946
rect 24446 24882 24498 24894
rect 32286 24882 32338 24894
rect 4958 24834 5010 24846
rect 4958 24770 5010 24782
rect 15262 24834 15314 24846
rect 20526 24834 20578 24846
rect 23998 24834 24050 24846
rect 18050 24782 18062 24834
rect 18114 24782 18126 24834
rect 23650 24782 23662 24834
rect 23714 24782 23726 24834
rect 15262 24770 15314 24782
rect 20526 24770 20578 24782
rect 23998 24770 24050 24782
rect 24334 24834 24386 24846
rect 27234 24782 27246 24834
rect 27298 24782 27310 24834
rect 24334 24770 24386 24782
rect 2942 24722 2994 24734
rect 8990 24722 9042 24734
rect 11566 24722 11618 24734
rect 18398 24722 18450 24734
rect 23214 24722 23266 24734
rect 3714 24670 3726 24722
rect 3778 24670 3790 24722
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 7746 24670 7758 24722
rect 7810 24670 7822 24722
rect 10210 24670 10222 24722
rect 10274 24670 10286 24722
rect 12114 24670 12126 24722
rect 12178 24670 12190 24722
rect 17490 24670 17502 24722
rect 17554 24670 17566 24722
rect 18946 24670 18958 24722
rect 19010 24670 19022 24722
rect 22866 24670 22878 24722
rect 22930 24670 22942 24722
rect 2942 24658 2994 24670
rect 8990 24658 9042 24670
rect 11566 24658 11618 24670
rect 18398 24658 18450 24670
rect 23214 24658 23266 24670
rect 28590 24722 28642 24734
rect 29250 24670 29262 24722
rect 29314 24670 29326 24722
rect 28590 24658 28642 24670
rect 1934 24610 1986 24622
rect 11342 24610 11394 24622
rect 25342 24610 25394 24622
rect 9762 24558 9774 24610
rect 9826 24558 9838 24610
rect 15922 24558 15934 24610
rect 15986 24558 15998 24610
rect 17602 24558 17614 24610
rect 17666 24558 17678 24610
rect 1934 24546 1986 24558
rect 11342 24546 11394 24558
rect 25342 24546 25394 24558
rect 25790 24610 25842 24622
rect 28030 24610 28082 24622
rect 26226 24558 26238 24610
rect 26290 24558 26302 24610
rect 28354 24558 28366 24610
rect 28418 24558 28430 24610
rect 25790 24546 25842 24558
rect 28030 24546 28082 24558
rect 2158 24498 2210 24510
rect 2158 24434 2210 24446
rect 4174 24498 4226 24510
rect 4174 24434 4226 24446
rect 1344 24330 32592 24364
rect 1344 24278 5120 24330
rect 5172 24278 5224 24330
rect 5276 24278 5328 24330
rect 5380 24278 12932 24330
rect 12984 24278 13036 24330
rect 13088 24278 13140 24330
rect 13192 24278 20744 24330
rect 20796 24278 20848 24330
rect 20900 24278 20952 24330
rect 21004 24278 28556 24330
rect 28608 24278 28660 24330
rect 28712 24278 28764 24330
rect 28816 24278 32592 24330
rect 1344 24244 32592 24278
rect 13022 24162 13074 24174
rect 13022 24098 13074 24110
rect 17054 24162 17106 24174
rect 17054 24098 17106 24110
rect 20862 24162 20914 24174
rect 20862 24098 20914 24110
rect 22990 24162 23042 24174
rect 22990 24098 23042 24110
rect 27134 24162 27186 24174
rect 27134 24098 27186 24110
rect 4510 24050 4562 24062
rect 6302 24050 6354 24062
rect 8654 24050 8706 24062
rect 4050 23998 4062 24050
rect 4114 23998 4126 24050
rect 5954 23998 5966 24050
rect 6018 23998 6030 24050
rect 8082 23998 8094 24050
rect 8146 23998 8158 24050
rect 4510 23986 4562 23998
rect 6302 23986 6354 23998
rect 8654 23986 8706 23998
rect 21646 24050 21698 24062
rect 27794 23998 27806 24050
rect 27858 23998 27870 24050
rect 30146 23998 30158 24050
rect 30210 23998 30222 24050
rect 21646 23986 21698 23998
rect 5070 23938 5122 23950
rect 2034 23886 2046 23938
rect 2098 23886 2110 23938
rect 5070 23874 5122 23886
rect 9550 23938 9602 23950
rect 17166 23938 17218 23950
rect 9986 23886 9998 23938
rect 10050 23886 10062 23938
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 22082 23886 22094 23938
rect 22146 23886 22158 23938
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 9550 23874 9602 23886
rect 17166 23874 17218 23886
rect 32062 23826 32114 23838
rect 3042 23774 3054 23826
rect 3106 23774 3118 23826
rect 7074 23774 7086 23826
rect 7138 23774 7150 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 31490 23774 31502 23826
rect 31554 23774 31566 23826
rect 32062 23762 32114 23774
rect 2270 23714 2322 23726
rect 2270 23650 2322 23662
rect 9102 23714 9154 23726
rect 27358 23714 27410 23726
rect 12450 23662 12462 23714
rect 12514 23662 12526 23714
rect 16370 23662 16382 23714
rect 16434 23662 16446 23714
rect 20290 23662 20302 23714
rect 20354 23662 20366 23714
rect 26562 23662 26574 23714
rect 26626 23662 26638 23714
rect 9102 23650 9154 23662
rect 27358 23650 27410 23662
rect 1344 23546 32752 23580
rect 1344 23494 9026 23546
rect 9078 23494 9130 23546
rect 9182 23494 9234 23546
rect 9286 23494 16838 23546
rect 16890 23494 16942 23546
rect 16994 23494 17046 23546
rect 17098 23494 24650 23546
rect 24702 23494 24754 23546
rect 24806 23494 24858 23546
rect 24910 23494 32462 23546
rect 32514 23494 32566 23546
rect 32618 23494 32670 23546
rect 32722 23494 32752 23546
rect 1344 23460 32752 23494
rect 4174 23378 4226 23390
rect 15150 23378 15202 23390
rect 7410 23326 7422 23378
rect 7474 23326 7486 23378
rect 13346 23326 13358 23378
rect 13410 23326 13422 23378
rect 4174 23314 4226 23326
rect 15150 23314 15202 23326
rect 17726 23378 17778 23390
rect 17726 23314 17778 23326
rect 8654 23266 8706 23278
rect 9886 23266 9938 23278
rect 18398 23266 18450 23278
rect 1810 23214 1822 23266
rect 1874 23214 1886 23266
rect 9538 23214 9550 23266
rect 9602 23214 9614 23266
rect 18050 23214 18062 23266
rect 18114 23214 18126 23266
rect 8654 23202 8706 23214
rect 9886 23202 9938 23214
rect 18398 23202 18450 23214
rect 18734 23266 18786 23278
rect 28914 23214 28926 23266
rect 28978 23214 28990 23266
rect 18734 23202 18786 23214
rect 4622 23154 4674 23166
rect 10222 23154 10274 23166
rect 4946 23102 4958 23154
rect 5010 23102 5022 23154
rect 10770 23102 10782 23154
rect 10834 23102 10846 23154
rect 14130 23102 14142 23154
rect 14194 23102 14206 23154
rect 17490 23102 17502 23154
rect 17554 23102 17566 23154
rect 20850 23102 20862 23154
rect 20914 23102 20926 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 32162 23102 32174 23154
rect 32226 23102 32238 23154
rect 4622 23090 4674 23102
rect 10222 23090 10274 23102
rect 3042 22990 3054 23042
rect 3106 22990 3118 23042
rect 8418 22990 8430 23042
rect 8482 22990 8494 23042
rect 18946 22990 18958 23042
rect 19010 22990 19022 23042
rect 22306 22990 22318 23042
rect 22370 22990 22382 23042
rect 31490 22990 31502 23042
rect 31554 22990 31566 23042
rect 8094 22930 8146 22942
rect 8094 22866 8146 22878
rect 13918 22930 13970 22942
rect 13918 22866 13970 22878
rect 1344 22762 32592 22796
rect 1344 22710 5120 22762
rect 5172 22710 5224 22762
rect 5276 22710 5328 22762
rect 5380 22710 12932 22762
rect 12984 22710 13036 22762
rect 13088 22710 13140 22762
rect 13192 22710 20744 22762
rect 20796 22710 20848 22762
rect 20900 22710 20952 22762
rect 21004 22710 28556 22762
rect 28608 22710 28660 22762
rect 28712 22710 28764 22762
rect 28816 22710 32592 22762
rect 1344 22676 32592 22710
rect 19630 22594 19682 22606
rect 19630 22530 19682 22542
rect 21198 22594 21250 22606
rect 21198 22530 21250 22542
rect 25006 22594 25058 22606
rect 25006 22530 25058 22542
rect 2270 22482 2322 22494
rect 5070 22482 5122 22494
rect 2034 22430 2046 22482
rect 2098 22430 2110 22482
rect 4050 22430 4062 22482
rect 4114 22430 4126 22482
rect 8530 22430 8542 22482
rect 8594 22430 8606 22482
rect 14018 22430 14030 22482
rect 14082 22430 14094 22482
rect 30146 22430 30158 22482
rect 30210 22430 30222 22482
rect 2270 22418 2322 22430
rect 5070 22418 5122 22430
rect 13582 22370 13634 22382
rect 11554 22318 11566 22370
rect 11618 22318 11630 22370
rect 12786 22318 12798 22370
rect 12850 22318 12862 22370
rect 13582 22306 13634 22318
rect 15038 22370 15090 22382
rect 15038 22306 15090 22318
rect 16158 22370 16210 22382
rect 24670 22370 24722 22382
rect 28702 22370 28754 22382
rect 16482 22318 16494 22370
rect 16546 22318 16558 22370
rect 20514 22318 20526 22370
rect 20578 22318 20590 22370
rect 24210 22318 24222 22370
rect 24274 22318 24286 22370
rect 28130 22318 28142 22370
rect 28194 22318 28206 22370
rect 16158 22306 16210 22318
rect 24670 22306 24722 22318
rect 28702 22306 28754 22318
rect 6190 22258 6242 22270
rect 2818 22206 2830 22258
rect 2882 22206 2894 22258
rect 5842 22206 5854 22258
rect 5906 22206 5918 22258
rect 12562 22206 12574 22258
rect 12626 22206 12638 22258
rect 15362 22206 15374 22258
rect 15426 22206 15438 22258
rect 20738 22206 20750 22258
rect 20802 22206 20814 22258
rect 31154 22206 31166 22258
rect 31218 22206 31230 22258
rect 6190 22194 6242 22206
rect 4622 22146 4674 22158
rect 4622 22082 4674 22094
rect 6526 22146 6578 22158
rect 6526 22082 6578 22094
rect 14702 22146 14754 22158
rect 19966 22146 20018 22158
rect 18946 22094 18958 22146
rect 19010 22094 19022 22146
rect 21970 22094 21982 22146
rect 22034 22094 22046 22146
rect 25554 22094 25566 22146
rect 25618 22094 25630 22146
rect 14702 22082 14754 22094
rect 19966 22082 20018 22094
rect 1344 21978 32752 22012
rect 1344 21926 9026 21978
rect 9078 21926 9130 21978
rect 9182 21926 9234 21978
rect 9286 21926 16838 21978
rect 16890 21926 16942 21978
rect 16994 21926 17046 21978
rect 17098 21926 24650 21978
rect 24702 21926 24754 21978
rect 24806 21926 24858 21978
rect 24910 21926 32462 21978
rect 32514 21926 32566 21978
rect 32618 21926 32670 21978
rect 32722 21926 32752 21978
rect 1344 21892 32752 21926
rect 10334 21810 10386 21822
rect 8530 21758 8542 21810
rect 8594 21758 8606 21810
rect 10334 21746 10386 21758
rect 16718 21810 16770 21822
rect 16718 21746 16770 21758
rect 18062 21810 18114 21822
rect 21982 21810 22034 21822
rect 21186 21758 21198 21810
rect 21250 21758 21262 21810
rect 18062 21746 18114 21758
rect 21982 21746 22034 21758
rect 25118 21810 25170 21822
rect 25666 21758 25678 21810
rect 25730 21758 25742 21810
rect 25118 21746 25170 21758
rect 2382 21698 2434 21710
rect 4622 21698 4674 21710
rect 3154 21646 3166 21698
rect 3218 21646 3230 21698
rect 2382 21634 2434 21646
rect 4622 21634 4674 21646
rect 9886 21698 9938 21710
rect 11778 21646 11790 21698
rect 11842 21646 11854 21698
rect 24434 21646 24446 21698
rect 24498 21646 24510 21698
rect 31042 21646 31054 21698
rect 31106 21646 31118 21698
rect 9886 21634 9938 21646
rect 5630 21586 5682 21598
rect 9102 21586 9154 21598
rect 2146 21534 2158 21586
rect 2210 21534 2222 21586
rect 5954 21534 5966 21586
rect 6018 21534 6030 21586
rect 9538 21534 9550 21586
rect 9602 21534 9614 21586
rect 10546 21534 10558 21586
rect 10610 21534 10622 21586
rect 16258 21534 16270 21586
rect 16322 21534 16334 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 18946 21534 18958 21586
rect 19010 21534 19022 21586
rect 28242 21534 28254 21586
rect 28306 21534 28318 21586
rect 28690 21534 28702 21586
rect 28754 21534 28766 21586
rect 5630 21522 5682 21534
rect 9102 21522 9154 21534
rect 22318 21474 22370 21486
rect 4162 21422 4174 21474
rect 4226 21422 4238 21474
rect 22318 21410 22370 21422
rect 22766 21474 22818 21486
rect 32174 21474 32226 21486
rect 23202 21422 23214 21474
rect 23266 21422 23278 21474
rect 30034 21422 30046 21474
rect 30098 21422 30110 21474
rect 31938 21422 31950 21474
rect 32002 21422 32014 21474
rect 22766 21410 22818 21422
rect 32174 21410 32226 21422
rect 1344 21194 32592 21228
rect 1344 21142 5120 21194
rect 5172 21142 5224 21194
rect 5276 21142 5328 21194
rect 5380 21142 12932 21194
rect 12984 21142 13036 21194
rect 13088 21142 13140 21194
rect 13192 21142 20744 21194
rect 20796 21142 20848 21194
rect 20900 21142 20952 21194
rect 21004 21142 28556 21194
rect 28608 21142 28660 21194
rect 28712 21142 28764 21194
rect 28816 21142 32592 21194
rect 1344 21108 32592 21142
rect 12238 21026 12290 21038
rect 12238 20962 12290 20974
rect 5742 20914 5794 20926
rect 14254 20914 14306 20926
rect 21870 20914 21922 20926
rect 26686 20914 26738 20926
rect 31502 20914 31554 20926
rect 4050 20862 4062 20914
rect 4114 20862 4126 20914
rect 6850 20862 6862 20914
rect 6914 20862 6926 20914
rect 20514 20862 20526 20914
rect 20578 20862 20590 20914
rect 22082 20862 22094 20914
rect 22146 20862 22158 20914
rect 27906 20862 27918 20914
rect 27970 20862 27982 20914
rect 30594 20862 30606 20914
rect 30658 20862 30670 20914
rect 5742 20850 5794 20862
rect 14254 20850 14306 20862
rect 21870 20850 21922 20862
rect 26686 20850 26738 20862
rect 31502 20850 31554 20862
rect 8766 20802 8818 20814
rect 13806 20802 13858 20814
rect 19070 20802 19122 20814
rect 2034 20750 2046 20802
rect 2098 20750 2110 20802
rect 9090 20750 9102 20802
rect 9154 20750 9166 20802
rect 12562 20750 12574 20802
rect 12626 20750 12638 20802
rect 15138 20750 15150 20802
rect 15202 20750 15214 20802
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 22978 20750 22990 20802
rect 23042 20750 23054 20802
rect 8766 20738 8818 20750
rect 13806 20738 13858 20750
rect 19070 20738 19122 20750
rect 2270 20690 2322 20702
rect 11454 20690 11506 20702
rect 3042 20638 3054 20690
rect 3106 20638 3118 20690
rect 8194 20638 8206 20690
rect 8258 20638 8270 20690
rect 2270 20626 2322 20638
rect 11454 20626 11506 20638
rect 12798 20690 12850 20702
rect 20750 20690 20802 20702
rect 13458 20638 13470 20690
rect 13522 20638 13534 20690
rect 12798 20626 12850 20638
rect 20750 20626 20802 20638
rect 21422 20690 21474 20702
rect 26338 20638 26350 20690
rect 26402 20638 26414 20690
rect 29474 20638 29486 20690
rect 29538 20638 29550 20690
rect 21422 20626 21474 20638
rect 4622 20578 4674 20590
rect 4622 20514 4674 20526
rect 6414 20578 6466 20590
rect 6414 20514 6466 20526
rect 17502 20578 17554 20590
rect 26126 20578 26178 20590
rect 25554 20526 25566 20578
rect 25618 20526 25630 20578
rect 17502 20514 17554 20526
rect 26126 20514 26178 20526
rect 27358 20578 27410 20590
rect 27358 20514 27410 20526
rect 1344 20410 32752 20444
rect 1344 20358 9026 20410
rect 9078 20358 9130 20410
rect 9182 20358 9234 20410
rect 9286 20358 16838 20410
rect 16890 20358 16942 20410
rect 16994 20358 17046 20410
rect 17098 20358 24650 20410
rect 24702 20358 24754 20410
rect 24806 20358 24858 20410
rect 24910 20358 32462 20410
rect 32514 20358 32566 20410
rect 32618 20358 32670 20410
rect 32722 20358 32752 20410
rect 1344 20324 32752 20358
rect 23102 20242 23154 20254
rect 8418 20190 8430 20242
rect 8482 20190 8494 20242
rect 15362 20190 15374 20242
rect 15426 20190 15438 20242
rect 23102 20178 23154 20190
rect 2382 20130 2434 20142
rect 12014 20130 12066 20142
rect 9650 20078 9662 20130
rect 9714 20078 9726 20130
rect 2382 20066 2434 20078
rect 12014 20066 12066 20078
rect 15934 20130 15986 20142
rect 25342 20130 25394 20142
rect 19394 20078 19406 20130
rect 19458 20078 19470 20130
rect 22194 20078 22206 20130
rect 22258 20078 22270 20130
rect 23426 20078 23438 20130
rect 23490 20078 23502 20130
rect 15934 20066 15986 20078
rect 25342 20066 25394 20078
rect 28478 20130 28530 20142
rect 28478 20066 28530 20078
rect 29262 20130 29314 20142
rect 31490 20078 31502 20130
rect 31554 20078 31566 20130
rect 29262 20066 29314 20078
rect 5294 20018 5346 20030
rect 4722 19966 4734 20018
rect 4786 19966 4798 20018
rect 5294 19954 5346 19966
rect 5630 20018 5682 20030
rect 12238 20018 12290 20030
rect 25566 20018 25618 20030
rect 5954 19966 5966 20018
rect 6018 19966 6030 20018
rect 12786 19966 12798 20018
rect 12850 19966 12862 20018
rect 26226 19966 26238 20018
rect 26290 19966 26302 20018
rect 5630 19954 5682 19966
rect 12238 19954 12290 19966
rect 25566 19954 25618 19966
rect 9102 19906 9154 19918
rect 11454 19906 11506 19918
rect 16830 19906 16882 19918
rect 10994 19854 11006 19906
rect 11058 19854 11070 19906
rect 16482 19854 16494 19906
rect 16546 19854 16558 19906
rect 9102 19842 9154 19854
rect 11454 19842 11506 19854
rect 16830 19842 16882 19854
rect 17502 19906 17554 19918
rect 20974 19906 21026 19918
rect 18386 19854 18398 19906
rect 18450 19854 18462 19906
rect 21186 19854 21198 19906
rect 21250 19854 21262 19906
rect 24322 19854 24334 19906
rect 24386 19854 24398 19906
rect 30482 19854 30494 19906
rect 30546 19854 30558 19906
rect 17502 19842 17554 19854
rect 20974 19842 21026 19854
rect 1598 19794 1650 19806
rect 1598 19730 1650 19742
rect 1344 19626 32592 19660
rect 1344 19574 5120 19626
rect 5172 19574 5224 19626
rect 5276 19574 5328 19626
rect 5380 19574 12932 19626
rect 12984 19574 13036 19626
rect 13088 19574 13140 19626
rect 13192 19574 20744 19626
rect 20796 19574 20848 19626
rect 20900 19574 20952 19626
rect 21004 19574 28556 19626
rect 28608 19574 28660 19626
rect 28712 19574 28764 19626
rect 28816 19574 32592 19626
rect 1344 19540 32592 19574
rect 14478 19458 14530 19470
rect 12226 19406 12238 19458
rect 12290 19455 12302 19458
rect 13010 19455 13022 19458
rect 12290 19409 13022 19455
rect 12290 19406 12302 19409
rect 13010 19406 13022 19409
rect 13074 19406 13086 19458
rect 14478 19394 14530 19406
rect 24894 19458 24946 19470
rect 24894 19394 24946 19406
rect 4510 19346 4562 19358
rect 4050 19294 4062 19346
rect 4114 19294 4126 19346
rect 4510 19282 4562 19294
rect 9774 19346 9826 19358
rect 12462 19346 12514 19358
rect 11890 19294 11902 19346
rect 11954 19294 11966 19346
rect 9774 19282 9826 19294
rect 12462 19282 12514 19294
rect 12910 19346 12962 19358
rect 30146 19294 30158 19346
rect 30210 19294 30222 19346
rect 12910 19282 12962 19294
rect 21198 19234 21250 19246
rect 25006 19234 25058 19246
rect 28702 19234 28754 19246
rect 2034 19182 2046 19234
rect 2098 19182 2110 19234
rect 5618 19182 5630 19234
rect 5682 19182 5694 19234
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 13682 19182 13694 19234
rect 13746 19182 13758 19234
rect 17602 19182 17614 19234
rect 17666 19182 17678 19234
rect 18050 19182 18062 19234
rect 18114 19182 18126 19234
rect 18946 19182 18958 19234
rect 19010 19182 19022 19234
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 21198 19170 21250 19182
rect 25006 19170 25058 19182
rect 28702 19170 28754 19182
rect 13470 19122 13522 19134
rect 2706 19070 2718 19122
rect 2770 19070 2782 19122
rect 10882 19070 10894 19122
rect 10946 19070 10958 19122
rect 13470 19058 13522 19070
rect 15262 19122 15314 19134
rect 15262 19058 15314 19070
rect 19182 19122 19234 19134
rect 20750 19122 20802 19134
rect 19506 19070 19518 19122
rect 19570 19070 19582 19122
rect 31154 19070 31166 19122
rect 31218 19070 31230 19122
rect 19182 19058 19234 19070
rect 20750 19058 20802 19070
rect 2046 19010 2098 19022
rect 9214 19010 9266 19022
rect 8642 18958 8654 19010
rect 8706 18958 8718 19010
rect 2046 18946 2098 18958
rect 9214 18946 9266 18958
rect 9886 19010 9938 19022
rect 9886 18946 9938 18958
rect 18510 19010 18562 19022
rect 29262 19010 29314 19022
rect 24322 18958 24334 19010
rect 24386 18958 24398 19010
rect 27906 18958 27918 19010
rect 27970 18958 27982 19010
rect 18510 18946 18562 18958
rect 29262 18946 29314 18958
rect 32062 19010 32114 19022
rect 32062 18946 32114 18958
rect 1344 18842 32752 18876
rect 1344 18790 9026 18842
rect 9078 18790 9130 18842
rect 9182 18790 9234 18842
rect 9286 18790 16838 18842
rect 16890 18790 16942 18842
rect 16994 18790 17046 18842
rect 17098 18790 24650 18842
rect 24702 18790 24754 18842
rect 24806 18790 24858 18842
rect 24910 18790 32462 18842
rect 32514 18790 32566 18842
rect 32618 18790 32670 18842
rect 32722 18790 32752 18842
rect 1344 18756 32752 18790
rect 1934 18674 1986 18686
rect 1934 18610 1986 18622
rect 2158 18674 2210 18686
rect 2158 18610 2210 18622
rect 9438 18674 9490 18686
rect 16370 18622 16382 18674
rect 16434 18622 16446 18674
rect 28130 18622 28142 18674
rect 28194 18622 28206 18674
rect 9438 18610 9490 18622
rect 6414 18562 6466 18574
rect 6414 18498 6466 18510
rect 10222 18562 10274 18574
rect 10222 18498 10274 18510
rect 17390 18562 17442 18574
rect 17390 18498 17442 18510
rect 21310 18562 21362 18574
rect 31838 18562 31890 18574
rect 24322 18510 24334 18562
rect 24386 18510 24398 18562
rect 26674 18510 26686 18562
rect 26738 18510 26750 18562
rect 27346 18510 27358 18562
rect 27410 18510 27422 18562
rect 21310 18498 21362 18510
rect 31838 18498 31890 18510
rect 2942 18450 2994 18462
rect 2942 18386 2994 18398
rect 3726 18450 3778 18462
rect 7422 18450 7474 18462
rect 4050 18398 4062 18450
rect 4114 18398 4126 18450
rect 3726 18386 3778 18398
rect 7422 18386 7474 18398
rect 8990 18450 9042 18462
rect 13246 18450 13298 18462
rect 22430 18450 22482 18462
rect 31278 18450 31330 18462
rect 12450 18398 12462 18450
rect 12514 18398 12526 18450
rect 13010 18398 13022 18450
rect 13074 18398 13086 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 17602 18398 17614 18450
rect 17666 18398 17678 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 19058 18398 19070 18450
rect 19122 18398 19134 18450
rect 22866 18398 22878 18450
rect 22930 18398 22942 18450
rect 24546 18398 24558 18450
rect 24610 18398 24622 18450
rect 25554 18398 25566 18450
rect 25618 18398 25630 18450
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 27122 18398 27134 18450
rect 27186 18398 27198 18450
rect 30594 18398 30606 18450
rect 30658 18398 30670 18450
rect 31490 18398 31502 18450
rect 31554 18398 31566 18450
rect 8990 18386 9042 18398
rect 13246 18386 13298 18398
rect 22430 18386 22482 18398
rect 31278 18386 31330 18398
rect 18174 18338 18226 18350
rect 27582 18338 27634 18350
rect 7858 18286 7870 18338
rect 7922 18286 7934 18338
rect 25666 18286 25678 18338
rect 25730 18286 25742 18338
rect 18174 18274 18226 18286
rect 27582 18274 27634 18286
rect 7198 18226 7250 18238
rect 7198 18162 7250 18174
rect 16942 18226 16994 18238
rect 16942 18162 16994 18174
rect 22094 18226 22146 18238
rect 22094 18162 22146 18174
rect 23326 18226 23378 18238
rect 23326 18162 23378 18174
rect 1344 18058 32592 18092
rect 1344 18006 5120 18058
rect 5172 18006 5224 18058
rect 5276 18006 5328 18058
rect 5380 18006 12932 18058
rect 12984 18006 13036 18058
rect 13088 18006 13140 18058
rect 13192 18006 20744 18058
rect 20796 18006 20848 18058
rect 20900 18006 20952 18058
rect 21004 18006 28556 18058
rect 28608 18006 28660 18058
rect 28712 18006 28764 18058
rect 28816 18006 32592 18058
rect 1344 17972 32592 18006
rect 20302 17890 20354 17902
rect 20302 17826 20354 17838
rect 1934 17778 1986 17790
rect 4510 17778 4562 17790
rect 3938 17726 3950 17778
rect 4002 17726 4014 17778
rect 1934 17714 1986 17726
rect 4510 17714 4562 17726
rect 5070 17778 5122 17790
rect 5070 17714 5122 17726
rect 5742 17778 5794 17790
rect 7422 17778 7474 17790
rect 6402 17726 6414 17778
rect 6466 17726 6478 17778
rect 5742 17714 5794 17726
rect 7422 17714 7474 17726
rect 11678 17778 11730 17790
rect 20750 17778 20802 17790
rect 26574 17778 26626 17790
rect 32062 17778 32114 17790
rect 12114 17726 12126 17778
rect 12178 17726 12190 17778
rect 15362 17726 15374 17778
rect 15426 17726 15438 17778
rect 21298 17726 21310 17778
rect 21362 17726 21374 17778
rect 30146 17726 30158 17778
rect 30210 17726 30222 17778
rect 11678 17714 11730 17726
rect 20750 17714 20802 17726
rect 26574 17714 26626 17726
rect 32062 17714 32114 17726
rect 7646 17666 7698 17678
rect 16606 17666 16658 17678
rect 22654 17666 22706 17678
rect 27358 17666 27410 17678
rect 29262 17666 29314 17678
rect 8194 17614 8206 17666
rect 8258 17614 8270 17666
rect 12338 17614 12350 17666
rect 12402 17614 12414 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 21522 17614 21534 17666
rect 21586 17614 21598 17666
rect 22194 17614 22206 17666
rect 22258 17614 22270 17666
rect 23314 17614 23326 17666
rect 23378 17614 23390 17666
rect 28578 17614 28590 17666
rect 28642 17614 28654 17666
rect 7646 17602 7698 17614
rect 16606 17602 16658 17614
rect 22654 17602 22706 17614
rect 27358 17602 27410 17614
rect 29262 17602 29314 17614
rect 10558 17554 10610 17566
rect 19518 17554 19570 17566
rect 26350 17554 26402 17566
rect 2258 17502 2270 17554
rect 2322 17502 2334 17554
rect 3042 17502 3054 17554
rect 3106 17502 3118 17554
rect 14354 17502 14366 17554
rect 14418 17502 14430 17554
rect 21970 17502 21982 17554
rect 22034 17502 22046 17554
rect 26898 17502 26910 17554
rect 26962 17502 26974 17554
rect 28354 17502 28366 17554
rect 28418 17502 28430 17554
rect 31154 17502 31166 17554
rect 31218 17502 31230 17554
rect 10558 17490 10610 17502
rect 19518 17490 19570 17502
rect 26350 17490 26402 17502
rect 6862 17442 6914 17454
rect 6862 17378 6914 17390
rect 11342 17442 11394 17454
rect 11342 17378 11394 17390
rect 12910 17442 12962 17454
rect 12910 17378 12962 17390
rect 13582 17442 13634 17454
rect 13582 17378 13634 17390
rect 15822 17442 15874 17454
rect 15822 17378 15874 17390
rect 16270 17442 16322 17454
rect 29710 17442 29762 17454
rect 25666 17390 25678 17442
rect 25730 17390 25742 17442
rect 16270 17378 16322 17390
rect 29710 17378 29762 17390
rect 1344 17274 32752 17308
rect 1344 17222 9026 17274
rect 9078 17222 9130 17274
rect 9182 17222 9234 17274
rect 9286 17222 16838 17274
rect 16890 17222 16942 17274
rect 16994 17222 17046 17274
rect 17098 17222 24650 17274
rect 24702 17222 24754 17274
rect 24806 17222 24858 17274
rect 24910 17222 32462 17274
rect 32514 17222 32566 17274
rect 32618 17222 32670 17274
rect 32722 17222 32752 17274
rect 1344 17188 32752 17222
rect 1598 17106 1650 17118
rect 5406 17106 5458 17118
rect 16830 17106 16882 17118
rect 29150 17106 29202 17118
rect 2258 17054 2270 17106
rect 2322 17054 2334 17106
rect 14354 17054 14366 17106
rect 14418 17054 14430 17106
rect 28018 17054 28030 17106
rect 28082 17054 28094 17106
rect 1598 17042 1650 17054
rect 5406 17042 5458 17054
rect 16830 17042 16882 17054
rect 29150 17042 29202 17054
rect 6190 16994 6242 17006
rect 11006 16994 11058 17006
rect 22990 16994 23042 17006
rect 10658 16942 10670 16994
rect 10722 16942 10734 16994
rect 15250 16942 15262 16994
rect 15314 16942 15326 16994
rect 6190 16930 6242 16942
rect 11006 16930 11058 16942
rect 22990 16930 23042 16942
rect 23326 16994 23378 17006
rect 23326 16930 23378 16942
rect 23662 16994 23714 17006
rect 23662 16930 23714 16942
rect 24334 16994 24386 17006
rect 31042 16942 31054 16994
rect 31106 16942 31118 16994
rect 31826 16942 31838 16994
rect 31890 16942 31902 16994
rect 24334 16930 24386 16942
rect 5294 16882 5346 16894
rect 8878 16882 8930 16894
rect 11454 16882 11506 16894
rect 25342 16882 25394 16894
rect 4722 16830 4734 16882
rect 4786 16830 4798 16882
rect 8418 16830 8430 16882
rect 8482 16830 8494 16882
rect 9762 16830 9774 16882
rect 9826 16830 9838 16882
rect 11778 16830 11790 16882
rect 11842 16830 11854 16882
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 16146 16830 16158 16882
rect 16210 16830 16222 16882
rect 17490 16830 17502 16882
rect 17554 16830 17566 16882
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 32050 16830 32062 16882
rect 32114 16830 32126 16882
rect 5294 16818 5346 16830
rect 8878 16818 8930 16830
rect 11454 16818 11506 16830
rect 25342 16818 25394 16830
rect 21634 16718 21646 16770
rect 21698 16718 21710 16770
rect 23986 16718 23998 16770
rect 24050 16718 24062 16770
rect 24658 16718 24670 16770
rect 24722 16718 24734 16770
rect 30034 16718 30046 16770
rect 30098 16718 30110 16770
rect 9662 16658 9714 16670
rect 9662 16594 9714 16606
rect 14926 16658 14978 16670
rect 14926 16594 14978 16606
rect 28814 16658 28866 16670
rect 28814 16594 28866 16606
rect 1344 16490 32592 16524
rect 1344 16438 5120 16490
rect 5172 16438 5224 16490
rect 5276 16438 5328 16490
rect 5380 16438 12932 16490
rect 12984 16438 13036 16490
rect 13088 16438 13140 16490
rect 13192 16438 20744 16490
rect 20796 16438 20848 16490
rect 20900 16438 20952 16490
rect 21004 16438 28556 16490
rect 28608 16438 28660 16490
rect 28712 16438 28764 16490
rect 28816 16438 32592 16490
rect 1344 16404 32592 16438
rect 13918 16322 13970 16334
rect 13918 16258 13970 16270
rect 25006 16322 25058 16334
rect 29810 16319 29822 16322
rect 25006 16258 25058 16270
rect 29153 16273 29822 16319
rect 4734 16210 4786 16222
rect 3938 16158 3950 16210
rect 4002 16158 4014 16210
rect 4734 16146 4786 16158
rect 5070 16210 5122 16222
rect 5070 16146 5122 16158
rect 6974 16210 7026 16222
rect 6974 16146 7026 16158
rect 13022 16210 13074 16222
rect 29153 16210 29199 16273
rect 29810 16270 29822 16273
rect 29874 16270 29886 16322
rect 29262 16210 29314 16222
rect 19394 16158 19406 16210
rect 19458 16158 19470 16210
rect 29138 16158 29150 16210
rect 29202 16158 29214 16210
rect 13022 16146 13074 16158
rect 29262 16146 29314 16158
rect 29822 16210 29874 16222
rect 32062 16210 32114 16222
rect 30146 16158 30158 16210
rect 30210 16158 30222 16210
rect 29822 16146 29874 16158
rect 32062 16146 32114 16158
rect 1934 16098 1986 16110
rect 11902 16098 11954 16110
rect 15486 16098 15538 16110
rect 21422 16098 21474 16110
rect 28702 16098 28754 16110
rect 5954 16046 5966 16098
rect 6018 16046 6030 16098
rect 7410 16046 7422 16098
rect 7474 16046 7486 16098
rect 11218 16046 11230 16098
rect 11282 16046 11294 16098
rect 14802 16046 14814 16098
rect 14866 16046 14878 16098
rect 16146 16046 16158 16098
rect 16210 16046 16222 16098
rect 19618 16046 19630 16098
rect 19682 16046 19694 16098
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 21858 16046 21870 16098
rect 21922 16046 21934 16098
rect 28130 16046 28142 16098
rect 28194 16046 28206 16098
rect 1934 16034 1986 16046
rect 11902 16034 11954 16046
rect 15486 16034 15538 16046
rect 21422 16034 21474 16046
rect 28702 16034 28754 16046
rect 12126 15986 12178 15998
rect 3042 15934 3054 15986
rect 3106 15934 3118 15986
rect 12126 15922 12178 15934
rect 12462 15986 12514 15998
rect 24894 15986 24946 15998
rect 20066 15934 20078 15986
rect 20130 15934 20142 15986
rect 31154 15934 31166 15986
rect 31218 15934 31230 15986
rect 12462 15922 12514 15934
rect 24894 15922 24946 15934
rect 2270 15874 2322 15886
rect 2270 15810 2322 15822
rect 5742 15874 5794 15886
rect 5742 15810 5794 15822
rect 7310 15874 7362 15886
rect 7310 15810 7362 15822
rect 8206 15874 8258 15886
rect 19182 15874 19234 15886
rect 8978 15822 8990 15874
rect 9042 15822 9054 15874
rect 18386 15822 18398 15874
rect 18450 15822 18462 15874
rect 24098 15822 24110 15874
rect 24162 15822 24174 15874
rect 25554 15822 25566 15874
rect 25618 15822 25630 15874
rect 8206 15810 8258 15822
rect 19182 15810 19234 15822
rect 1344 15706 32752 15740
rect 1344 15654 9026 15706
rect 9078 15654 9130 15706
rect 9182 15654 9234 15706
rect 9286 15654 16838 15706
rect 16890 15654 16942 15706
rect 16994 15654 17046 15706
rect 17098 15654 24650 15706
rect 24702 15654 24754 15706
rect 24806 15654 24858 15706
rect 24910 15654 32462 15706
rect 32514 15654 32566 15706
rect 32618 15654 32670 15706
rect 32722 15654 32752 15706
rect 1344 15620 32752 15654
rect 8990 15538 9042 15550
rect 2146 15486 2158 15538
rect 2210 15486 2222 15538
rect 8990 15474 9042 15486
rect 9886 15538 9938 15550
rect 18062 15538 18114 15550
rect 22542 15538 22594 15550
rect 12562 15486 12574 15538
rect 12626 15486 12638 15538
rect 21522 15486 21534 15538
rect 21586 15486 21598 15538
rect 9886 15474 9938 15486
rect 18062 15474 18114 15486
rect 22542 15474 22594 15486
rect 24110 15538 24162 15550
rect 24110 15474 24162 15486
rect 26126 15538 26178 15550
rect 26898 15486 26910 15538
rect 26962 15486 26974 15538
rect 26126 15474 26178 15486
rect 18174 15426 18226 15438
rect 6178 15374 6190 15426
rect 6242 15374 6254 15426
rect 6626 15374 6638 15426
rect 6690 15374 6702 15426
rect 10882 15374 10894 15426
rect 10946 15374 10958 15426
rect 18174 15362 18226 15374
rect 22878 15426 22930 15438
rect 22878 15362 22930 15374
rect 23214 15426 23266 15438
rect 24334 15426 24386 15438
rect 23538 15374 23550 15426
rect 23602 15374 23614 15426
rect 23214 15362 23266 15374
rect 24334 15362 24386 15374
rect 24670 15426 24722 15438
rect 24670 15362 24722 15374
rect 5070 15314 5122 15326
rect 8542 15314 8594 15326
rect 15486 15314 15538 15326
rect 18622 15314 18674 15326
rect 29822 15314 29874 15326
rect 4610 15262 4622 15314
rect 4674 15262 4686 15314
rect 5954 15262 5966 15314
rect 6018 15262 6030 15314
rect 9762 15262 9774 15314
rect 9826 15262 9838 15314
rect 11106 15262 11118 15314
rect 11170 15262 11182 15314
rect 14802 15262 14814 15314
rect 14866 15262 14878 15314
rect 16482 15262 16494 15314
rect 16546 15262 16558 15314
rect 19058 15262 19070 15314
rect 19122 15262 19134 15314
rect 25442 15262 25454 15314
rect 25506 15262 25518 15314
rect 29362 15262 29374 15314
rect 29426 15262 29438 15314
rect 30706 15262 30718 15314
rect 30770 15262 30782 15314
rect 31602 15262 31614 15314
rect 31666 15262 31678 15314
rect 5070 15250 5122 15262
rect 8542 15250 8594 15262
rect 15486 15250 15538 15262
rect 18622 15250 18674 15262
rect 29822 15250 29874 15262
rect 17502 15202 17554 15214
rect 7970 15150 7982 15202
rect 8034 15150 8046 15202
rect 16034 15150 16046 15202
rect 16098 15150 16110 15202
rect 25218 15150 25230 15202
rect 25282 15150 25294 15202
rect 30818 15150 30830 15202
rect 30882 15150 30894 15202
rect 17502 15138 17554 15150
rect 1598 15090 1650 15102
rect 1598 15026 1650 15038
rect 11790 15090 11842 15102
rect 11790 15026 11842 15038
rect 22094 15090 22146 15102
rect 22094 15026 22146 15038
rect 26350 15090 26402 15102
rect 26350 15026 26402 15038
rect 31502 15090 31554 15102
rect 31502 15026 31554 15038
rect 1344 14922 32592 14956
rect 1344 14870 5120 14922
rect 5172 14870 5224 14922
rect 5276 14870 5328 14922
rect 5380 14870 12932 14922
rect 12984 14870 13036 14922
rect 13088 14870 13140 14922
rect 13192 14870 20744 14922
rect 20796 14870 20848 14922
rect 20900 14870 20952 14922
rect 21004 14870 28556 14922
rect 28608 14870 28660 14922
rect 28712 14870 28764 14922
rect 28816 14870 32592 14922
rect 1344 14836 32592 14870
rect 25678 14754 25730 14766
rect 25678 14690 25730 14702
rect 5182 14642 5234 14654
rect 26126 14642 26178 14654
rect 4050 14590 4062 14642
rect 4114 14590 4126 14642
rect 14802 14590 14814 14642
rect 14866 14590 14878 14642
rect 5182 14578 5234 14590
rect 26126 14578 26178 14590
rect 26462 14642 26514 14654
rect 26898 14590 26910 14642
rect 26962 14590 26974 14642
rect 30146 14590 30158 14642
rect 30210 14590 30222 14642
rect 26462 14578 26514 14590
rect 5518 14530 5570 14542
rect 9214 14530 9266 14542
rect 8530 14478 8542 14530
rect 8594 14478 8606 14530
rect 5518 14466 5570 14478
rect 9214 14466 9266 14478
rect 9550 14530 9602 14542
rect 21982 14530 22034 14542
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 17154 14478 17166 14530
rect 17218 14478 17230 14530
rect 21522 14478 21534 14530
rect 21586 14478 21598 14530
rect 22642 14478 22654 14530
rect 22706 14478 22718 14530
rect 9550 14466 9602 14478
rect 21982 14466 22034 14478
rect 2270 14418 2322 14430
rect 6302 14418 6354 14430
rect 20414 14418 20466 14430
rect 2706 14366 2718 14418
rect 2770 14366 2782 14418
rect 15810 14366 15822 14418
rect 15874 14366 15886 14418
rect 2270 14354 2322 14366
rect 6302 14354 6354 14366
rect 20414 14354 20466 14366
rect 20750 14418 20802 14430
rect 20750 14354 20802 14366
rect 21758 14418 21810 14430
rect 27906 14366 27918 14418
rect 27970 14366 27982 14418
rect 31490 14366 31502 14418
rect 31554 14366 31566 14418
rect 21758 14354 21810 14366
rect 1934 14306 1986 14318
rect 1934 14242 1986 14254
rect 4622 14306 4674 14318
rect 13022 14306 13074 14318
rect 12450 14254 12462 14306
rect 12514 14254 12526 14306
rect 4622 14242 4674 14254
rect 13022 14242 13074 14254
rect 13582 14306 13634 14318
rect 13582 14242 13634 14254
rect 14030 14306 14082 14318
rect 14030 14242 14082 14254
rect 14478 14306 14530 14318
rect 20190 14306 20242 14318
rect 29822 14306 29874 14318
rect 19618 14254 19630 14306
rect 19682 14254 19694 14306
rect 25106 14254 25118 14306
rect 25170 14254 25182 14306
rect 14478 14242 14530 14254
rect 20190 14242 20242 14254
rect 29822 14242 29874 14254
rect 32062 14306 32114 14318
rect 32062 14242 32114 14254
rect 1344 14138 32752 14172
rect 1344 14086 9026 14138
rect 9078 14086 9130 14138
rect 9182 14086 9234 14138
rect 9286 14086 16838 14138
rect 16890 14086 16942 14138
rect 16994 14086 17046 14138
rect 17098 14086 24650 14138
rect 24702 14086 24754 14138
rect 24806 14086 24858 14138
rect 24910 14086 32462 14138
rect 32514 14086 32566 14138
rect 32618 14086 32670 14138
rect 32722 14086 32752 14138
rect 1344 14052 32752 14086
rect 9886 13970 9938 13982
rect 2370 13918 2382 13970
rect 2434 13918 2446 13970
rect 9886 13906 9938 13918
rect 12350 13970 12402 13982
rect 17390 13970 17442 13982
rect 16034 13918 16046 13970
rect 16098 13918 16110 13970
rect 12350 13906 12402 13918
rect 17390 13906 17442 13918
rect 18062 13970 18114 13982
rect 18062 13906 18114 13918
rect 23326 13970 23378 13982
rect 23326 13906 23378 13918
rect 24110 13970 24162 13982
rect 24110 13906 24162 13918
rect 5406 13858 5458 13870
rect 5406 13794 5458 13806
rect 6190 13858 6242 13870
rect 6190 13794 6242 13806
rect 9550 13858 9602 13870
rect 10770 13806 10782 13858
rect 10834 13806 10846 13858
rect 29698 13806 29710 13858
rect 29762 13806 29774 13858
rect 9550 13794 9602 13806
rect 5294 13746 5346 13758
rect 8878 13746 8930 13758
rect 4610 13694 4622 13746
rect 4674 13694 4686 13746
rect 8418 13694 8430 13746
rect 8482 13694 8494 13746
rect 5294 13682 5346 13694
rect 8878 13682 8930 13694
rect 13358 13746 13410 13758
rect 17726 13746 17778 13758
rect 13682 13694 13694 13746
rect 13746 13694 13758 13746
rect 18274 13694 18286 13746
rect 18338 13694 18350 13746
rect 18834 13694 18846 13746
rect 18898 13694 18910 13746
rect 25666 13694 25678 13746
rect 25730 13694 25742 13746
rect 26450 13694 26462 13746
rect 26514 13694 26526 13746
rect 13358 13682 13410 13694
rect 17726 13682 17778 13694
rect 12798 13634 12850 13646
rect 11778 13582 11790 13634
rect 11842 13582 11854 13634
rect 12798 13570 12850 13582
rect 22542 13634 22594 13646
rect 22542 13570 22594 13582
rect 24670 13634 24722 13646
rect 24670 13570 24722 13582
rect 1598 13522 1650 13534
rect 1598 13458 1650 13470
rect 16830 13522 16882 13534
rect 16830 13458 16882 13470
rect 25902 13522 25954 13534
rect 25902 13458 25954 13470
rect 1344 13354 32592 13388
rect 1344 13302 5120 13354
rect 5172 13302 5224 13354
rect 5276 13302 5328 13354
rect 5380 13302 12932 13354
rect 12984 13302 13036 13354
rect 13088 13302 13140 13354
rect 13192 13302 20744 13354
rect 20796 13302 20848 13354
rect 20900 13302 20952 13354
rect 21004 13302 28556 13354
rect 28608 13302 28660 13354
rect 28712 13302 28764 13354
rect 28816 13302 32592 13354
rect 1344 13268 32592 13302
rect 2494 13074 2546 13086
rect 6974 13074 7026 13086
rect 9998 13074 10050 13086
rect 15374 13074 15426 13086
rect 18510 13074 18562 13086
rect 3826 13022 3838 13074
rect 3890 13022 3902 13074
rect 6178 13022 6190 13074
rect 6242 13022 6254 13074
rect 8082 13022 8094 13074
rect 8146 13022 8158 13074
rect 11890 13022 11902 13074
rect 11954 13022 11966 13074
rect 13570 13022 13582 13074
rect 13634 13022 13646 13074
rect 16706 13022 16718 13074
rect 16770 13022 16782 13074
rect 2494 13010 2546 13022
rect 6974 13010 7026 13022
rect 9998 13010 10050 13022
rect 15374 13010 15426 13022
rect 18510 13010 18562 13022
rect 18958 13074 19010 13086
rect 21422 13074 21474 13086
rect 19282 13022 19294 13074
rect 19346 13022 19358 13074
rect 18958 13010 19010 13022
rect 21422 13010 21474 13022
rect 21870 13074 21922 13086
rect 30370 13022 30382 13074
rect 30434 13022 30446 13074
rect 21870 13010 21922 13022
rect 1710 12962 1762 12974
rect 1710 12898 1762 12910
rect 2942 12962 2994 12974
rect 5954 12910 5966 12962
rect 6018 12910 6030 12962
rect 13682 12910 13694 12962
rect 13746 12910 13758 12962
rect 14802 12910 14814 12962
rect 14866 12910 14878 12962
rect 26450 12910 26462 12962
rect 26514 12910 26526 12962
rect 27794 12910 27806 12962
rect 27858 12910 27870 12962
rect 2942 12898 2994 12910
rect 2046 12850 2098 12862
rect 14590 12850 14642 12862
rect 4946 12798 4958 12850
rect 5010 12798 5022 12850
rect 9090 12798 9102 12850
rect 9154 12798 9166 12850
rect 10882 12798 10894 12850
rect 10946 12798 10958 12850
rect 17490 12798 17502 12850
rect 17554 12798 17566 12850
rect 20514 12798 20526 12850
rect 20578 12798 20590 12850
rect 23650 12798 23662 12850
rect 23714 12798 23726 12850
rect 29474 12798 29486 12850
rect 29538 12798 29550 12850
rect 2046 12786 2098 12798
rect 14590 12786 14642 12798
rect 7422 12738 7474 12750
rect 7422 12674 7474 12686
rect 12462 12738 12514 12750
rect 12462 12674 12514 12686
rect 12910 12738 12962 12750
rect 12910 12674 12962 12686
rect 16158 12738 16210 12750
rect 16158 12674 16210 12686
rect 27918 12738 27970 12750
rect 27918 12674 27970 12686
rect 1344 12570 32752 12604
rect 1344 12518 9026 12570
rect 9078 12518 9130 12570
rect 9182 12518 9234 12570
rect 9286 12518 16838 12570
rect 16890 12518 16942 12570
rect 16994 12518 17046 12570
rect 17098 12518 24650 12570
rect 24702 12518 24754 12570
rect 24806 12518 24858 12570
rect 24910 12518 32462 12570
rect 32514 12518 32566 12570
rect 32618 12518 32670 12570
rect 32722 12518 32752 12570
rect 1344 12484 32752 12518
rect 5518 12402 5570 12414
rect 5518 12338 5570 12350
rect 8990 12402 9042 12414
rect 8990 12338 9042 12350
rect 16270 12402 16322 12414
rect 29598 12402 29650 12414
rect 25890 12350 25902 12402
rect 25954 12350 25966 12402
rect 16270 12338 16322 12350
rect 29598 12338 29650 12350
rect 2382 12290 2434 12302
rect 17390 12290 17442 12302
rect 6850 12238 6862 12290
rect 6914 12238 6926 12290
rect 2382 12226 2434 12238
rect 17390 12226 17442 12238
rect 20862 12290 20914 12302
rect 23874 12238 23886 12290
rect 23938 12238 23950 12290
rect 31266 12238 31278 12290
rect 31330 12238 31342 12290
rect 20862 12226 20914 12238
rect 5070 12178 5122 12190
rect 14366 12178 14418 12190
rect 18174 12178 18226 12190
rect 28814 12178 28866 12190
rect 4610 12126 4622 12178
rect 4674 12126 4686 12178
rect 5730 12126 5742 12178
rect 5794 12126 5806 12178
rect 12786 12126 12798 12178
rect 12850 12126 12862 12178
rect 15138 12126 15150 12178
rect 15202 12126 15214 12178
rect 16482 12126 16494 12178
rect 16546 12126 16558 12178
rect 17602 12126 17614 12178
rect 17666 12126 17678 12178
rect 18610 12126 18622 12178
rect 18674 12126 18686 12178
rect 28242 12126 28254 12178
rect 28306 12126 28318 12178
rect 5070 12114 5122 12126
rect 14366 12114 14418 12126
rect 18174 12114 18226 12126
rect 28814 12114 28866 12126
rect 29150 12178 29202 12190
rect 29150 12114 29202 12126
rect 14030 12066 14082 12078
rect 7970 12014 7982 12066
rect 8034 12014 8046 12066
rect 10434 12014 10446 12066
rect 10498 12014 10510 12066
rect 14030 12002 14082 12014
rect 14926 12066 14978 12078
rect 22866 12014 22878 12066
rect 22930 12014 22942 12066
rect 30258 12014 30270 12066
rect 30322 12014 30334 12066
rect 14926 12002 14978 12014
rect 1598 11954 1650 11966
rect 1598 11890 1650 11902
rect 15262 11954 15314 11966
rect 15262 11890 15314 11902
rect 21646 11954 21698 11966
rect 21646 11890 21698 11902
rect 25118 11954 25170 11966
rect 25118 11890 25170 11902
rect 1344 11786 32592 11820
rect 1344 11734 5120 11786
rect 5172 11734 5224 11786
rect 5276 11734 5328 11786
rect 5380 11734 12932 11786
rect 12984 11734 13036 11786
rect 13088 11734 13140 11786
rect 13192 11734 20744 11786
rect 20796 11734 20848 11786
rect 20900 11734 20952 11786
rect 21004 11734 28556 11786
rect 28608 11734 28660 11786
rect 28712 11734 28764 11786
rect 28816 11734 32592 11786
rect 1344 11700 32592 11734
rect 5742 11618 5794 11630
rect 20414 11618 20466 11630
rect 18946 11566 18958 11618
rect 19010 11615 19022 11618
rect 19010 11569 19343 11615
rect 19010 11566 19022 11569
rect 5742 11554 5794 11566
rect 4510 11506 4562 11518
rect 3826 11454 3838 11506
rect 3890 11454 3902 11506
rect 4510 11442 4562 11454
rect 5070 11506 5122 11518
rect 11666 11454 11678 11506
rect 11730 11454 11742 11506
rect 5070 11442 5122 11454
rect 1934 11394 1986 11406
rect 12910 11394 12962 11406
rect 5954 11342 5966 11394
rect 6018 11342 6030 11394
rect 9426 11342 9438 11394
rect 9490 11342 9502 11394
rect 13458 11342 13470 11394
rect 13522 11342 13534 11394
rect 19297 11391 19343 11569
rect 20414 11554 20466 11566
rect 29262 11506 29314 11518
rect 32062 11506 32114 11518
rect 30146 11454 30158 11506
rect 30210 11454 30222 11506
rect 29262 11442 29314 11454
rect 32062 11442 32114 11454
rect 21198 11394 21250 11406
rect 25230 11394 25282 11406
rect 19730 11391 19742 11394
rect 19297 11345 19742 11391
rect 19730 11342 19742 11345
rect 19794 11342 19806 11394
rect 20514 11342 20526 11394
rect 20578 11342 20590 11394
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 25666 11342 25678 11394
rect 25730 11342 25742 11394
rect 1934 11330 1986 11342
rect 12910 11330 12962 11342
rect 21198 11330 21250 11342
rect 25230 11330 25282 11342
rect 2270 11282 2322 11294
rect 27918 11282 27970 11294
rect 3042 11230 3054 11282
rect 3106 11230 3118 11282
rect 15810 11230 15822 11282
rect 15874 11230 15886 11282
rect 31154 11230 31166 11282
rect 31218 11230 31230 11282
rect 2270 11218 2322 11230
rect 27918 11218 27970 11230
rect 6750 11170 6802 11182
rect 6750 11106 6802 11118
rect 7310 11170 7362 11182
rect 7310 11106 7362 11118
rect 19182 11170 19234 11182
rect 24894 11170 24946 11182
rect 24098 11118 24110 11170
rect 24162 11118 24174 11170
rect 19182 11106 19234 11118
rect 24894 11106 24946 11118
rect 28702 11170 28754 11182
rect 28702 11106 28754 11118
rect 1344 11002 32752 11036
rect 1344 10950 9026 11002
rect 9078 10950 9130 11002
rect 9182 10950 9234 11002
rect 9286 10950 16838 11002
rect 16890 10950 16942 11002
rect 16994 10950 17046 11002
rect 17098 10950 24650 11002
rect 24702 10950 24754 11002
rect 24806 10950 24858 11002
rect 24910 10950 32462 11002
rect 32514 10950 32566 11002
rect 32618 10950 32670 11002
rect 32722 10950 32752 11002
rect 1344 10916 32752 10950
rect 9662 10834 9714 10846
rect 4722 10782 4734 10834
rect 4786 10782 4798 10834
rect 6178 10782 6190 10834
rect 6242 10782 6254 10834
rect 9662 10770 9714 10782
rect 10110 10834 10162 10846
rect 10110 10770 10162 10782
rect 10558 10834 10610 10846
rect 10558 10770 10610 10782
rect 22318 10834 22370 10846
rect 22318 10770 22370 10782
rect 30270 10834 30322 10846
rect 30270 10770 30322 10782
rect 16270 10722 16322 10734
rect 25566 10722 25618 10734
rect 20962 10670 20974 10722
rect 21026 10670 21038 10722
rect 23874 10670 23886 10722
rect 23938 10670 23950 10722
rect 16270 10658 16322 10670
rect 25566 10658 25618 10670
rect 29038 10722 29090 10734
rect 29038 10658 29090 10670
rect 30606 10722 30658 10734
rect 30606 10658 30658 10670
rect 32286 10722 32338 10734
rect 32286 10658 32338 10670
rect 9102 10610 9154 10622
rect 19406 10610 19458 10622
rect 1698 10558 1710 10610
rect 1762 10558 1774 10610
rect 2146 10558 2158 10610
rect 2210 10558 2222 10610
rect 8530 10558 8542 10610
rect 8594 10558 8606 10610
rect 10882 10558 10894 10610
rect 10946 10558 10958 10610
rect 15138 10558 15150 10610
rect 15202 10558 15214 10610
rect 16482 10558 16494 10610
rect 16546 10558 16558 10610
rect 18162 10558 18174 10610
rect 18226 10558 18238 10610
rect 9102 10546 9154 10558
rect 19406 10546 19458 10558
rect 25902 10610 25954 10622
rect 25902 10546 25954 10558
rect 26350 10610 26402 10622
rect 30942 10610 30994 10622
rect 26786 10558 26798 10610
rect 26850 10558 26862 10610
rect 26350 10546 26402 10558
rect 30942 10546 30994 10558
rect 18958 10498 19010 10510
rect 21870 10498 21922 10510
rect 15250 10446 15262 10498
rect 15314 10446 15326 10498
rect 19954 10446 19966 10498
rect 20018 10446 20030 10498
rect 22866 10446 22878 10498
rect 22930 10446 22942 10498
rect 18958 10434 19010 10446
rect 21870 10434 21922 10446
rect 5294 10386 5346 10398
rect 5294 10322 5346 10334
rect 5406 10386 5458 10398
rect 13694 10386 13746 10398
rect 9650 10334 9662 10386
rect 9714 10383 9726 10386
rect 10658 10383 10670 10386
rect 9714 10337 10670 10383
rect 9714 10334 9726 10337
rect 10658 10334 10670 10337
rect 10722 10334 10734 10386
rect 5406 10322 5458 10334
rect 13694 10322 13746 10334
rect 18062 10386 18114 10398
rect 18062 10322 18114 10334
rect 29822 10386 29874 10398
rect 29822 10322 29874 10334
rect 31726 10386 31778 10398
rect 31726 10322 31778 10334
rect 1344 10218 32592 10252
rect 1344 10166 5120 10218
rect 5172 10166 5224 10218
rect 5276 10166 5328 10218
rect 5380 10166 12932 10218
rect 12984 10166 13036 10218
rect 13088 10166 13140 10218
rect 13192 10166 20744 10218
rect 20796 10166 20848 10218
rect 20900 10166 20952 10218
rect 21004 10166 28556 10218
rect 28608 10166 28660 10218
rect 28712 10166 28764 10218
rect 28816 10166 32592 10218
rect 1344 10132 32592 10166
rect 18958 10050 19010 10062
rect 18958 9986 19010 9998
rect 23102 10050 23154 10062
rect 23102 9986 23154 9998
rect 4622 9938 4674 9950
rect 29822 9938 29874 9950
rect 32174 9938 32226 9950
rect 3938 9886 3950 9938
rect 4002 9886 4014 9938
rect 9090 9886 9102 9938
rect 9154 9886 9166 9938
rect 30146 9886 30158 9938
rect 30210 9886 30222 9938
rect 4622 9874 4674 9886
rect 29822 9874 29874 9886
rect 32174 9874 32226 9886
rect 15262 9826 15314 9838
rect 23662 9826 23714 9838
rect 2034 9774 2046 9826
rect 2098 9774 2110 9826
rect 6626 9774 6638 9826
rect 6690 9774 6702 9826
rect 8306 9774 8318 9826
rect 8370 9774 8382 9826
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 14802 9774 14814 9826
rect 14866 9774 14878 9826
rect 15922 9774 15934 9826
rect 15986 9774 15998 9826
rect 19394 9774 19406 9826
rect 19458 9774 19470 9826
rect 20738 9774 20750 9826
rect 20802 9774 20814 9826
rect 21522 9774 21534 9826
rect 21586 9774 21598 9826
rect 22978 9774 22990 9826
rect 23042 9774 23054 9826
rect 23986 9774 23998 9826
rect 24050 9774 24062 9826
rect 27346 9774 27358 9826
rect 27410 9774 27422 9826
rect 15262 9762 15314 9774
rect 23662 9762 23714 9774
rect 2270 9714 2322 9726
rect 18174 9714 18226 9726
rect 3042 9662 3054 9714
rect 3106 9662 3118 9714
rect 31154 9662 31166 9714
rect 31218 9662 31230 9714
rect 2270 9650 2322 9662
rect 18174 9650 18226 9662
rect 5070 9602 5122 9614
rect 5070 9538 5122 9550
rect 6638 9602 6690 9614
rect 6638 9538 6690 9550
rect 12686 9602 12738 9614
rect 12686 9538 12738 9550
rect 13582 9602 13634 9614
rect 13582 9538 13634 9550
rect 14590 9602 14642 9614
rect 14590 9538 14642 9550
rect 19182 9602 19234 9614
rect 19182 9538 19234 9550
rect 20638 9602 20690 9614
rect 20638 9538 20690 9550
rect 21422 9602 21474 9614
rect 27134 9602 27186 9614
rect 26450 9550 26462 9602
rect 26514 9550 26526 9602
rect 21422 9538 21474 9550
rect 27134 9538 27186 9550
rect 27470 9602 27522 9614
rect 27470 9538 27522 9550
rect 28590 9602 28642 9614
rect 28590 9538 28642 9550
rect 1344 9434 32752 9468
rect 1344 9382 9026 9434
rect 9078 9382 9130 9434
rect 9182 9382 9234 9434
rect 9286 9382 16838 9434
rect 16890 9382 16942 9434
rect 16994 9382 17046 9434
rect 17098 9382 24650 9434
rect 24702 9382 24754 9434
rect 24806 9382 24858 9434
rect 24910 9382 32462 9434
rect 32514 9382 32566 9434
rect 32618 9382 32670 9434
rect 32722 9382 32752 9434
rect 1344 9348 32752 9382
rect 10446 9266 10498 9278
rect 4498 9214 4510 9266
rect 4562 9214 4574 9266
rect 8306 9214 8318 9266
rect 8370 9214 8382 9266
rect 10446 9202 10498 9214
rect 10894 9266 10946 9278
rect 10894 9202 10946 9214
rect 11230 9266 11282 9278
rect 22318 9266 22370 9278
rect 21186 9214 21198 9266
rect 21250 9214 21262 9266
rect 11230 9202 11282 9214
rect 22318 9202 22370 9214
rect 22878 9266 22930 9278
rect 22878 9202 22930 9214
rect 26462 9266 26514 9278
rect 26462 9202 26514 9214
rect 27582 9266 27634 9278
rect 31502 9266 31554 9278
rect 30818 9214 30830 9266
rect 30882 9214 30894 9266
rect 27582 9202 27634 9214
rect 31502 9202 31554 9214
rect 31726 9266 31778 9278
rect 31726 9202 31778 9214
rect 9550 9154 9602 9166
rect 16158 9154 16210 9166
rect 12786 9102 12798 9154
rect 12850 9102 12862 9154
rect 9550 9090 9602 9102
rect 16158 9090 16210 9102
rect 17390 9154 17442 9166
rect 17390 9090 17442 9102
rect 17726 9154 17778 9166
rect 32062 9154 32114 9166
rect 24210 9102 24222 9154
rect 24274 9102 24286 9154
rect 17726 9090 17778 9102
rect 32062 9090 32114 9102
rect 1822 9042 1874 9054
rect 5406 9042 5458 9054
rect 13246 9042 13298 9054
rect 18286 9042 18338 9054
rect 28030 9042 28082 9054
rect 2258 8990 2270 9042
rect 2322 8990 2334 9042
rect 6066 8990 6078 9042
rect 6130 8990 6142 9042
rect 9762 8990 9774 9042
rect 9826 8990 9838 9042
rect 13906 8990 13918 9042
rect 13970 8990 13982 9042
rect 18946 8990 18958 9042
rect 19010 8990 19022 9042
rect 25218 8990 25230 9042
rect 25282 8990 25294 9042
rect 26338 8990 26350 9042
rect 26402 8990 26414 9042
rect 28354 8990 28366 9042
rect 28418 8990 28430 9042
rect 1822 8978 1874 8990
rect 5406 8978 5458 8990
rect 13246 8978 13298 8990
rect 18286 8978 18338 8990
rect 28030 8978 28082 8990
rect 11666 8878 11678 8930
rect 11730 8878 11742 8930
rect 23202 8878 23214 8930
rect 23266 8878 23278 8930
rect 5294 8818 5346 8830
rect 5294 8754 5346 8766
rect 9102 8818 9154 8830
rect 9102 8754 9154 8766
rect 16942 8818 16994 8830
rect 16942 8754 16994 8766
rect 21982 8818 22034 8830
rect 21982 8754 22034 8766
rect 25342 8818 25394 8830
rect 25342 8754 25394 8766
rect 1344 8650 32592 8684
rect 1344 8598 5120 8650
rect 5172 8598 5224 8650
rect 5276 8598 5328 8650
rect 5380 8598 12932 8650
rect 12984 8598 13036 8650
rect 13088 8598 13140 8650
rect 13192 8598 20744 8650
rect 20796 8598 20848 8650
rect 20900 8598 20952 8650
rect 21004 8598 28556 8650
rect 28608 8598 28660 8650
rect 28712 8598 28764 8650
rect 28816 8598 32592 8650
rect 1344 8564 32592 8598
rect 13022 8482 13074 8494
rect 13022 8418 13074 8430
rect 5070 8370 5122 8382
rect 19294 8370 19346 8382
rect 4050 8318 4062 8370
rect 4114 8318 4126 8370
rect 14802 8318 14814 8370
rect 14866 8318 14878 8370
rect 5070 8306 5122 8318
rect 19294 8306 19346 8318
rect 29710 8370 29762 8382
rect 30258 8318 30270 8370
rect 30322 8318 30334 8370
rect 29710 8306 29762 8318
rect 5518 8258 5570 8270
rect 15822 8258 15874 8270
rect 21198 8258 21250 8270
rect 24894 8258 24946 8270
rect 28702 8258 28754 8270
rect 6066 8206 6078 8258
rect 6130 8206 6142 8258
rect 9426 8206 9438 8258
rect 9490 8206 9502 8258
rect 9874 8206 9886 8258
rect 9938 8206 9950 8258
rect 14242 8206 14254 8258
rect 14306 8206 14318 8258
rect 15026 8206 15038 8258
rect 15090 8206 15102 8258
rect 16258 8206 16270 8258
rect 16322 8206 16334 8258
rect 19506 8206 19518 8258
rect 19570 8206 19582 8258
rect 21858 8206 21870 8258
rect 21922 8206 21934 8258
rect 28130 8206 28142 8258
rect 28194 8206 28206 8258
rect 5518 8194 5570 8206
rect 15822 8194 15874 8206
rect 21198 8194 21250 8206
rect 24894 8194 24946 8206
rect 28702 8194 28754 8206
rect 1934 8146 1986 8158
rect 1934 8082 1986 8094
rect 2270 8146 2322 8158
rect 25790 8146 25842 8158
rect 2706 8094 2718 8146
rect 2770 8094 2782 8146
rect 31154 8094 31166 8146
rect 31218 8094 31230 8146
rect 2270 8082 2322 8094
rect 25790 8082 25842 8094
rect 9214 8034 9266 8046
rect 14142 8034 14194 8046
rect 19630 8034 19682 8046
rect 8642 7982 8654 8034
rect 8706 7982 8718 8034
rect 12450 7982 12462 8034
rect 12514 7982 12526 8034
rect 18722 7982 18734 8034
rect 18786 7982 18798 8034
rect 9214 7970 9266 7982
rect 14142 7970 14194 7982
rect 19630 7970 19682 7982
rect 20750 8034 20802 8046
rect 25006 8034 25058 8046
rect 24322 7982 24334 8034
rect 24386 7982 24398 8034
rect 20750 7970 20802 7982
rect 25006 7970 25058 7982
rect 29262 8034 29314 8046
rect 29262 7970 29314 7982
rect 32062 8034 32114 8046
rect 32062 7970 32114 7982
rect 1344 7866 32752 7900
rect 1344 7814 9026 7866
rect 9078 7814 9130 7866
rect 9182 7814 9234 7866
rect 9286 7814 16838 7866
rect 16890 7814 16942 7866
rect 16994 7814 17046 7866
rect 17098 7814 24650 7866
rect 24702 7814 24754 7866
rect 24806 7814 24858 7866
rect 24910 7814 32462 7866
rect 32514 7814 32566 7866
rect 32618 7814 32670 7866
rect 32722 7814 32752 7866
rect 1344 7780 32752 7814
rect 1822 7698 1874 7710
rect 8654 7698 8706 7710
rect 7410 7646 7422 7698
rect 7474 7646 7486 7698
rect 1822 7634 1874 7646
rect 8654 7634 8706 7646
rect 9662 7698 9714 7710
rect 9662 7634 9714 7646
rect 10782 7698 10834 7710
rect 15262 7698 15314 7710
rect 14130 7646 14142 7698
rect 14194 7646 14206 7698
rect 10782 7634 10834 7646
rect 15262 7634 15314 7646
rect 16830 7698 16882 7710
rect 16830 7634 16882 7646
rect 17950 7698 18002 7710
rect 17950 7634 18002 7646
rect 24670 7698 24722 7710
rect 31154 7646 31166 7698
rect 31218 7646 31230 7698
rect 24670 7634 24722 7646
rect 20862 7586 20914 7598
rect 3938 7534 3950 7586
rect 4002 7534 4014 7586
rect 19394 7534 19406 7586
rect 19458 7534 19470 7586
rect 27570 7534 27582 7586
rect 27634 7534 27646 7586
rect 20862 7522 20914 7534
rect 4622 7474 4674 7486
rect 11118 7474 11170 7486
rect 23550 7474 23602 7486
rect 5058 7422 5070 7474
rect 5122 7422 5134 7474
rect 8418 7422 8430 7474
rect 8482 7422 8494 7474
rect 11666 7422 11678 7474
rect 11730 7422 11742 7474
rect 16034 7422 16046 7474
rect 16098 7422 16110 7474
rect 23202 7422 23214 7474
rect 23266 7422 23278 7474
rect 4622 7410 4674 7422
rect 11118 7410 11170 7422
rect 23550 7410 23602 7422
rect 24334 7474 24386 7486
rect 24334 7410 24386 7422
rect 28478 7474 28530 7486
rect 28914 7422 28926 7474
rect 28978 7422 28990 7474
rect 28478 7410 28530 7422
rect 17502 7362 17554 7374
rect 2706 7310 2718 7362
rect 2770 7310 2782 7362
rect 10098 7310 10110 7362
rect 10162 7310 10174 7362
rect 16146 7310 16158 7362
rect 16210 7310 16222 7362
rect 18386 7310 18398 7362
rect 18450 7310 18462 7362
rect 26226 7310 26238 7362
rect 26290 7310 26302 7362
rect 17502 7298 17554 7310
rect 8094 7250 8146 7262
rect 8094 7186 8146 7198
rect 14814 7250 14866 7262
rect 14814 7186 14866 7198
rect 20078 7250 20130 7262
rect 20078 7186 20130 7198
rect 31950 7250 32002 7262
rect 31950 7186 32002 7198
rect 1344 7082 32592 7116
rect 1344 7030 5120 7082
rect 5172 7030 5224 7082
rect 5276 7030 5328 7082
rect 5380 7030 12932 7082
rect 12984 7030 13036 7082
rect 13088 7030 13140 7082
rect 13192 7030 20744 7082
rect 20796 7030 20848 7082
rect 20900 7030 20952 7082
rect 21004 7030 28556 7082
rect 28608 7030 28660 7082
rect 28712 7030 28764 7082
rect 28816 7030 32592 7082
rect 1344 6996 32592 7030
rect 5070 6802 5122 6814
rect 14254 6802 14306 6814
rect 4050 6750 4062 6802
rect 4114 6750 4126 6802
rect 11218 6750 11230 6802
rect 11282 6750 11294 6802
rect 15474 6750 15486 6802
rect 15538 6750 15550 6802
rect 19170 6750 19182 6802
rect 19234 6750 19246 6802
rect 23090 6750 23102 6802
rect 23154 6750 23166 6802
rect 25890 6750 25902 6802
rect 25954 6750 25966 6802
rect 30146 6750 30158 6802
rect 30210 6750 30222 6802
rect 5070 6738 5122 6750
rect 14254 6738 14306 6750
rect 6302 6690 6354 6702
rect 10334 6690 10386 6702
rect 1810 6638 1822 6690
rect 1874 6638 1886 6690
rect 6850 6638 6862 6690
rect 6914 6638 6926 6690
rect 6302 6626 6354 6638
rect 10334 6626 10386 6638
rect 10782 6690 10834 6702
rect 10782 6626 10834 6638
rect 18846 6690 18898 6702
rect 21522 6638 21534 6690
rect 21586 6638 21598 6690
rect 28242 6638 28254 6690
rect 28306 6638 28318 6690
rect 18846 6626 18898 6638
rect 2046 6578 2098 6590
rect 5630 6578 5682 6590
rect 3042 6526 3054 6578
rect 3106 6526 3118 6578
rect 2046 6514 2098 6526
rect 5630 6514 5682 6526
rect 5966 6578 6018 6590
rect 13470 6578 13522 6590
rect 12226 6526 12238 6578
rect 12290 6526 12302 6578
rect 5966 6514 6018 6526
rect 13470 6514 13522 6526
rect 13806 6578 13858 6590
rect 13806 6514 13858 6526
rect 14702 6578 14754 6590
rect 17502 6578 17554 6590
rect 16706 6526 16718 6578
rect 16770 6526 16782 6578
rect 20178 6526 20190 6578
rect 20242 6526 20254 6578
rect 24098 6526 24110 6578
rect 24162 6526 24174 6578
rect 26898 6526 26910 6578
rect 26962 6526 26974 6578
rect 28466 6526 28478 6578
rect 28530 6526 28542 6578
rect 31490 6526 31502 6578
rect 31554 6526 31566 6578
rect 14702 6514 14754 6526
rect 17502 6514 17554 6526
rect 4510 6466 4562 6478
rect 9998 6466 10050 6478
rect 9426 6414 9438 6466
rect 9490 6414 9502 6466
rect 4510 6402 4562 6414
rect 9998 6402 10050 6414
rect 15150 6466 15202 6478
rect 15150 6402 15202 6414
rect 17838 6466 17890 6478
rect 17838 6402 17890 6414
rect 18286 6466 18338 6478
rect 18286 6402 18338 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 22318 6466 22370 6478
rect 22318 6402 22370 6414
rect 32062 6466 32114 6478
rect 32062 6402 32114 6414
rect 1344 6298 32752 6332
rect 1344 6246 9026 6298
rect 9078 6246 9130 6298
rect 9182 6246 9234 6298
rect 9286 6246 16838 6298
rect 16890 6246 16942 6298
rect 16994 6246 17046 6298
rect 17098 6246 24650 6298
rect 24702 6246 24754 6298
rect 24806 6246 24858 6298
rect 24910 6246 32462 6298
rect 32514 6246 32566 6298
rect 32618 6246 32670 6298
rect 32722 6246 32752 6298
rect 1344 6212 32752 6246
rect 3614 6130 3666 6142
rect 3614 6066 3666 6078
rect 4062 6130 4114 6142
rect 4062 6066 4114 6078
rect 8094 6130 8146 6142
rect 8094 6066 8146 6078
rect 9550 6130 9602 6142
rect 9550 6066 9602 6078
rect 14926 6130 14978 6142
rect 14926 6066 14978 6078
rect 27582 6130 27634 6142
rect 27582 6066 27634 6078
rect 28366 6130 28418 6142
rect 29138 6078 29150 6130
rect 29202 6078 29214 6130
rect 28366 6066 28418 6078
rect 4846 6018 4898 6030
rect 4846 5954 4898 5966
rect 13358 6018 13410 6030
rect 13358 5954 13410 5966
rect 14478 6018 14530 6030
rect 20190 6018 20242 6030
rect 16370 5966 16382 6018
rect 16434 5966 16446 6018
rect 14478 5954 14530 5966
rect 20190 5954 20242 5966
rect 20974 6018 21026 6030
rect 20974 5954 21026 5966
rect 21870 6018 21922 6030
rect 25342 6018 25394 6030
rect 22306 5966 22318 6018
rect 22370 5966 22382 6018
rect 25778 5966 25790 6018
rect 25842 5966 25854 6018
rect 21870 5954 21922 5966
rect 25342 5954 25394 5966
rect 7534 5906 7586 5918
rect 10670 5906 10722 5918
rect 17502 5906 17554 5918
rect 32062 5906 32114 5918
rect 2930 5854 2942 5906
rect 2994 5854 3006 5906
rect 3378 5854 3390 5906
rect 3442 5854 3454 5906
rect 7186 5854 7198 5906
rect 7250 5854 7262 5906
rect 8082 5854 8094 5906
rect 8146 5854 8158 5906
rect 9762 5854 9774 5906
rect 9826 5854 9838 5906
rect 11106 5854 11118 5906
rect 11170 5854 11182 5906
rect 17826 5854 17838 5906
rect 17890 5854 17902 5906
rect 21634 5854 21646 5906
rect 21698 5854 21710 5906
rect 31378 5854 31390 5906
rect 31442 5854 31454 5906
rect 7534 5842 7586 5854
rect 10670 5842 10722 5854
rect 17502 5842 17554 5854
rect 32062 5842 32114 5854
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 15362 5742 15374 5794
rect 15426 5742 15438 5794
rect 23426 5742 23438 5794
rect 23490 5742 23502 5794
rect 27122 5742 27134 5794
rect 27186 5742 27198 5794
rect 14142 5682 14194 5694
rect 14142 5618 14194 5630
rect 1344 5514 32592 5548
rect 1344 5462 5120 5514
rect 5172 5462 5224 5514
rect 5276 5462 5328 5514
rect 5380 5462 12932 5514
rect 12984 5462 13036 5514
rect 13088 5462 13140 5514
rect 13192 5462 20744 5514
rect 20796 5462 20848 5514
rect 20900 5462 20952 5514
rect 21004 5462 28556 5514
rect 28608 5462 28660 5514
rect 28712 5462 28764 5514
rect 28816 5462 32592 5514
rect 1344 5428 32592 5462
rect 12798 5346 12850 5358
rect 12798 5282 12850 5294
rect 18174 5346 18226 5358
rect 18174 5282 18226 5294
rect 19742 5346 19794 5358
rect 19742 5282 19794 5294
rect 21982 5346 22034 5358
rect 21982 5282 22034 5294
rect 23774 5346 23826 5358
rect 23774 5282 23826 5294
rect 3950 5234 4002 5246
rect 2146 5182 2158 5234
rect 2210 5182 2222 5234
rect 3950 5170 4002 5182
rect 4734 5234 4786 5246
rect 4734 5170 4786 5182
rect 6974 5234 7026 5246
rect 6974 5170 7026 5182
rect 24334 5234 24386 5246
rect 29822 5234 29874 5246
rect 32062 5234 32114 5246
rect 25330 5182 25342 5234
rect 25394 5182 25406 5234
rect 27570 5182 27582 5234
rect 27634 5182 27646 5234
rect 30146 5182 30158 5234
rect 30210 5182 30222 5234
rect 24334 5170 24386 5182
rect 29822 5170 29874 5182
rect 32062 5170 32114 5182
rect 11678 5122 11730 5134
rect 14702 5122 14754 5134
rect 20414 5122 20466 5134
rect 24670 5122 24722 5134
rect 6402 5070 6414 5122
rect 6466 5070 6478 5122
rect 11218 5070 11230 5122
rect 11282 5070 11294 5122
rect 12562 5070 12574 5122
rect 12626 5070 12638 5122
rect 13906 5070 13918 5122
rect 13970 5070 13982 5122
rect 15138 5070 15150 5122
rect 15202 5070 15214 5122
rect 18498 5070 18510 5122
rect 18562 5070 18574 5122
rect 19842 5070 19854 5122
rect 19906 5070 19918 5122
rect 22082 5070 22094 5122
rect 22146 5070 22158 5122
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 11678 5058 11730 5070
rect 14702 5058 14754 5070
rect 20414 5058 20466 5070
rect 24670 5058 24722 5070
rect 17390 5010 17442 5022
rect 3266 4958 3278 5010
rect 3330 4958 3342 5010
rect 6290 4958 6302 5010
rect 6354 4958 6366 5010
rect 17390 4946 17442 4958
rect 18734 5010 18786 5022
rect 26562 4958 26574 5010
rect 26626 4958 26638 5010
rect 31154 4958 31166 5010
rect 31218 4958 31230 5010
rect 18734 4946 18786 4958
rect 5070 4898 5122 4910
rect 5070 4834 5122 4846
rect 7198 4898 7250 4910
rect 7198 4834 7250 4846
rect 7982 4898 8034 4910
rect 7982 4834 8034 4846
rect 8206 4898 8258 4910
rect 14142 4898 14194 4910
rect 8754 4846 8766 4898
rect 8818 4846 8830 4898
rect 8206 4834 8258 4846
rect 14142 4834 14194 4846
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 21422 4898 21474 4910
rect 21422 4834 21474 4846
rect 25790 4898 25842 4910
rect 25790 4834 25842 4846
rect 1344 4730 32752 4764
rect 1344 4678 9026 4730
rect 9078 4678 9130 4730
rect 9182 4678 9234 4730
rect 9286 4678 16838 4730
rect 16890 4678 16942 4730
rect 16994 4678 17046 4730
rect 17098 4678 24650 4730
rect 24702 4678 24754 4730
rect 24806 4678 24858 4730
rect 24910 4678 32462 4730
rect 32514 4678 32566 4730
rect 32618 4678 32670 4730
rect 32722 4678 32752 4730
rect 1344 4644 32752 4678
rect 5518 4562 5570 4574
rect 5518 4498 5570 4510
rect 8430 4562 8482 4574
rect 8430 4498 8482 4510
rect 8990 4562 9042 4574
rect 8990 4498 9042 4510
rect 11902 4562 11954 4574
rect 11902 4498 11954 4510
rect 12350 4562 12402 4574
rect 17726 4562 17778 4574
rect 15474 4510 15486 4562
rect 15538 4510 15550 4562
rect 12350 4498 12402 4510
rect 17726 4498 17778 4510
rect 18062 4562 18114 4574
rect 18062 4498 18114 4510
rect 20302 4562 20354 4574
rect 20302 4498 20354 4510
rect 21422 4562 21474 4574
rect 21422 4498 21474 4510
rect 23102 4562 23154 4574
rect 23102 4498 23154 4510
rect 26014 4562 26066 4574
rect 26014 4498 26066 4510
rect 26798 4562 26850 4574
rect 26798 4498 26850 4510
rect 28142 4562 28194 4574
rect 28690 4510 28702 4562
rect 28754 4510 28766 4562
rect 28142 4498 28194 4510
rect 2382 4450 2434 4462
rect 16270 4450 16322 4462
rect 7746 4398 7758 4450
rect 7810 4398 7822 4450
rect 10098 4398 10110 4450
rect 10162 4398 10174 4450
rect 2382 4386 2434 4398
rect 16270 4386 16322 4398
rect 16830 4450 16882 4462
rect 22766 4450 22818 4462
rect 19394 4398 19406 4450
rect 19458 4398 19470 4450
rect 16830 4386 16882 4398
rect 22766 4386 22818 4398
rect 25566 4450 25618 4462
rect 25566 4386 25618 4398
rect 32174 4450 32226 4462
rect 32174 4386 32226 4398
rect 5294 4338 5346 4350
rect 4722 4286 4734 4338
rect 4786 4286 4798 4338
rect 5294 4274 5346 4286
rect 5854 4338 5906 4350
rect 5854 4274 5906 4286
rect 12798 4338 12850 4350
rect 25230 4338 25282 4350
rect 27918 4338 27970 4350
rect 31614 4338 31666 4350
rect 13234 4286 13246 4338
rect 13298 4286 13310 4338
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 20178 4286 20190 4338
rect 20242 4286 20254 4338
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 23538 4286 23550 4338
rect 23602 4286 23614 4338
rect 26226 4286 26238 4338
rect 26290 4286 26302 4338
rect 31154 4286 31166 4338
rect 31218 4286 31230 4338
rect 12798 4274 12850 4286
rect 25230 4274 25282 4286
rect 27918 4274 27970 4286
rect 31614 4274 31666 4286
rect 24670 4226 24722 4238
rect 6514 4174 6526 4226
rect 6578 4174 6590 4226
rect 11106 4174 11118 4226
rect 11170 4174 11182 4226
rect 18386 4174 18398 4226
rect 18450 4174 18462 4226
rect 27346 4174 27358 4226
rect 27410 4174 27422 4226
rect 24670 4162 24722 4174
rect 1598 4114 1650 4126
rect 1598 4050 1650 4062
rect 24222 4114 24274 4126
rect 24222 4050 24274 4062
rect 1344 3946 32592 3980
rect 1344 3894 5120 3946
rect 5172 3894 5224 3946
rect 5276 3894 5328 3946
rect 5380 3894 12932 3946
rect 12984 3894 13036 3946
rect 13088 3894 13140 3946
rect 13192 3894 20744 3946
rect 20796 3894 20848 3946
rect 20900 3894 20952 3946
rect 21004 3894 28556 3946
rect 28608 3894 28660 3946
rect 28712 3894 28764 3946
rect 28816 3894 32592 3946
rect 1344 3860 32592 3894
rect 20862 3778 20914 3790
rect 20862 3714 20914 3726
rect 27694 3778 27746 3790
rect 27694 3714 27746 3726
rect 4622 3666 4674 3678
rect 3826 3614 3838 3666
rect 3890 3614 3902 3666
rect 4622 3602 4674 3614
rect 5070 3666 5122 3678
rect 5070 3602 5122 3614
rect 5742 3666 5794 3678
rect 5742 3602 5794 3614
rect 6302 3666 6354 3678
rect 14030 3666 14082 3678
rect 6626 3614 6638 3666
rect 6690 3614 6702 3666
rect 10994 3614 11006 3666
rect 11058 3614 11070 3666
rect 6302 3602 6354 3614
rect 14030 3602 14082 3614
rect 14590 3666 14642 3678
rect 17166 3666 17218 3678
rect 14802 3614 14814 3666
rect 14866 3614 14878 3666
rect 14590 3602 14642 3614
rect 17166 3602 17218 3614
rect 17726 3666 17778 3678
rect 24110 3666 24162 3678
rect 29934 3666 29986 3678
rect 18162 3614 18174 3666
rect 18226 3614 18238 3666
rect 23426 3614 23438 3666
rect 23490 3614 23502 3666
rect 26002 3614 26014 3666
rect 26066 3614 26078 3666
rect 30146 3614 30158 3666
rect 30210 3614 30222 3666
rect 17726 3602 17778 3614
rect 24110 3602 24162 3614
rect 29934 3602 29986 3614
rect 12126 3554 12178 3566
rect 19854 3554 19906 3566
rect 22766 3554 22818 3566
rect 1810 3502 1822 3554
rect 1874 3502 1886 3554
rect 13346 3502 13358 3554
rect 13410 3502 13422 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 22194 3502 22206 3554
rect 22258 3502 22270 3554
rect 12126 3490 12178 3502
rect 19854 3490 19906 3502
rect 22766 3490 22818 3502
rect 25118 3554 25170 3566
rect 25118 3490 25170 3502
rect 25566 3554 25618 3566
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 25566 3490 25618 3502
rect 2046 3442 2098 3454
rect 8318 3442 8370 3454
rect 2594 3390 2606 3442
rect 2658 3390 2670 3442
rect 7522 3390 7534 3442
rect 7586 3390 7598 3442
rect 2046 3378 2098 3390
rect 8318 3378 8370 3390
rect 8654 3442 8706 3454
rect 13134 3442 13186 3454
rect 20190 3442 20242 3454
rect 9986 3390 9998 3442
rect 10050 3390 10062 3442
rect 15810 3390 15822 3442
rect 15874 3390 15886 3442
rect 18946 3390 18958 3442
rect 19010 3390 19022 3442
rect 8654 3378 8706 3390
rect 13134 3378 13186 3390
rect 20190 3378 20242 3390
rect 22430 3442 22482 3454
rect 22430 3378 22482 3390
rect 28366 3442 28418 3454
rect 31154 3390 31166 3442
rect 31218 3390 31230 3442
rect 28366 3378 28418 3390
rect 12350 3330 12402 3342
rect 12350 3266 12402 3278
rect 24558 3330 24610 3342
rect 24558 3266 24610 3278
rect 1344 3162 32752 3196
rect 1344 3110 9026 3162
rect 9078 3110 9130 3162
rect 9182 3110 9234 3162
rect 9286 3110 16838 3162
rect 16890 3110 16942 3162
rect 16994 3110 17046 3162
rect 17098 3110 24650 3162
rect 24702 3110 24754 3162
rect 24806 3110 24858 3162
rect 24910 3110 32462 3162
rect 32514 3110 32566 3162
rect 32618 3110 32670 3162
rect 32722 3110 32752 3162
rect 1344 3076 32752 3110
<< via1 >>
rect 29262 30718 29314 30770
rect 30158 30718 30210 30770
rect 5120 30550 5172 30602
rect 5224 30550 5276 30602
rect 5328 30550 5380 30602
rect 12932 30550 12984 30602
rect 13036 30550 13088 30602
rect 13140 30550 13192 30602
rect 20744 30550 20796 30602
rect 20848 30550 20900 30602
rect 20952 30550 21004 30602
rect 28556 30550 28608 30602
rect 28660 30550 28712 30602
rect 28764 30550 28816 30602
rect 7422 30270 7474 30322
rect 11566 30270 11618 30322
rect 14926 30270 14978 30322
rect 17950 30270 18002 30322
rect 21758 30270 21810 30322
rect 30158 30270 30210 30322
rect 2158 30158 2210 30210
rect 13582 30158 13634 30210
rect 14030 30158 14082 30210
rect 19966 30158 20018 30210
rect 21422 30158 21474 30210
rect 25230 30158 25282 30210
rect 26910 30158 26962 30210
rect 3390 30046 3442 30098
rect 4958 30046 5010 30098
rect 5630 30046 5682 30098
rect 5966 30046 6018 30098
rect 8654 30046 8706 30098
rect 9438 30046 9490 30098
rect 9774 30046 9826 30098
rect 10558 30046 10610 30098
rect 12014 30046 12066 30098
rect 13246 30046 13298 30098
rect 16270 30046 16322 30098
rect 19182 30046 19234 30098
rect 22766 30046 22818 30098
rect 23550 30046 23602 30098
rect 23886 30046 23938 30098
rect 24782 30046 24834 30098
rect 26686 30046 26738 30098
rect 27358 30046 27410 30098
rect 28478 30046 28530 30098
rect 28814 30046 28866 30098
rect 31278 30046 31330 30098
rect 1934 29934 1986 29986
rect 2942 29934 2994 29986
rect 3838 29934 3890 29986
rect 4174 29934 4226 29986
rect 6414 29934 6466 29986
rect 6974 29934 7026 29986
rect 19742 29934 19794 29986
rect 21086 29934 21138 29986
rect 25902 29934 25954 29986
rect 27470 29934 27522 29986
rect 9026 29766 9078 29818
rect 9130 29766 9182 29818
rect 9234 29766 9286 29818
rect 16838 29766 16890 29818
rect 16942 29766 16994 29818
rect 17046 29766 17098 29818
rect 24650 29766 24702 29818
rect 24754 29766 24806 29818
rect 24858 29766 24910 29818
rect 32462 29766 32514 29818
rect 32566 29766 32618 29818
rect 32670 29766 32722 29818
rect 1822 29598 1874 29650
rect 9550 29598 9602 29650
rect 10782 29598 10834 29650
rect 19070 29598 19122 29650
rect 19406 29598 19458 29650
rect 20190 29598 20242 29650
rect 23998 29598 24050 29650
rect 28142 29598 28194 29650
rect 5182 29486 5234 29538
rect 8990 29486 9042 29538
rect 12014 29486 12066 29538
rect 16606 29486 16658 29538
rect 27246 29486 27298 29538
rect 30270 29486 30322 29538
rect 2606 29374 2658 29426
rect 2942 29374 2994 29426
rect 7422 29374 7474 29426
rect 8094 29374 8146 29426
rect 8766 29374 8818 29426
rect 10110 29374 10162 29426
rect 17502 29374 17554 29426
rect 22542 29374 22594 29426
rect 23102 29374 23154 29426
rect 24334 29374 24386 29426
rect 25342 29374 25394 29426
rect 30942 29374 30994 29426
rect 3614 29262 3666 29314
rect 4174 29262 4226 29314
rect 11342 29262 11394 29314
rect 13022 29262 13074 29314
rect 15374 29262 15426 29314
rect 17838 29262 17890 29314
rect 26238 29262 26290 29314
rect 29038 29262 29090 29314
rect 32174 29262 32226 29314
rect 4398 29150 4450 29202
rect 31726 29150 31778 29202
rect 5120 28982 5172 29034
rect 5224 28982 5276 29034
rect 5328 28982 5380 29034
rect 12932 28982 12984 29034
rect 13036 28982 13088 29034
rect 13140 28982 13192 29034
rect 20744 28982 20796 29034
rect 20848 28982 20900 29034
rect 20952 28982 21004 29034
rect 28556 28982 28608 29034
rect 28660 28982 28712 29034
rect 28764 28982 28816 29034
rect 9326 28814 9378 28866
rect 9998 28814 10050 28866
rect 17054 28814 17106 28866
rect 20862 28814 20914 28866
rect 4062 28702 4114 28754
rect 6862 28702 6914 28754
rect 9102 28702 9154 28754
rect 9550 28702 9602 28754
rect 10110 28702 10162 28754
rect 11678 28702 11730 28754
rect 21870 28702 21922 28754
rect 27582 28702 27634 28754
rect 30158 28702 30210 28754
rect 2046 28590 2098 28642
rect 6190 28590 6242 28642
rect 7310 28590 7362 28642
rect 13470 28590 13522 28642
rect 13918 28590 13970 28642
rect 17278 28590 17330 28642
rect 17726 28590 17778 28642
rect 22542 28590 22594 28642
rect 25902 28590 25954 28642
rect 26238 28590 26290 28642
rect 2270 28478 2322 28530
rect 3054 28478 3106 28530
rect 5742 28478 5794 28530
rect 7758 28478 7810 28530
rect 12798 28478 12850 28530
rect 21310 28478 21362 28530
rect 23550 28478 23602 28530
rect 26798 28478 26850 28530
rect 31166 28478 31218 28530
rect 31950 28478 32002 28530
rect 16494 28366 16546 28418
rect 20078 28366 20130 28418
rect 22766 28366 22818 28418
rect 27134 28366 27186 28418
rect 9026 28198 9078 28250
rect 9130 28198 9182 28250
rect 9234 28198 9286 28250
rect 16838 28198 16890 28250
rect 16942 28198 16994 28250
rect 17046 28198 17098 28250
rect 24650 28198 24702 28250
rect 24754 28198 24806 28250
rect 24858 28198 24910 28250
rect 32462 28198 32514 28250
rect 32566 28198 32618 28250
rect 32670 28198 32722 28250
rect 8990 28030 9042 28082
rect 12574 28030 12626 28082
rect 16382 28030 16434 28082
rect 16942 28030 16994 28082
rect 23326 28030 23378 28082
rect 31502 28030 31554 28082
rect 2158 27918 2210 27970
rect 5182 27918 5234 27970
rect 8654 27918 8706 27970
rect 20078 27918 20130 27970
rect 24110 27918 24162 27970
rect 24334 27918 24386 27970
rect 27246 27918 27298 27970
rect 7422 27806 7474 27858
rect 8094 27806 8146 27858
rect 9662 27806 9714 27858
rect 10110 27806 10162 27858
rect 13358 27806 13410 27858
rect 13806 27806 13858 27858
rect 20638 27806 20690 27858
rect 21086 27806 21138 27858
rect 24558 27806 24610 27858
rect 28590 27806 28642 27858
rect 29262 27806 29314 27858
rect 3166 27694 3218 27746
rect 18734 27694 18786 27746
rect 25342 27694 25394 27746
rect 26238 27694 26290 27746
rect 28030 27694 28082 27746
rect 28366 27694 28418 27746
rect 4398 27582 4450 27634
rect 13134 27582 13186 27634
rect 32286 27582 32338 27634
rect 5120 27414 5172 27466
rect 5224 27414 5276 27466
rect 5328 27414 5380 27466
rect 12932 27414 12984 27466
rect 13036 27414 13088 27466
rect 13140 27414 13192 27466
rect 20744 27414 20796 27466
rect 20848 27414 20900 27466
rect 20952 27414 21004 27466
rect 28556 27414 28608 27466
rect 28660 27414 28712 27466
rect 28764 27414 28816 27466
rect 8766 27246 8818 27298
rect 19742 27246 19794 27298
rect 22206 27246 22258 27298
rect 4062 27134 4114 27186
rect 4510 27134 4562 27186
rect 7534 27134 7586 27186
rect 7982 27134 8034 27186
rect 13694 27134 13746 27186
rect 14814 27134 14866 27186
rect 19966 27134 20018 27186
rect 20750 27134 20802 27186
rect 21646 27134 21698 27186
rect 27582 27134 27634 27186
rect 30718 27134 30770 27186
rect 2046 27022 2098 27074
rect 11902 27022 11954 27074
rect 12462 27022 12514 27074
rect 15598 27022 15650 27074
rect 16270 27022 16322 27074
rect 16606 27022 16658 27074
rect 25230 27022 25282 27074
rect 25678 27022 25730 27074
rect 2270 26910 2322 26962
rect 3054 26910 3106 26962
rect 6526 26910 6578 26962
rect 9550 26910 9602 26962
rect 14030 26910 14082 26962
rect 14366 26910 14418 26962
rect 20302 26910 20354 26962
rect 21310 26910 21362 26962
rect 22990 26910 23042 26962
rect 26574 26910 26626 26962
rect 31950 26910 32002 26962
rect 5742 26798 5794 26850
rect 8542 26798 8594 26850
rect 12686 26798 12738 26850
rect 18958 26798 19010 26850
rect 29374 26798 29426 26850
rect 9026 26630 9078 26682
rect 9130 26630 9182 26682
rect 9234 26630 9286 26682
rect 16838 26630 16890 26682
rect 16942 26630 16994 26682
rect 17046 26630 17098 26682
rect 24650 26630 24702 26682
rect 24754 26630 24806 26682
rect 24858 26630 24910 26682
rect 32462 26630 32514 26682
rect 32566 26630 32618 26682
rect 32670 26630 32722 26682
rect 10222 26462 10274 26514
rect 16382 26462 16434 26514
rect 16942 26462 16994 26514
rect 21310 26462 21362 26514
rect 24110 26462 24162 26514
rect 24558 26462 24610 26514
rect 31278 26462 31330 26514
rect 32174 26462 32226 26514
rect 2382 26350 2434 26402
rect 3166 26350 3218 26402
rect 8318 26350 8370 26402
rect 9102 26350 9154 26402
rect 9886 26350 9938 26402
rect 11006 26350 11058 26402
rect 17390 26350 17442 26402
rect 21982 26350 22034 26402
rect 22318 26350 22370 26402
rect 27246 26350 27298 26402
rect 2158 26238 2210 26290
rect 5630 26238 5682 26290
rect 5966 26238 6018 26290
rect 13022 26238 13074 26290
rect 13358 26238 13410 26290
rect 13918 26238 13970 26290
rect 18286 26238 18338 26290
rect 18846 26238 18898 26290
rect 28366 26238 28418 26290
rect 28814 26238 28866 26290
rect 4174 26126 4226 26178
rect 4734 26126 4786 26178
rect 5070 26126 5122 26178
rect 11902 26126 11954 26178
rect 12462 26126 12514 26178
rect 17726 26126 17778 26178
rect 23438 26126 23490 26178
rect 25454 26126 25506 26178
rect 26238 26126 26290 26178
rect 31838 26014 31890 26066
rect 5120 25846 5172 25898
rect 5224 25846 5276 25898
rect 5328 25846 5380 25898
rect 12932 25846 12984 25898
rect 13036 25846 13088 25898
rect 13140 25846 13192 25898
rect 20744 25846 20796 25898
rect 20848 25846 20900 25898
rect 20952 25846 21004 25898
rect 28556 25846 28608 25898
rect 28660 25846 28712 25898
rect 28764 25846 28816 25898
rect 6078 25678 6130 25730
rect 14590 25678 14642 25730
rect 1934 25566 1986 25618
rect 3838 25566 3890 25618
rect 4734 25566 4786 25618
rect 22654 25678 22706 25730
rect 24894 25678 24946 25730
rect 8094 25566 8146 25618
rect 12574 25566 12626 25618
rect 16494 25566 16546 25618
rect 19294 25566 19346 25618
rect 21758 25566 21810 25618
rect 22094 25566 22146 25618
rect 22654 25566 22706 25618
rect 24334 25566 24386 25618
rect 30158 25566 30210 25618
rect 2942 25454 2994 25506
rect 3390 25454 3442 25506
rect 11118 25454 11170 25506
rect 11790 25454 11842 25506
rect 13806 25454 13858 25506
rect 15262 25454 15314 25506
rect 21534 25454 21586 25506
rect 27918 25454 27970 25506
rect 28366 25454 28418 25506
rect 4958 25342 5010 25394
rect 7422 25342 7474 25394
rect 7758 25342 7810 25394
rect 12014 25342 12066 25394
rect 12798 25342 12850 25394
rect 17502 25342 17554 25394
rect 20302 25342 20354 25394
rect 23214 25342 23266 25394
rect 25678 25342 25730 25394
rect 31502 25342 31554 25394
rect 32174 25342 32226 25394
rect 5742 25230 5794 25282
rect 6862 25230 6914 25282
rect 8878 25230 8930 25282
rect 22206 25230 22258 25282
rect 9026 25062 9078 25114
rect 9130 25062 9182 25114
rect 9234 25062 9286 25114
rect 16838 25062 16890 25114
rect 16942 25062 16994 25114
rect 17046 25062 17098 25114
rect 24650 25062 24702 25114
rect 24754 25062 24806 25114
rect 24858 25062 24910 25114
rect 32462 25062 32514 25114
rect 32566 25062 32618 25114
rect 32670 25062 32722 25114
rect 3726 24894 3778 24946
rect 8094 24894 8146 24946
rect 8878 24894 8930 24946
rect 10782 24894 10834 24946
rect 14702 24894 14754 24946
rect 15486 24894 15538 24946
rect 16830 24894 16882 24946
rect 18958 24894 19010 24946
rect 19742 24894 19794 24946
rect 24446 24894 24498 24946
rect 31726 24894 31778 24946
rect 32286 24894 32338 24946
rect 4958 24782 5010 24834
rect 15262 24782 15314 24834
rect 18062 24782 18114 24834
rect 20526 24782 20578 24834
rect 23662 24782 23714 24834
rect 23998 24782 24050 24834
rect 24334 24782 24386 24834
rect 27246 24782 27298 24834
rect 2942 24670 2994 24722
rect 3726 24670 3778 24722
rect 7310 24670 7362 24722
rect 7758 24670 7810 24722
rect 8990 24670 9042 24722
rect 10222 24670 10274 24722
rect 11566 24670 11618 24722
rect 12126 24670 12178 24722
rect 17502 24670 17554 24722
rect 18398 24670 18450 24722
rect 18958 24670 19010 24722
rect 22878 24670 22930 24722
rect 23214 24670 23266 24722
rect 28590 24670 28642 24722
rect 29262 24670 29314 24722
rect 1934 24558 1986 24610
rect 9774 24558 9826 24610
rect 11342 24558 11394 24610
rect 15934 24558 15986 24610
rect 17614 24558 17666 24610
rect 25342 24558 25394 24610
rect 25790 24558 25842 24610
rect 26238 24558 26290 24610
rect 28030 24558 28082 24610
rect 28366 24558 28418 24610
rect 2158 24446 2210 24498
rect 4174 24446 4226 24498
rect 5120 24278 5172 24330
rect 5224 24278 5276 24330
rect 5328 24278 5380 24330
rect 12932 24278 12984 24330
rect 13036 24278 13088 24330
rect 13140 24278 13192 24330
rect 20744 24278 20796 24330
rect 20848 24278 20900 24330
rect 20952 24278 21004 24330
rect 28556 24278 28608 24330
rect 28660 24278 28712 24330
rect 28764 24278 28816 24330
rect 13022 24110 13074 24162
rect 17054 24110 17106 24162
rect 20862 24110 20914 24162
rect 22990 24110 23042 24162
rect 27134 24110 27186 24162
rect 4062 23998 4114 24050
rect 4510 23998 4562 24050
rect 5966 23998 6018 24050
rect 6302 23998 6354 24050
rect 8094 23998 8146 24050
rect 8654 23998 8706 24050
rect 21646 23998 21698 24050
rect 27806 23998 27858 24050
rect 30158 23998 30210 24050
rect 2046 23886 2098 23938
rect 5070 23886 5122 23938
rect 9550 23886 9602 23938
rect 9998 23886 10050 23938
rect 13470 23886 13522 23938
rect 13918 23886 13970 23938
rect 17166 23886 17218 23938
rect 17838 23886 17890 23938
rect 22094 23886 22146 23938
rect 23550 23886 23602 23938
rect 24110 23886 24162 23938
rect 3054 23774 3106 23826
rect 7086 23774 7138 23826
rect 21310 23774 21362 23826
rect 31502 23774 31554 23826
rect 32062 23774 32114 23826
rect 2270 23662 2322 23714
rect 9102 23662 9154 23714
rect 12462 23662 12514 23714
rect 16382 23662 16434 23714
rect 20302 23662 20354 23714
rect 26574 23662 26626 23714
rect 27358 23662 27410 23714
rect 9026 23494 9078 23546
rect 9130 23494 9182 23546
rect 9234 23494 9286 23546
rect 16838 23494 16890 23546
rect 16942 23494 16994 23546
rect 17046 23494 17098 23546
rect 24650 23494 24702 23546
rect 24754 23494 24806 23546
rect 24858 23494 24910 23546
rect 32462 23494 32514 23546
rect 32566 23494 32618 23546
rect 32670 23494 32722 23546
rect 4174 23326 4226 23378
rect 7422 23326 7474 23378
rect 13358 23326 13410 23378
rect 15150 23326 15202 23378
rect 17726 23326 17778 23378
rect 1822 23214 1874 23266
rect 8654 23214 8706 23266
rect 9550 23214 9602 23266
rect 9886 23214 9938 23266
rect 18062 23214 18114 23266
rect 18398 23214 18450 23266
rect 18734 23214 18786 23266
rect 28926 23214 28978 23266
rect 4622 23102 4674 23154
rect 4958 23102 5010 23154
rect 10222 23102 10274 23154
rect 10782 23102 10834 23154
rect 14142 23102 14194 23154
rect 17502 23102 17554 23154
rect 20862 23102 20914 23154
rect 26686 23102 26738 23154
rect 32174 23102 32226 23154
rect 3054 22990 3106 23042
rect 8430 22990 8482 23042
rect 18958 22990 19010 23042
rect 22318 22990 22370 23042
rect 31502 22990 31554 23042
rect 8094 22878 8146 22930
rect 13918 22878 13970 22930
rect 5120 22710 5172 22762
rect 5224 22710 5276 22762
rect 5328 22710 5380 22762
rect 12932 22710 12984 22762
rect 13036 22710 13088 22762
rect 13140 22710 13192 22762
rect 20744 22710 20796 22762
rect 20848 22710 20900 22762
rect 20952 22710 21004 22762
rect 28556 22710 28608 22762
rect 28660 22710 28712 22762
rect 28764 22710 28816 22762
rect 19630 22542 19682 22594
rect 21198 22542 21250 22594
rect 25006 22542 25058 22594
rect 2046 22430 2098 22482
rect 2270 22430 2322 22482
rect 4062 22430 4114 22482
rect 5070 22430 5122 22482
rect 8542 22430 8594 22482
rect 14030 22430 14082 22482
rect 30158 22430 30210 22482
rect 11566 22318 11618 22370
rect 12798 22318 12850 22370
rect 13582 22318 13634 22370
rect 15038 22318 15090 22370
rect 16158 22318 16210 22370
rect 16494 22318 16546 22370
rect 20526 22318 20578 22370
rect 24222 22318 24274 22370
rect 24670 22318 24722 22370
rect 28142 22318 28194 22370
rect 28702 22318 28754 22370
rect 2830 22206 2882 22258
rect 5854 22206 5906 22258
rect 6190 22206 6242 22258
rect 12574 22206 12626 22258
rect 15374 22206 15426 22258
rect 20750 22206 20802 22258
rect 31166 22206 31218 22258
rect 4622 22094 4674 22146
rect 6526 22094 6578 22146
rect 14702 22094 14754 22146
rect 18958 22094 19010 22146
rect 19966 22094 20018 22146
rect 21982 22094 22034 22146
rect 25566 22094 25618 22146
rect 9026 21926 9078 21978
rect 9130 21926 9182 21978
rect 9234 21926 9286 21978
rect 16838 21926 16890 21978
rect 16942 21926 16994 21978
rect 17046 21926 17098 21978
rect 24650 21926 24702 21978
rect 24754 21926 24806 21978
rect 24858 21926 24910 21978
rect 32462 21926 32514 21978
rect 32566 21926 32618 21978
rect 32670 21926 32722 21978
rect 8542 21758 8594 21810
rect 10334 21758 10386 21810
rect 16718 21758 16770 21810
rect 18062 21758 18114 21810
rect 21198 21758 21250 21810
rect 21982 21758 22034 21810
rect 25118 21758 25170 21810
rect 25678 21758 25730 21810
rect 2382 21646 2434 21698
rect 3166 21646 3218 21698
rect 4622 21646 4674 21698
rect 9886 21646 9938 21698
rect 11790 21646 11842 21698
rect 24446 21646 24498 21698
rect 31054 21646 31106 21698
rect 2158 21534 2210 21586
rect 5630 21534 5682 21586
rect 5966 21534 6018 21586
rect 9102 21534 9154 21586
rect 9550 21534 9602 21586
rect 10558 21534 10610 21586
rect 16270 21534 16322 21586
rect 17838 21534 17890 21586
rect 18398 21534 18450 21586
rect 18958 21534 19010 21586
rect 28254 21534 28306 21586
rect 28702 21534 28754 21586
rect 4174 21422 4226 21474
rect 22318 21422 22370 21474
rect 22766 21422 22818 21474
rect 23214 21422 23266 21474
rect 30046 21422 30098 21474
rect 31950 21422 32002 21474
rect 32174 21422 32226 21474
rect 5120 21142 5172 21194
rect 5224 21142 5276 21194
rect 5328 21142 5380 21194
rect 12932 21142 12984 21194
rect 13036 21142 13088 21194
rect 13140 21142 13192 21194
rect 20744 21142 20796 21194
rect 20848 21142 20900 21194
rect 20952 21142 21004 21194
rect 28556 21142 28608 21194
rect 28660 21142 28712 21194
rect 28764 21142 28816 21194
rect 12238 20974 12290 21026
rect 4062 20862 4114 20914
rect 5742 20862 5794 20914
rect 6862 20862 6914 20914
rect 14254 20862 14306 20914
rect 20526 20862 20578 20914
rect 21870 20862 21922 20914
rect 22094 20862 22146 20914
rect 26686 20862 26738 20914
rect 27918 20862 27970 20914
rect 30606 20862 30658 20914
rect 31502 20862 31554 20914
rect 2046 20750 2098 20802
rect 8766 20750 8818 20802
rect 9102 20750 9154 20802
rect 12574 20750 12626 20802
rect 13806 20750 13858 20802
rect 15150 20750 15202 20802
rect 19070 20750 19122 20802
rect 22542 20750 22594 20802
rect 22990 20750 23042 20802
rect 2270 20638 2322 20690
rect 3054 20638 3106 20690
rect 8206 20638 8258 20690
rect 11454 20638 11506 20690
rect 12798 20638 12850 20690
rect 13470 20638 13522 20690
rect 20750 20638 20802 20690
rect 21422 20638 21474 20690
rect 26350 20638 26402 20690
rect 29486 20638 29538 20690
rect 4622 20526 4674 20578
rect 6414 20526 6466 20578
rect 17502 20526 17554 20578
rect 25566 20526 25618 20578
rect 26126 20526 26178 20578
rect 27358 20526 27410 20578
rect 9026 20358 9078 20410
rect 9130 20358 9182 20410
rect 9234 20358 9286 20410
rect 16838 20358 16890 20410
rect 16942 20358 16994 20410
rect 17046 20358 17098 20410
rect 24650 20358 24702 20410
rect 24754 20358 24806 20410
rect 24858 20358 24910 20410
rect 32462 20358 32514 20410
rect 32566 20358 32618 20410
rect 32670 20358 32722 20410
rect 8430 20190 8482 20242
rect 15374 20190 15426 20242
rect 23102 20190 23154 20242
rect 2382 20078 2434 20130
rect 9662 20078 9714 20130
rect 12014 20078 12066 20130
rect 15934 20078 15986 20130
rect 19406 20078 19458 20130
rect 22206 20078 22258 20130
rect 23438 20078 23490 20130
rect 25342 20078 25394 20130
rect 28478 20078 28530 20130
rect 29262 20078 29314 20130
rect 31502 20078 31554 20130
rect 4734 19966 4786 20018
rect 5294 19966 5346 20018
rect 5630 19966 5682 20018
rect 5966 19966 6018 20018
rect 12238 19966 12290 20018
rect 12798 19966 12850 20018
rect 25566 19966 25618 20018
rect 26238 19966 26290 20018
rect 9102 19854 9154 19906
rect 11006 19854 11058 19906
rect 11454 19854 11506 19906
rect 16494 19854 16546 19906
rect 16830 19854 16882 19906
rect 17502 19854 17554 19906
rect 18398 19854 18450 19906
rect 20974 19854 21026 19906
rect 21198 19854 21250 19906
rect 24334 19854 24386 19906
rect 30494 19854 30546 19906
rect 1598 19742 1650 19794
rect 5120 19574 5172 19626
rect 5224 19574 5276 19626
rect 5328 19574 5380 19626
rect 12932 19574 12984 19626
rect 13036 19574 13088 19626
rect 13140 19574 13192 19626
rect 20744 19574 20796 19626
rect 20848 19574 20900 19626
rect 20952 19574 21004 19626
rect 28556 19574 28608 19626
rect 28660 19574 28712 19626
rect 28764 19574 28816 19626
rect 12238 19406 12290 19458
rect 13022 19406 13074 19458
rect 14478 19406 14530 19458
rect 24894 19406 24946 19458
rect 4062 19294 4114 19346
rect 4510 19294 4562 19346
rect 9774 19294 9826 19346
rect 11902 19294 11954 19346
rect 12462 19294 12514 19346
rect 12910 19294 12962 19346
rect 30158 19294 30210 19346
rect 2046 19182 2098 19234
rect 5630 19182 5682 19234
rect 6078 19182 6130 19234
rect 13694 19182 13746 19234
rect 17614 19182 17666 19234
rect 18062 19182 18114 19234
rect 18958 19182 19010 19234
rect 19742 19182 19794 19234
rect 20526 19182 20578 19234
rect 21198 19182 21250 19234
rect 21870 19182 21922 19234
rect 25006 19182 25058 19234
rect 25678 19182 25730 19234
rect 28702 19182 28754 19234
rect 2718 19070 2770 19122
rect 10894 19070 10946 19122
rect 13470 19070 13522 19122
rect 15262 19070 15314 19122
rect 19182 19070 19234 19122
rect 19518 19070 19570 19122
rect 20750 19070 20802 19122
rect 31166 19070 31218 19122
rect 2046 18958 2098 19010
rect 8654 18958 8706 19010
rect 9214 18958 9266 19010
rect 9886 18958 9938 19010
rect 18510 18958 18562 19010
rect 24334 18958 24386 19010
rect 27918 18958 27970 19010
rect 29262 18958 29314 19010
rect 32062 18958 32114 19010
rect 9026 18790 9078 18842
rect 9130 18790 9182 18842
rect 9234 18790 9286 18842
rect 16838 18790 16890 18842
rect 16942 18790 16994 18842
rect 17046 18790 17098 18842
rect 24650 18790 24702 18842
rect 24754 18790 24806 18842
rect 24858 18790 24910 18842
rect 32462 18790 32514 18842
rect 32566 18790 32618 18842
rect 32670 18790 32722 18842
rect 1934 18622 1986 18674
rect 2158 18622 2210 18674
rect 9438 18622 9490 18674
rect 16382 18622 16434 18674
rect 28142 18622 28194 18674
rect 6414 18510 6466 18562
rect 10222 18510 10274 18562
rect 17390 18510 17442 18562
rect 21310 18510 21362 18562
rect 24334 18510 24386 18562
rect 26686 18510 26738 18562
rect 27358 18510 27410 18562
rect 31838 18510 31890 18562
rect 2942 18398 2994 18450
rect 3726 18398 3778 18450
rect 4062 18398 4114 18450
rect 7422 18398 7474 18450
rect 8990 18398 9042 18450
rect 12462 18398 12514 18450
rect 13022 18398 13074 18450
rect 13246 18398 13298 18450
rect 13918 18398 13970 18450
rect 17614 18398 17666 18450
rect 18510 18398 18562 18450
rect 19070 18398 19122 18450
rect 22430 18398 22482 18450
rect 22878 18398 22930 18450
rect 24558 18398 24610 18450
rect 25566 18398 25618 18450
rect 26462 18398 26514 18450
rect 27134 18398 27186 18450
rect 30606 18398 30658 18450
rect 31278 18398 31330 18450
rect 31502 18398 31554 18450
rect 7870 18286 7922 18338
rect 18174 18286 18226 18338
rect 25678 18286 25730 18338
rect 27582 18286 27634 18338
rect 7198 18174 7250 18226
rect 16942 18174 16994 18226
rect 22094 18174 22146 18226
rect 23326 18174 23378 18226
rect 5120 18006 5172 18058
rect 5224 18006 5276 18058
rect 5328 18006 5380 18058
rect 12932 18006 12984 18058
rect 13036 18006 13088 18058
rect 13140 18006 13192 18058
rect 20744 18006 20796 18058
rect 20848 18006 20900 18058
rect 20952 18006 21004 18058
rect 28556 18006 28608 18058
rect 28660 18006 28712 18058
rect 28764 18006 28816 18058
rect 20302 17838 20354 17890
rect 1934 17726 1986 17778
rect 3950 17726 4002 17778
rect 4510 17726 4562 17778
rect 5070 17726 5122 17778
rect 5742 17726 5794 17778
rect 6414 17726 6466 17778
rect 7422 17726 7474 17778
rect 11678 17726 11730 17778
rect 12126 17726 12178 17778
rect 15374 17726 15426 17778
rect 20750 17726 20802 17778
rect 21310 17726 21362 17778
rect 26574 17726 26626 17778
rect 30158 17726 30210 17778
rect 32062 17726 32114 17778
rect 7646 17614 7698 17666
rect 8206 17614 8258 17666
rect 12350 17614 12402 17666
rect 16606 17614 16658 17666
rect 17166 17614 17218 17666
rect 21534 17614 21586 17666
rect 22206 17614 22258 17666
rect 22654 17614 22706 17666
rect 23326 17614 23378 17666
rect 27358 17614 27410 17666
rect 28590 17614 28642 17666
rect 29262 17614 29314 17666
rect 2270 17502 2322 17554
rect 3054 17502 3106 17554
rect 10558 17502 10610 17554
rect 14366 17502 14418 17554
rect 19518 17502 19570 17554
rect 21982 17502 22034 17554
rect 26350 17502 26402 17554
rect 26910 17502 26962 17554
rect 28366 17502 28418 17554
rect 31166 17502 31218 17554
rect 6862 17390 6914 17442
rect 11342 17390 11394 17442
rect 12910 17390 12962 17442
rect 13582 17390 13634 17442
rect 15822 17390 15874 17442
rect 16270 17390 16322 17442
rect 25678 17390 25730 17442
rect 29710 17390 29762 17442
rect 9026 17222 9078 17274
rect 9130 17222 9182 17274
rect 9234 17222 9286 17274
rect 16838 17222 16890 17274
rect 16942 17222 16994 17274
rect 17046 17222 17098 17274
rect 24650 17222 24702 17274
rect 24754 17222 24806 17274
rect 24858 17222 24910 17274
rect 32462 17222 32514 17274
rect 32566 17222 32618 17274
rect 32670 17222 32722 17274
rect 1598 17054 1650 17106
rect 2270 17054 2322 17106
rect 5406 17054 5458 17106
rect 14366 17054 14418 17106
rect 16830 17054 16882 17106
rect 28030 17054 28082 17106
rect 29150 17054 29202 17106
rect 6190 16942 6242 16994
rect 10670 16942 10722 16994
rect 11006 16942 11058 16994
rect 15262 16942 15314 16994
rect 22990 16942 23042 16994
rect 23326 16942 23378 16994
rect 23662 16942 23714 16994
rect 24334 16942 24386 16994
rect 31054 16942 31106 16994
rect 31838 16942 31890 16994
rect 4734 16830 4786 16882
rect 5294 16830 5346 16882
rect 8430 16830 8482 16882
rect 8878 16830 8930 16882
rect 9774 16830 9826 16882
rect 11454 16830 11506 16882
rect 11790 16830 11842 16882
rect 15486 16830 15538 16882
rect 15934 16830 15986 16882
rect 16158 16830 16210 16882
rect 17502 16830 17554 16882
rect 25342 16830 25394 16882
rect 25790 16830 25842 16882
rect 32062 16830 32114 16882
rect 21646 16718 21698 16770
rect 23998 16718 24050 16770
rect 24670 16718 24722 16770
rect 30046 16718 30098 16770
rect 9662 16606 9714 16658
rect 14926 16606 14978 16658
rect 28814 16606 28866 16658
rect 5120 16438 5172 16490
rect 5224 16438 5276 16490
rect 5328 16438 5380 16490
rect 12932 16438 12984 16490
rect 13036 16438 13088 16490
rect 13140 16438 13192 16490
rect 20744 16438 20796 16490
rect 20848 16438 20900 16490
rect 20952 16438 21004 16490
rect 28556 16438 28608 16490
rect 28660 16438 28712 16490
rect 28764 16438 28816 16490
rect 13918 16270 13970 16322
rect 25006 16270 25058 16322
rect 3950 16158 4002 16210
rect 4734 16158 4786 16210
rect 5070 16158 5122 16210
rect 6974 16158 7026 16210
rect 29822 16270 29874 16322
rect 13022 16158 13074 16210
rect 19406 16158 19458 16210
rect 29150 16158 29202 16210
rect 29262 16158 29314 16210
rect 29822 16158 29874 16210
rect 30158 16158 30210 16210
rect 32062 16158 32114 16210
rect 1934 16046 1986 16098
rect 5966 16046 6018 16098
rect 7422 16046 7474 16098
rect 11230 16046 11282 16098
rect 11902 16046 11954 16098
rect 14814 16046 14866 16098
rect 15486 16046 15538 16098
rect 16158 16046 16210 16098
rect 19630 16046 19682 16098
rect 20302 16046 20354 16098
rect 21422 16046 21474 16098
rect 21870 16046 21922 16098
rect 28142 16046 28194 16098
rect 28702 16046 28754 16098
rect 3054 15934 3106 15986
rect 12126 15934 12178 15986
rect 12462 15934 12514 15986
rect 20078 15934 20130 15986
rect 24894 15934 24946 15986
rect 31166 15934 31218 15986
rect 2270 15822 2322 15874
rect 5742 15822 5794 15874
rect 7310 15822 7362 15874
rect 8206 15822 8258 15874
rect 8990 15822 9042 15874
rect 18398 15822 18450 15874
rect 19182 15822 19234 15874
rect 24110 15822 24162 15874
rect 25566 15822 25618 15874
rect 9026 15654 9078 15706
rect 9130 15654 9182 15706
rect 9234 15654 9286 15706
rect 16838 15654 16890 15706
rect 16942 15654 16994 15706
rect 17046 15654 17098 15706
rect 24650 15654 24702 15706
rect 24754 15654 24806 15706
rect 24858 15654 24910 15706
rect 32462 15654 32514 15706
rect 32566 15654 32618 15706
rect 32670 15654 32722 15706
rect 2158 15486 2210 15538
rect 8990 15486 9042 15538
rect 9886 15486 9938 15538
rect 12574 15486 12626 15538
rect 18062 15486 18114 15538
rect 21534 15486 21586 15538
rect 22542 15486 22594 15538
rect 24110 15486 24162 15538
rect 26126 15486 26178 15538
rect 26910 15486 26962 15538
rect 6190 15374 6242 15426
rect 6638 15374 6690 15426
rect 10894 15374 10946 15426
rect 18174 15374 18226 15426
rect 22878 15374 22930 15426
rect 23214 15374 23266 15426
rect 23550 15374 23602 15426
rect 24334 15374 24386 15426
rect 24670 15374 24722 15426
rect 4622 15262 4674 15314
rect 5070 15262 5122 15314
rect 5966 15262 6018 15314
rect 8542 15262 8594 15314
rect 9774 15262 9826 15314
rect 11118 15262 11170 15314
rect 14814 15262 14866 15314
rect 15486 15262 15538 15314
rect 16494 15262 16546 15314
rect 18622 15262 18674 15314
rect 19070 15262 19122 15314
rect 25454 15262 25506 15314
rect 29374 15262 29426 15314
rect 29822 15262 29874 15314
rect 30718 15262 30770 15314
rect 31614 15262 31666 15314
rect 7982 15150 8034 15202
rect 16046 15150 16098 15202
rect 17502 15150 17554 15202
rect 25230 15150 25282 15202
rect 30830 15150 30882 15202
rect 1598 15038 1650 15090
rect 11790 15038 11842 15090
rect 22094 15038 22146 15090
rect 26350 15038 26402 15090
rect 31502 15038 31554 15090
rect 5120 14870 5172 14922
rect 5224 14870 5276 14922
rect 5328 14870 5380 14922
rect 12932 14870 12984 14922
rect 13036 14870 13088 14922
rect 13140 14870 13192 14922
rect 20744 14870 20796 14922
rect 20848 14870 20900 14922
rect 20952 14870 21004 14922
rect 28556 14870 28608 14922
rect 28660 14870 28712 14922
rect 28764 14870 28816 14922
rect 25678 14702 25730 14754
rect 4062 14590 4114 14642
rect 5182 14590 5234 14642
rect 14814 14590 14866 14642
rect 26126 14590 26178 14642
rect 26462 14590 26514 14642
rect 26910 14590 26962 14642
rect 30158 14590 30210 14642
rect 5518 14478 5570 14530
rect 8542 14478 8594 14530
rect 9214 14478 9266 14530
rect 9550 14478 9602 14530
rect 9886 14478 9938 14530
rect 16606 14478 16658 14530
rect 17166 14478 17218 14530
rect 21534 14478 21586 14530
rect 21982 14478 22034 14530
rect 22654 14478 22706 14530
rect 2270 14366 2322 14418
rect 2718 14366 2770 14418
rect 6302 14366 6354 14418
rect 15822 14366 15874 14418
rect 20414 14366 20466 14418
rect 20750 14366 20802 14418
rect 21758 14366 21810 14418
rect 27918 14366 27970 14418
rect 31502 14366 31554 14418
rect 1934 14254 1986 14306
rect 4622 14254 4674 14306
rect 12462 14254 12514 14306
rect 13022 14254 13074 14306
rect 13582 14254 13634 14306
rect 14030 14254 14082 14306
rect 14478 14254 14530 14306
rect 19630 14254 19682 14306
rect 20190 14254 20242 14306
rect 25118 14254 25170 14306
rect 29822 14254 29874 14306
rect 32062 14254 32114 14306
rect 9026 14086 9078 14138
rect 9130 14086 9182 14138
rect 9234 14086 9286 14138
rect 16838 14086 16890 14138
rect 16942 14086 16994 14138
rect 17046 14086 17098 14138
rect 24650 14086 24702 14138
rect 24754 14086 24806 14138
rect 24858 14086 24910 14138
rect 32462 14086 32514 14138
rect 32566 14086 32618 14138
rect 32670 14086 32722 14138
rect 2382 13918 2434 13970
rect 9886 13918 9938 13970
rect 12350 13918 12402 13970
rect 16046 13918 16098 13970
rect 17390 13918 17442 13970
rect 18062 13918 18114 13970
rect 23326 13918 23378 13970
rect 24110 13918 24162 13970
rect 5406 13806 5458 13858
rect 6190 13806 6242 13858
rect 9550 13806 9602 13858
rect 10782 13806 10834 13858
rect 29710 13806 29762 13858
rect 4622 13694 4674 13746
rect 5294 13694 5346 13746
rect 8430 13694 8482 13746
rect 8878 13694 8930 13746
rect 13358 13694 13410 13746
rect 13694 13694 13746 13746
rect 17726 13694 17778 13746
rect 18286 13694 18338 13746
rect 18846 13694 18898 13746
rect 25678 13694 25730 13746
rect 26462 13694 26514 13746
rect 11790 13582 11842 13634
rect 12798 13582 12850 13634
rect 22542 13582 22594 13634
rect 24670 13582 24722 13634
rect 1598 13470 1650 13522
rect 16830 13470 16882 13522
rect 25902 13470 25954 13522
rect 5120 13302 5172 13354
rect 5224 13302 5276 13354
rect 5328 13302 5380 13354
rect 12932 13302 12984 13354
rect 13036 13302 13088 13354
rect 13140 13302 13192 13354
rect 20744 13302 20796 13354
rect 20848 13302 20900 13354
rect 20952 13302 21004 13354
rect 28556 13302 28608 13354
rect 28660 13302 28712 13354
rect 28764 13302 28816 13354
rect 2494 13022 2546 13074
rect 3838 13022 3890 13074
rect 6190 13022 6242 13074
rect 6974 13022 7026 13074
rect 8094 13022 8146 13074
rect 9998 13022 10050 13074
rect 11902 13022 11954 13074
rect 13582 13022 13634 13074
rect 15374 13022 15426 13074
rect 16718 13022 16770 13074
rect 18510 13022 18562 13074
rect 18958 13022 19010 13074
rect 19294 13022 19346 13074
rect 21422 13022 21474 13074
rect 21870 13022 21922 13074
rect 30382 13022 30434 13074
rect 1710 12910 1762 12962
rect 2942 12910 2994 12962
rect 5966 12910 6018 12962
rect 13694 12910 13746 12962
rect 14814 12910 14866 12962
rect 26462 12910 26514 12962
rect 27806 12910 27858 12962
rect 2046 12798 2098 12850
rect 4958 12798 5010 12850
rect 9102 12798 9154 12850
rect 10894 12798 10946 12850
rect 14590 12798 14642 12850
rect 17502 12798 17554 12850
rect 20526 12798 20578 12850
rect 23662 12798 23714 12850
rect 29486 12798 29538 12850
rect 7422 12686 7474 12738
rect 12462 12686 12514 12738
rect 12910 12686 12962 12738
rect 16158 12686 16210 12738
rect 27918 12686 27970 12738
rect 9026 12518 9078 12570
rect 9130 12518 9182 12570
rect 9234 12518 9286 12570
rect 16838 12518 16890 12570
rect 16942 12518 16994 12570
rect 17046 12518 17098 12570
rect 24650 12518 24702 12570
rect 24754 12518 24806 12570
rect 24858 12518 24910 12570
rect 32462 12518 32514 12570
rect 32566 12518 32618 12570
rect 32670 12518 32722 12570
rect 5518 12350 5570 12402
rect 8990 12350 9042 12402
rect 16270 12350 16322 12402
rect 25902 12350 25954 12402
rect 29598 12350 29650 12402
rect 2382 12238 2434 12290
rect 6862 12238 6914 12290
rect 17390 12238 17442 12290
rect 20862 12238 20914 12290
rect 23886 12238 23938 12290
rect 31278 12238 31330 12290
rect 4622 12126 4674 12178
rect 5070 12126 5122 12178
rect 5742 12126 5794 12178
rect 12798 12126 12850 12178
rect 14366 12126 14418 12178
rect 15150 12126 15202 12178
rect 16494 12126 16546 12178
rect 17614 12126 17666 12178
rect 18174 12126 18226 12178
rect 18622 12126 18674 12178
rect 28254 12126 28306 12178
rect 28814 12126 28866 12178
rect 29150 12126 29202 12178
rect 7982 12014 8034 12066
rect 10446 12014 10498 12066
rect 14030 12014 14082 12066
rect 14926 12014 14978 12066
rect 22878 12014 22930 12066
rect 30270 12014 30322 12066
rect 1598 11902 1650 11954
rect 15262 11902 15314 11954
rect 21646 11902 21698 11954
rect 25118 11902 25170 11954
rect 5120 11734 5172 11786
rect 5224 11734 5276 11786
rect 5328 11734 5380 11786
rect 12932 11734 12984 11786
rect 13036 11734 13088 11786
rect 13140 11734 13192 11786
rect 20744 11734 20796 11786
rect 20848 11734 20900 11786
rect 20952 11734 21004 11786
rect 28556 11734 28608 11786
rect 28660 11734 28712 11786
rect 28764 11734 28816 11786
rect 5742 11566 5794 11618
rect 18958 11566 19010 11618
rect 3838 11454 3890 11506
rect 4510 11454 4562 11506
rect 5070 11454 5122 11506
rect 11678 11454 11730 11506
rect 1934 11342 1986 11394
rect 5966 11342 6018 11394
rect 9438 11342 9490 11394
rect 12910 11342 12962 11394
rect 13470 11342 13522 11394
rect 20414 11566 20466 11618
rect 29262 11454 29314 11506
rect 30158 11454 30210 11506
rect 32062 11454 32114 11506
rect 19742 11342 19794 11394
rect 20526 11342 20578 11394
rect 21198 11342 21250 11394
rect 21870 11342 21922 11394
rect 25230 11342 25282 11394
rect 25678 11342 25730 11394
rect 2270 11230 2322 11282
rect 3054 11230 3106 11282
rect 15822 11230 15874 11282
rect 27918 11230 27970 11282
rect 31166 11230 31218 11282
rect 6750 11118 6802 11170
rect 7310 11118 7362 11170
rect 19182 11118 19234 11170
rect 24110 11118 24162 11170
rect 24894 11118 24946 11170
rect 28702 11118 28754 11170
rect 9026 10950 9078 11002
rect 9130 10950 9182 11002
rect 9234 10950 9286 11002
rect 16838 10950 16890 11002
rect 16942 10950 16994 11002
rect 17046 10950 17098 11002
rect 24650 10950 24702 11002
rect 24754 10950 24806 11002
rect 24858 10950 24910 11002
rect 32462 10950 32514 11002
rect 32566 10950 32618 11002
rect 32670 10950 32722 11002
rect 4734 10782 4786 10834
rect 6190 10782 6242 10834
rect 9662 10782 9714 10834
rect 10110 10782 10162 10834
rect 10558 10782 10610 10834
rect 22318 10782 22370 10834
rect 30270 10782 30322 10834
rect 16270 10670 16322 10722
rect 20974 10670 21026 10722
rect 23886 10670 23938 10722
rect 25566 10670 25618 10722
rect 29038 10670 29090 10722
rect 30606 10670 30658 10722
rect 32286 10670 32338 10722
rect 1710 10558 1762 10610
rect 2158 10558 2210 10610
rect 8542 10558 8594 10610
rect 9102 10558 9154 10610
rect 10894 10558 10946 10610
rect 15150 10558 15202 10610
rect 16494 10558 16546 10610
rect 18174 10558 18226 10610
rect 19406 10558 19458 10610
rect 25902 10558 25954 10610
rect 26350 10558 26402 10610
rect 26798 10558 26850 10610
rect 30942 10558 30994 10610
rect 15262 10446 15314 10498
rect 18958 10446 19010 10498
rect 19966 10446 20018 10498
rect 21870 10446 21922 10498
rect 22878 10446 22930 10498
rect 5294 10334 5346 10386
rect 5406 10334 5458 10386
rect 9662 10334 9714 10386
rect 10670 10334 10722 10386
rect 13694 10334 13746 10386
rect 18062 10334 18114 10386
rect 29822 10334 29874 10386
rect 31726 10334 31778 10386
rect 5120 10166 5172 10218
rect 5224 10166 5276 10218
rect 5328 10166 5380 10218
rect 12932 10166 12984 10218
rect 13036 10166 13088 10218
rect 13140 10166 13192 10218
rect 20744 10166 20796 10218
rect 20848 10166 20900 10218
rect 20952 10166 21004 10218
rect 28556 10166 28608 10218
rect 28660 10166 28712 10218
rect 28764 10166 28816 10218
rect 18958 9998 19010 10050
rect 23102 9998 23154 10050
rect 3950 9886 4002 9938
rect 4622 9886 4674 9938
rect 9102 9886 9154 9938
rect 29822 9886 29874 9938
rect 30158 9886 30210 9938
rect 32174 9886 32226 9938
rect 2046 9774 2098 9826
rect 6638 9774 6690 9826
rect 8318 9774 8370 9826
rect 13470 9774 13522 9826
rect 14814 9774 14866 9826
rect 15262 9774 15314 9826
rect 15934 9774 15986 9826
rect 19406 9774 19458 9826
rect 20750 9774 20802 9826
rect 21534 9774 21586 9826
rect 22990 9774 23042 9826
rect 23662 9774 23714 9826
rect 23998 9774 24050 9826
rect 27358 9774 27410 9826
rect 2270 9662 2322 9714
rect 3054 9662 3106 9714
rect 18174 9662 18226 9714
rect 31166 9662 31218 9714
rect 5070 9550 5122 9602
rect 6638 9550 6690 9602
rect 12686 9550 12738 9602
rect 13582 9550 13634 9602
rect 14590 9550 14642 9602
rect 19182 9550 19234 9602
rect 20638 9550 20690 9602
rect 21422 9550 21474 9602
rect 26462 9550 26514 9602
rect 27134 9550 27186 9602
rect 27470 9550 27522 9602
rect 28590 9550 28642 9602
rect 9026 9382 9078 9434
rect 9130 9382 9182 9434
rect 9234 9382 9286 9434
rect 16838 9382 16890 9434
rect 16942 9382 16994 9434
rect 17046 9382 17098 9434
rect 24650 9382 24702 9434
rect 24754 9382 24806 9434
rect 24858 9382 24910 9434
rect 32462 9382 32514 9434
rect 32566 9382 32618 9434
rect 32670 9382 32722 9434
rect 4510 9214 4562 9266
rect 8318 9214 8370 9266
rect 10446 9214 10498 9266
rect 10894 9214 10946 9266
rect 11230 9214 11282 9266
rect 21198 9214 21250 9266
rect 22318 9214 22370 9266
rect 22878 9214 22930 9266
rect 26462 9214 26514 9266
rect 27582 9214 27634 9266
rect 30830 9214 30882 9266
rect 31502 9214 31554 9266
rect 31726 9214 31778 9266
rect 9550 9102 9602 9154
rect 12798 9102 12850 9154
rect 16158 9102 16210 9154
rect 17390 9102 17442 9154
rect 17726 9102 17778 9154
rect 24222 9102 24274 9154
rect 32062 9102 32114 9154
rect 1822 8990 1874 9042
rect 2270 8990 2322 9042
rect 5406 8990 5458 9042
rect 6078 8990 6130 9042
rect 9774 8990 9826 9042
rect 13246 8990 13298 9042
rect 13918 8990 13970 9042
rect 18286 8990 18338 9042
rect 18958 8990 19010 9042
rect 25230 8990 25282 9042
rect 26350 8990 26402 9042
rect 28030 8990 28082 9042
rect 28366 8990 28418 9042
rect 11678 8878 11730 8930
rect 23214 8878 23266 8930
rect 5294 8766 5346 8818
rect 9102 8766 9154 8818
rect 16942 8766 16994 8818
rect 21982 8766 22034 8818
rect 25342 8766 25394 8818
rect 5120 8598 5172 8650
rect 5224 8598 5276 8650
rect 5328 8598 5380 8650
rect 12932 8598 12984 8650
rect 13036 8598 13088 8650
rect 13140 8598 13192 8650
rect 20744 8598 20796 8650
rect 20848 8598 20900 8650
rect 20952 8598 21004 8650
rect 28556 8598 28608 8650
rect 28660 8598 28712 8650
rect 28764 8598 28816 8650
rect 13022 8430 13074 8482
rect 4062 8318 4114 8370
rect 5070 8318 5122 8370
rect 14814 8318 14866 8370
rect 19294 8318 19346 8370
rect 29710 8318 29762 8370
rect 30270 8318 30322 8370
rect 5518 8206 5570 8258
rect 6078 8206 6130 8258
rect 9438 8206 9490 8258
rect 9886 8206 9938 8258
rect 14254 8206 14306 8258
rect 15038 8206 15090 8258
rect 15822 8206 15874 8258
rect 16270 8206 16322 8258
rect 19518 8206 19570 8258
rect 21198 8206 21250 8258
rect 21870 8206 21922 8258
rect 24894 8206 24946 8258
rect 28142 8206 28194 8258
rect 28702 8206 28754 8258
rect 1934 8094 1986 8146
rect 2270 8094 2322 8146
rect 2718 8094 2770 8146
rect 25790 8094 25842 8146
rect 31166 8094 31218 8146
rect 8654 7982 8706 8034
rect 9214 7982 9266 8034
rect 12462 7982 12514 8034
rect 14142 7982 14194 8034
rect 18734 7982 18786 8034
rect 19630 7982 19682 8034
rect 20750 7982 20802 8034
rect 24334 7982 24386 8034
rect 25006 7982 25058 8034
rect 29262 7982 29314 8034
rect 32062 7982 32114 8034
rect 9026 7814 9078 7866
rect 9130 7814 9182 7866
rect 9234 7814 9286 7866
rect 16838 7814 16890 7866
rect 16942 7814 16994 7866
rect 17046 7814 17098 7866
rect 24650 7814 24702 7866
rect 24754 7814 24806 7866
rect 24858 7814 24910 7866
rect 32462 7814 32514 7866
rect 32566 7814 32618 7866
rect 32670 7814 32722 7866
rect 1822 7646 1874 7698
rect 7422 7646 7474 7698
rect 8654 7646 8706 7698
rect 9662 7646 9714 7698
rect 10782 7646 10834 7698
rect 14142 7646 14194 7698
rect 15262 7646 15314 7698
rect 16830 7646 16882 7698
rect 17950 7646 18002 7698
rect 24670 7646 24722 7698
rect 31166 7646 31218 7698
rect 3950 7534 4002 7586
rect 19406 7534 19458 7586
rect 20862 7534 20914 7586
rect 27582 7534 27634 7586
rect 4622 7422 4674 7474
rect 5070 7422 5122 7474
rect 8430 7422 8482 7474
rect 11118 7422 11170 7474
rect 11678 7422 11730 7474
rect 16046 7422 16098 7474
rect 23214 7422 23266 7474
rect 23550 7422 23602 7474
rect 24334 7422 24386 7474
rect 28478 7422 28530 7474
rect 28926 7422 28978 7474
rect 2718 7310 2770 7362
rect 10110 7310 10162 7362
rect 16158 7310 16210 7362
rect 17502 7310 17554 7362
rect 18398 7310 18450 7362
rect 26238 7310 26290 7362
rect 8094 7198 8146 7250
rect 14814 7198 14866 7250
rect 20078 7198 20130 7250
rect 31950 7198 32002 7250
rect 5120 7030 5172 7082
rect 5224 7030 5276 7082
rect 5328 7030 5380 7082
rect 12932 7030 12984 7082
rect 13036 7030 13088 7082
rect 13140 7030 13192 7082
rect 20744 7030 20796 7082
rect 20848 7030 20900 7082
rect 20952 7030 21004 7082
rect 28556 7030 28608 7082
rect 28660 7030 28712 7082
rect 28764 7030 28816 7082
rect 4062 6750 4114 6802
rect 5070 6750 5122 6802
rect 11230 6750 11282 6802
rect 14254 6750 14306 6802
rect 15486 6750 15538 6802
rect 19182 6750 19234 6802
rect 23102 6750 23154 6802
rect 25902 6750 25954 6802
rect 30158 6750 30210 6802
rect 1822 6638 1874 6690
rect 6302 6638 6354 6690
rect 6862 6638 6914 6690
rect 10334 6638 10386 6690
rect 10782 6638 10834 6690
rect 18846 6638 18898 6690
rect 21534 6638 21586 6690
rect 28254 6638 28306 6690
rect 2046 6526 2098 6578
rect 3054 6526 3106 6578
rect 5630 6526 5682 6578
rect 5966 6526 6018 6578
rect 12238 6526 12290 6578
rect 13470 6526 13522 6578
rect 13806 6526 13858 6578
rect 14702 6526 14754 6578
rect 16718 6526 16770 6578
rect 17502 6526 17554 6578
rect 20190 6526 20242 6578
rect 24110 6526 24162 6578
rect 26910 6526 26962 6578
rect 28478 6526 28530 6578
rect 31502 6526 31554 6578
rect 4510 6414 4562 6466
rect 9438 6414 9490 6466
rect 9998 6414 10050 6466
rect 15150 6414 15202 6466
rect 17838 6414 17890 6466
rect 18286 6414 18338 6466
rect 21758 6414 21810 6466
rect 22318 6414 22370 6466
rect 32062 6414 32114 6466
rect 9026 6246 9078 6298
rect 9130 6246 9182 6298
rect 9234 6246 9286 6298
rect 16838 6246 16890 6298
rect 16942 6246 16994 6298
rect 17046 6246 17098 6298
rect 24650 6246 24702 6298
rect 24754 6246 24806 6298
rect 24858 6246 24910 6298
rect 32462 6246 32514 6298
rect 32566 6246 32618 6298
rect 32670 6246 32722 6298
rect 3614 6078 3666 6130
rect 4062 6078 4114 6130
rect 8094 6078 8146 6130
rect 9550 6078 9602 6130
rect 14926 6078 14978 6130
rect 27582 6078 27634 6130
rect 28366 6078 28418 6130
rect 29150 6078 29202 6130
rect 4846 5966 4898 6018
rect 13358 5966 13410 6018
rect 14478 5966 14530 6018
rect 16382 5966 16434 6018
rect 20190 5966 20242 6018
rect 20974 5966 21026 6018
rect 21870 5966 21922 6018
rect 22318 5966 22370 6018
rect 25342 5966 25394 6018
rect 25790 5966 25842 6018
rect 2942 5854 2994 5906
rect 3390 5854 3442 5906
rect 7198 5854 7250 5906
rect 7534 5854 7586 5906
rect 8094 5854 8146 5906
rect 9774 5854 9826 5906
rect 10670 5854 10722 5906
rect 11118 5854 11170 5906
rect 17502 5854 17554 5906
rect 17838 5854 17890 5906
rect 21646 5854 21698 5906
rect 31390 5854 31442 5906
rect 32062 5854 32114 5906
rect 1934 5742 1986 5794
rect 15374 5742 15426 5794
rect 23438 5742 23490 5794
rect 27134 5742 27186 5794
rect 14142 5630 14194 5682
rect 5120 5462 5172 5514
rect 5224 5462 5276 5514
rect 5328 5462 5380 5514
rect 12932 5462 12984 5514
rect 13036 5462 13088 5514
rect 13140 5462 13192 5514
rect 20744 5462 20796 5514
rect 20848 5462 20900 5514
rect 20952 5462 21004 5514
rect 28556 5462 28608 5514
rect 28660 5462 28712 5514
rect 28764 5462 28816 5514
rect 12798 5294 12850 5346
rect 18174 5294 18226 5346
rect 19742 5294 19794 5346
rect 21982 5294 22034 5346
rect 23774 5294 23826 5346
rect 2158 5182 2210 5234
rect 3950 5182 4002 5234
rect 4734 5182 4786 5234
rect 6974 5182 7026 5234
rect 24334 5182 24386 5234
rect 25342 5182 25394 5234
rect 27582 5182 27634 5234
rect 29822 5182 29874 5234
rect 30158 5182 30210 5234
rect 32062 5182 32114 5234
rect 6414 5070 6466 5122
rect 11230 5070 11282 5122
rect 11678 5070 11730 5122
rect 12574 5070 12626 5122
rect 13918 5070 13970 5122
rect 14702 5070 14754 5122
rect 15150 5070 15202 5122
rect 18510 5070 18562 5122
rect 19854 5070 19906 5122
rect 20414 5070 20466 5122
rect 22094 5070 22146 5122
rect 23102 5070 23154 5122
rect 24670 5070 24722 5122
rect 3278 4958 3330 5010
rect 6302 4958 6354 5010
rect 17390 4958 17442 5010
rect 18734 4958 18786 5010
rect 26574 4958 26626 5010
rect 31166 4958 31218 5010
rect 5070 4846 5122 4898
rect 7198 4846 7250 4898
rect 7982 4846 8034 4898
rect 8206 4846 8258 4898
rect 8766 4846 8818 4898
rect 14142 4846 14194 4898
rect 20750 4846 20802 4898
rect 21422 4846 21474 4898
rect 25790 4846 25842 4898
rect 9026 4678 9078 4730
rect 9130 4678 9182 4730
rect 9234 4678 9286 4730
rect 16838 4678 16890 4730
rect 16942 4678 16994 4730
rect 17046 4678 17098 4730
rect 24650 4678 24702 4730
rect 24754 4678 24806 4730
rect 24858 4678 24910 4730
rect 32462 4678 32514 4730
rect 32566 4678 32618 4730
rect 32670 4678 32722 4730
rect 5518 4510 5570 4562
rect 8430 4510 8482 4562
rect 8990 4510 9042 4562
rect 11902 4510 11954 4562
rect 12350 4510 12402 4562
rect 15486 4510 15538 4562
rect 17726 4510 17778 4562
rect 18062 4510 18114 4562
rect 20302 4510 20354 4562
rect 21422 4510 21474 4562
rect 23102 4510 23154 4562
rect 26014 4510 26066 4562
rect 26798 4510 26850 4562
rect 28142 4510 28194 4562
rect 28702 4510 28754 4562
rect 2382 4398 2434 4450
rect 7758 4398 7810 4450
rect 10110 4398 10162 4450
rect 16270 4398 16322 4450
rect 16830 4398 16882 4450
rect 19406 4398 19458 4450
rect 22766 4398 22818 4450
rect 25566 4398 25618 4450
rect 32174 4398 32226 4450
rect 4734 4286 4786 4338
rect 5294 4286 5346 4338
rect 5854 4286 5906 4338
rect 12798 4286 12850 4338
rect 13246 4286 13298 4338
rect 16606 4286 16658 4338
rect 20190 4286 20242 4338
rect 21310 4286 21362 4338
rect 23550 4286 23602 4338
rect 25230 4286 25282 4338
rect 26238 4286 26290 4338
rect 27918 4286 27970 4338
rect 31166 4286 31218 4338
rect 31614 4286 31666 4338
rect 6526 4174 6578 4226
rect 11118 4174 11170 4226
rect 18398 4174 18450 4226
rect 24670 4174 24722 4226
rect 27358 4174 27410 4226
rect 1598 4062 1650 4114
rect 24222 4062 24274 4114
rect 5120 3894 5172 3946
rect 5224 3894 5276 3946
rect 5328 3894 5380 3946
rect 12932 3894 12984 3946
rect 13036 3894 13088 3946
rect 13140 3894 13192 3946
rect 20744 3894 20796 3946
rect 20848 3894 20900 3946
rect 20952 3894 21004 3946
rect 28556 3894 28608 3946
rect 28660 3894 28712 3946
rect 28764 3894 28816 3946
rect 20862 3726 20914 3778
rect 27694 3726 27746 3778
rect 3838 3614 3890 3666
rect 4622 3614 4674 3666
rect 5070 3614 5122 3666
rect 5742 3614 5794 3666
rect 6302 3614 6354 3666
rect 6638 3614 6690 3666
rect 11006 3614 11058 3666
rect 14030 3614 14082 3666
rect 14590 3614 14642 3666
rect 14814 3614 14866 3666
rect 17166 3614 17218 3666
rect 17726 3614 17778 3666
rect 18174 3614 18226 3666
rect 23438 3614 23490 3666
rect 24110 3614 24162 3666
rect 26014 3614 26066 3666
rect 29934 3614 29986 3666
rect 30158 3614 30210 3666
rect 1822 3502 1874 3554
rect 12126 3502 12178 3554
rect 13358 3502 13410 3554
rect 19854 3502 19906 3554
rect 21086 3502 21138 3554
rect 22206 3502 22258 3554
rect 22766 3502 22818 3554
rect 25118 3502 25170 3554
rect 25566 3502 25618 3554
rect 27470 3502 27522 3554
rect 28590 3502 28642 3554
rect 2046 3390 2098 3442
rect 2606 3390 2658 3442
rect 7534 3390 7586 3442
rect 8318 3390 8370 3442
rect 8654 3390 8706 3442
rect 9998 3390 10050 3442
rect 13134 3390 13186 3442
rect 15822 3390 15874 3442
rect 18958 3390 19010 3442
rect 20190 3390 20242 3442
rect 22430 3390 22482 3442
rect 28366 3390 28418 3442
rect 31166 3390 31218 3442
rect 12350 3278 12402 3330
rect 24558 3278 24610 3330
rect 9026 3110 9078 3162
rect 9130 3110 9182 3162
rect 9234 3110 9286 3162
rect 16838 3110 16890 3162
rect 16942 3110 16994 3162
rect 17046 3110 17098 3162
rect 24650 3110 24702 3162
rect 24754 3110 24806 3162
rect 24858 3110 24910 3162
rect 32462 3110 32514 3162
rect 32566 3110 32618 3162
rect 32670 3110 32722 3162
<< metal2 >>
rect 672 33200 784 34000
rect 1344 33200 1456 34000
rect 2016 33200 2128 34000
rect 2688 33200 2800 34000
rect 3360 33200 3472 34000
rect 4032 33200 4144 34000
rect 4704 33200 4816 34000
rect 5376 33200 5488 34000
rect 6048 33200 6160 34000
rect 6720 33200 6832 34000
rect 7392 33200 7504 34000
rect 8064 33200 8176 34000
rect 8736 33200 8848 34000
rect 9408 33200 9520 34000
rect 10080 33200 10192 34000
rect 10752 33200 10864 34000
rect 11424 33200 11536 34000
rect 12096 33200 12208 34000
rect 12768 33200 12880 34000
rect 13440 33200 13552 34000
rect 14112 33200 14224 34000
rect 14784 33200 14896 34000
rect 15456 33200 15568 34000
rect 16128 33200 16240 34000
rect 16800 33200 16912 34000
rect 17472 33200 17584 34000
rect 18144 33200 18256 34000
rect 18816 33200 18928 34000
rect 24864 33200 24976 34000
rect 25536 33200 25648 34000
rect 26208 33200 26320 34000
rect 26880 33200 26992 34000
rect 27552 33200 27664 34000
rect 28224 33200 28336 34000
rect 28896 33200 29008 34000
rect 700 31948 756 33200
rect 700 31892 868 31948
rect 140 28756 196 28766
rect 140 18228 196 28700
rect 812 25172 868 31892
rect 1372 28868 1428 33200
rect 1820 32900 1876 32910
rect 1820 29650 1876 32844
rect 2044 31948 2100 33200
rect 2044 31892 2436 31948
rect 2156 30996 2212 31006
rect 2044 30324 2100 30334
rect 1820 29598 1822 29650
rect 1874 29598 1876 29650
rect 1820 29586 1876 29598
rect 1932 29986 1988 29998
rect 1932 29934 1934 29986
rect 1986 29934 1988 29986
rect 1932 29428 1988 29934
rect 1932 29362 1988 29372
rect 1372 28802 1428 28812
rect 2044 28642 2100 30268
rect 2156 30210 2212 30940
rect 2156 30158 2158 30210
rect 2210 30158 2212 30210
rect 2156 30146 2212 30158
rect 2044 28590 2046 28642
rect 2098 28590 2100 28642
rect 2044 28578 2100 28590
rect 2268 29540 2324 29550
rect 2268 28530 2324 29484
rect 2268 28478 2270 28530
rect 2322 28478 2324 28530
rect 2268 28466 2324 28478
rect 2156 27972 2212 27982
rect 2156 27878 2212 27916
rect 2044 27188 2100 27198
rect 2044 27074 2100 27132
rect 2044 27022 2046 27074
rect 2098 27022 2100 27074
rect 2044 27010 2100 27022
rect 2268 27076 2324 27086
rect 2268 26962 2324 27020
rect 2268 26910 2270 26962
rect 2322 26910 2324 26962
rect 2268 26898 2324 26910
rect 2380 26908 2436 31892
rect 2604 29426 2660 29438
rect 2604 29374 2606 29426
rect 2658 29374 2660 29426
rect 2604 29316 2660 29374
rect 2604 29250 2660 29260
rect 2380 26852 2548 26908
rect 2380 26402 2436 26414
rect 2380 26350 2382 26402
rect 2434 26350 2436 26402
rect 2156 26290 2212 26302
rect 2156 26238 2158 26290
rect 2210 26238 2212 26290
rect 2156 26068 2212 26238
rect 2156 26002 2212 26012
rect 2380 25732 2436 26350
rect 2380 25666 2436 25676
rect 1932 25620 1988 25630
rect 1932 25526 1988 25564
rect 812 25106 868 25116
rect 2044 25060 2100 25070
rect 1932 24612 1988 24622
rect 1932 24518 1988 24556
rect 2044 24388 2100 25004
rect 1932 24332 2100 24388
rect 2156 24498 2212 24510
rect 2156 24446 2158 24498
rect 2210 24446 2212 24498
rect 1820 23268 1876 23278
rect 140 18162 196 18172
rect 1484 23266 1876 23268
rect 1484 23214 1822 23266
rect 1874 23214 1876 23266
rect 1484 23212 1876 23214
rect 1484 17108 1540 23212
rect 1820 23202 1876 23212
rect 1820 22932 1876 22942
rect 1708 21252 1764 21262
rect 1596 19796 1652 19806
rect 1596 19702 1652 19740
rect 1596 17108 1652 17118
rect 1484 17106 1652 17108
rect 1484 17054 1598 17106
rect 1650 17054 1652 17106
rect 1484 17052 1652 17054
rect 1596 17042 1652 17052
rect 1260 15876 1316 15886
rect 1260 6468 1316 15820
rect 1596 15090 1652 15102
rect 1596 15038 1598 15090
rect 1650 15038 1652 15090
rect 1596 14420 1652 15038
rect 1596 14354 1652 14364
rect 1596 13524 1652 13534
rect 1484 13522 1652 13524
rect 1484 13470 1598 13522
rect 1650 13470 1652 13522
rect 1484 13468 1652 13470
rect 1484 10052 1540 13468
rect 1596 13458 1652 13468
rect 1708 12964 1764 21196
rect 1820 15148 1876 22876
rect 1932 22484 1988 24332
rect 2044 24052 2100 24062
rect 2044 23938 2100 23996
rect 2044 23886 2046 23938
rect 2098 23886 2100 23938
rect 2044 23874 2100 23886
rect 2044 22484 2100 22494
rect 1932 22482 2100 22484
rect 1932 22430 2046 22482
rect 2098 22430 2100 22482
rect 1932 22428 2100 22430
rect 2044 22418 2100 22428
rect 2156 22484 2212 24446
rect 2268 23716 2324 23726
rect 2268 23714 2436 23716
rect 2268 23662 2270 23714
rect 2322 23662 2436 23714
rect 2268 23660 2436 23662
rect 2268 23650 2324 23660
rect 2156 22418 2212 22428
rect 2268 22596 2324 22606
rect 2268 22482 2324 22540
rect 2268 22430 2270 22482
rect 2322 22430 2324 22482
rect 2268 22418 2324 22430
rect 2156 22148 2212 22158
rect 2156 21700 2212 22092
rect 2156 21586 2212 21644
rect 2156 21534 2158 21586
rect 2210 21534 2212 21586
rect 2156 21522 2212 21534
rect 2268 22036 2324 22046
rect 2156 20916 2212 20926
rect 2044 20804 2100 20814
rect 2044 20710 2100 20748
rect 2044 19348 2100 19358
rect 2044 19236 2100 19292
rect 1932 19234 2100 19236
rect 1932 19182 2046 19234
rect 2098 19182 2100 19234
rect 1932 19180 2100 19182
rect 1932 18674 1988 19180
rect 2044 19170 2100 19180
rect 1932 18622 1934 18674
rect 1986 18622 1988 18674
rect 1932 17778 1988 18622
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 17714 1988 17726
rect 2044 19010 2100 19022
rect 2044 18958 2046 19010
rect 2098 18958 2100 19010
rect 1932 17556 1988 17566
rect 1932 16098 1988 17500
rect 1932 16046 1934 16098
rect 1986 16046 1988 16098
rect 1932 16034 1988 16046
rect 2044 15540 2100 18958
rect 2156 18674 2212 20860
rect 2268 20690 2324 21980
rect 2380 21924 2436 23660
rect 2492 22484 2548 26852
rect 2604 25284 2660 25294
rect 2604 22484 2660 25228
rect 2716 23548 2772 33200
rect 3388 31948 3444 33200
rect 3724 32340 3780 32350
rect 3388 31892 3556 31948
rect 3388 30212 3444 30222
rect 3388 30098 3444 30156
rect 3388 30046 3390 30098
rect 3442 30046 3444 30098
rect 3388 30034 3444 30046
rect 2940 29986 2996 29998
rect 2940 29934 2942 29986
rect 2994 29934 2996 29986
rect 2940 29764 2996 29934
rect 3276 29764 3332 29774
rect 2940 29708 3276 29764
rect 2940 29428 2996 29438
rect 2940 26740 2996 29372
rect 3052 29204 3108 29214
rect 3052 28530 3108 29148
rect 3052 28478 3054 28530
rect 3106 28478 3108 28530
rect 3052 28466 3108 28478
rect 3164 27860 3220 27870
rect 3164 27746 3220 27804
rect 3164 27694 3166 27746
rect 3218 27694 3220 27746
rect 3164 27682 3220 27694
rect 3052 27636 3108 27646
rect 3052 26962 3108 27580
rect 3052 26910 3054 26962
rect 3106 26910 3108 26962
rect 3052 26898 3108 26910
rect 2940 26684 3108 26740
rect 2940 25620 2996 25630
rect 2940 25506 2996 25564
rect 2940 25454 2942 25506
rect 2994 25454 2996 25506
rect 2940 25442 2996 25454
rect 2940 25284 2996 25294
rect 3052 25284 3108 26684
rect 3164 26404 3220 26414
rect 3164 26310 3220 26348
rect 2996 25228 3108 25284
rect 2940 25218 2996 25228
rect 2940 24722 2996 24734
rect 2940 24670 2942 24722
rect 2994 24670 2996 24722
rect 2940 24612 2996 24670
rect 2940 24546 2996 24556
rect 3052 24500 3108 24510
rect 3052 23826 3108 24444
rect 3052 23774 3054 23826
rect 3106 23774 3108 23826
rect 3052 23762 3108 23774
rect 2716 23492 2884 23548
rect 2828 22708 2884 23492
rect 3052 23042 3108 23054
rect 3052 22990 3054 23042
rect 3106 22990 3108 23042
rect 2828 22652 2996 22708
rect 2604 22428 2772 22484
rect 2492 22418 2548 22428
rect 2380 21868 2660 21924
rect 2380 21700 2436 21710
rect 2380 21698 2548 21700
rect 2380 21646 2382 21698
rect 2434 21646 2548 21698
rect 2380 21644 2548 21646
rect 2380 21634 2436 21644
rect 2268 20638 2270 20690
rect 2322 20638 2324 20690
rect 2268 20626 2324 20638
rect 2380 20132 2436 20142
rect 2380 20038 2436 20076
rect 2156 18622 2158 18674
rect 2210 18622 2212 18674
rect 2156 18610 2212 18622
rect 2268 17554 2324 17566
rect 2268 17502 2270 17554
rect 2322 17502 2324 17554
rect 2268 17106 2324 17502
rect 2268 17054 2270 17106
rect 2322 17054 2324 17106
rect 2268 17042 2324 17054
rect 2268 15876 2324 15886
rect 2268 15782 2324 15820
rect 2156 15540 2212 15550
rect 2044 15538 2212 15540
rect 2044 15486 2158 15538
rect 2210 15486 2212 15538
rect 2044 15484 2212 15486
rect 2156 15474 2212 15484
rect 1820 15092 2324 15148
rect 2268 14418 2324 15092
rect 2492 14532 2548 21644
rect 2604 21476 2660 21868
rect 2604 21410 2660 21420
rect 2716 21028 2772 22428
rect 2492 14466 2548 14476
rect 2604 20972 2772 21028
rect 2828 22258 2884 22270
rect 2828 22206 2830 22258
rect 2882 22206 2884 22258
rect 2268 14366 2270 14418
rect 2322 14366 2324 14418
rect 1708 12870 1764 12908
rect 1932 14306 1988 14318
rect 1932 14254 1934 14306
rect 1986 14254 1988 14306
rect 1484 9986 1540 9996
rect 1596 11954 1652 11966
rect 1596 11902 1598 11954
rect 1650 11902 1652 11954
rect 1596 8372 1652 11902
rect 1932 11620 1988 14254
rect 2044 13188 2100 13198
rect 2044 12850 2100 13132
rect 2268 13076 2324 14366
rect 2380 13972 2436 13982
rect 2380 13878 2436 13916
rect 2492 13076 2548 13086
rect 2268 13074 2548 13076
rect 2268 13022 2494 13074
rect 2546 13022 2548 13074
rect 2268 13020 2548 13022
rect 2492 13010 2548 13020
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 2044 12786 2100 12798
rect 2492 12404 2548 12414
rect 1820 11564 1988 11620
rect 2380 12290 2436 12302
rect 2380 12238 2382 12290
rect 2434 12238 2436 12290
rect 2380 11620 2436 12238
rect 1820 10724 1876 11564
rect 2380 11554 2436 11564
rect 2268 11508 2324 11518
rect 1932 11396 1988 11406
rect 1932 11302 1988 11340
rect 2268 11282 2324 11452
rect 2268 11230 2270 11282
rect 2322 11230 2324 11282
rect 2268 11218 2324 11230
rect 2492 11060 2548 12348
rect 2268 11004 2548 11060
rect 1820 10668 2100 10724
rect 1708 10612 1764 10622
rect 1708 10610 1876 10612
rect 1708 10558 1710 10610
rect 1762 10558 1876 10610
rect 1708 10556 1876 10558
rect 1708 10546 1764 10556
rect 1820 9604 1876 10556
rect 1820 9042 1876 9548
rect 1820 8990 1822 9042
rect 1874 8990 1876 9042
rect 1820 8978 1876 8990
rect 1932 10500 1988 10510
rect 1596 8306 1652 8316
rect 1820 8820 1876 8830
rect 1820 7698 1876 8764
rect 1932 8146 1988 10444
rect 2044 9826 2100 10668
rect 2044 9774 2046 9826
rect 2098 9774 2100 9826
rect 2044 9762 2100 9774
rect 2156 10610 2212 10622
rect 2156 10558 2158 10610
rect 2210 10558 2212 10610
rect 1932 8094 1934 8146
rect 1986 8094 1988 8146
rect 1932 8082 1988 8094
rect 2044 9380 2100 9390
rect 2044 7924 2100 9324
rect 1820 7646 1822 7698
rect 1874 7646 1876 7698
rect 1820 6690 1876 7646
rect 1820 6638 1822 6690
rect 1874 6638 1876 6690
rect 1820 6626 1876 6638
rect 1932 7868 2100 7924
rect 1260 6402 1316 6412
rect 1932 6356 1988 7868
rect 2044 7700 2100 7710
rect 2044 6578 2100 7644
rect 2044 6526 2046 6578
rect 2098 6526 2100 6578
rect 2044 6514 2100 6526
rect 1932 6300 2100 6356
rect 1820 6244 1876 6254
rect 1596 4114 1652 4126
rect 1596 4062 1598 4114
rect 1650 4062 1652 4114
rect 1596 3444 1652 4062
rect 1820 3554 1876 6188
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5460 1988 5742
rect 1932 5394 1988 5404
rect 1820 3502 1822 3554
rect 1874 3502 1876 3554
rect 1820 3490 1876 3502
rect 1596 3378 1652 3388
rect 2044 3442 2100 6300
rect 2156 5234 2212 10558
rect 2268 9714 2324 11004
rect 2604 10948 2660 20972
rect 2828 19908 2884 22206
rect 2828 19842 2884 19852
rect 2716 19796 2772 19806
rect 2716 19122 2772 19740
rect 2716 19070 2718 19122
rect 2770 19070 2772 19122
rect 2716 19058 2772 19070
rect 2940 18676 2996 22652
rect 3052 20916 3108 22990
rect 3164 21698 3220 21710
rect 3164 21646 3166 21698
rect 3218 21646 3220 21698
rect 3164 21588 3220 21646
rect 3164 21522 3220 21532
rect 3052 20860 3220 20916
rect 3052 20692 3108 20702
rect 3052 20598 3108 20636
rect 2940 18620 3108 18676
rect 2940 18452 2996 18462
rect 2940 18358 2996 18396
rect 3052 17892 3108 18620
rect 3052 17826 3108 17836
rect 3052 17556 3108 17566
rect 3052 17462 3108 17500
rect 2828 16884 2884 16894
rect 2716 14420 2772 14430
rect 2716 14326 2772 14364
rect 2604 10882 2660 10892
rect 2268 9662 2270 9714
rect 2322 9662 2324 9714
rect 2268 9650 2324 9662
rect 2716 10052 2772 10062
rect 2268 9044 2324 9054
rect 2268 9042 2436 9044
rect 2268 8990 2270 9042
rect 2322 8990 2436 9042
rect 2268 8988 2436 8990
rect 2268 8978 2324 8988
rect 2268 8146 2324 8158
rect 2268 8094 2270 8146
rect 2322 8094 2324 8146
rect 2268 5908 2324 8094
rect 2380 7364 2436 8988
rect 2716 8146 2772 9996
rect 2828 8820 2884 16828
rect 3052 15986 3108 15998
rect 3052 15934 3054 15986
rect 3106 15934 3108 15986
rect 3052 14756 3108 15934
rect 3164 15316 3220 20860
rect 3164 15250 3220 15260
rect 3052 14690 3108 14700
rect 3052 13524 3108 13534
rect 2940 12964 2996 12974
rect 2940 12870 2996 12908
rect 3052 11282 3108 13468
rect 3276 12404 3332 29708
rect 3388 25506 3444 25518
rect 3388 25454 3390 25506
rect 3442 25454 3444 25506
rect 3388 22036 3444 25454
rect 3500 24724 3556 31892
rect 3612 31668 3668 31678
rect 3612 29314 3668 31612
rect 3724 29428 3780 32284
rect 3836 29986 3892 29998
rect 3836 29934 3838 29986
rect 3890 29934 3892 29986
rect 3836 29764 3892 29934
rect 3836 29698 3892 29708
rect 3948 29652 4004 29662
rect 3724 29372 3892 29428
rect 3612 29262 3614 29314
rect 3666 29262 3668 29314
rect 3612 29250 3668 29262
rect 3724 25732 3780 25742
rect 3724 24946 3780 25676
rect 3836 25618 3892 29372
rect 3836 25566 3838 25618
rect 3890 25566 3892 25618
rect 3836 25554 3892 25566
rect 3724 24894 3726 24946
rect 3778 24894 3780 24946
rect 3724 24882 3780 24894
rect 3948 24948 4004 29596
rect 4060 29092 4116 33200
rect 4620 33012 4676 33022
rect 4172 29988 4228 29998
rect 4172 29894 4228 29932
rect 4172 29316 4228 29326
rect 4228 29260 4340 29316
rect 4172 29222 4228 29260
rect 4060 29026 4116 29036
rect 4060 28756 4116 28766
rect 4060 28662 4116 28700
rect 4172 28308 4228 28318
rect 4060 27186 4116 27198
rect 4060 27134 4062 27186
rect 4114 27134 4116 27186
rect 4060 26292 4116 27134
rect 4172 26516 4228 28252
rect 4284 27412 4340 29260
rect 4396 29204 4452 29214
rect 4396 29110 4452 29148
rect 4508 28420 4564 28430
rect 4620 28420 4676 32956
rect 4732 31948 4788 33200
rect 5404 31948 5460 33200
rect 4732 31892 4900 31948
rect 5404 31892 5908 31948
rect 4844 28644 4900 31892
rect 5118 30604 5382 30614
rect 5174 30548 5222 30604
rect 5278 30548 5326 30604
rect 5118 30538 5382 30548
rect 4956 30100 5012 30110
rect 4956 30006 5012 30044
rect 5628 30098 5684 30110
rect 5628 30046 5630 30098
rect 5682 30046 5684 30098
rect 5628 29876 5684 30046
rect 5628 29810 5684 29820
rect 5740 29764 5796 29774
rect 5180 29538 5236 29550
rect 5180 29486 5182 29538
rect 5234 29486 5236 29538
rect 5180 29204 5236 29486
rect 5180 29138 5236 29148
rect 5118 29036 5382 29046
rect 5174 28980 5222 29036
rect 5278 28980 5326 29036
rect 5118 28970 5382 28980
rect 4844 28578 4900 28588
rect 5628 28644 5684 28654
rect 4620 28364 5012 28420
rect 4396 27636 4452 27646
rect 4396 27542 4452 27580
rect 4284 27356 4452 27412
rect 4172 26450 4228 26460
rect 4060 26226 4116 26236
rect 4172 26178 4228 26190
rect 4172 26126 4174 26178
rect 4226 26126 4228 26178
rect 4172 25508 4228 26126
rect 4172 25442 4228 25452
rect 3948 24892 4340 24948
rect 3500 24658 3556 24668
rect 3724 24722 3780 24734
rect 3724 24670 3726 24722
rect 3778 24670 3780 24722
rect 3724 23940 3780 24670
rect 4172 24500 4228 24510
rect 4172 24406 4228 24444
rect 3724 23874 3780 23884
rect 3948 24276 4004 24286
rect 3388 21970 3444 21980
rect 3500 23604 3556 23614
rect 3500 16884 3556 23548
rect 3948 19796 4004 24220
rect 4060 24050 4116 24062
rect 4060 23998 4062 24050
rect 4114 23998 4116 24050
rect 4060 23156 4116 23998
rect 4060 23090 4116 23100
rect 4172 23940 4228 23950
rect 4172 23378 4228 23884
rect 4172 23326 4174 23378
rect 4226 23326 4228 23378
rect 4172 22596 4228 23326
rect 4060 22482 4116 22494
rect 4060 22430 4062 22482
rect 4114 22430 4116 22482
rect 4060 21588 4116 22430
rect 4172 22148 4228 22540
rect 4172 22082 4228 22092
rect 4060 21522 4116 21532
rect 4172 21474 4228 21486
rect 4172 21422 4174 21474
rect 4226 21422 4228 21474
rect 4060 20914 4116 20926
rect 4060 20862 4062 20914
rect 4114 20862 4116 20914
rect 4060 20020 4116 20862
rect 4172 20804 4228 21422
rect 4172 20738 4228 20748
rect 4060 19954 4116 19964
rect 3948 19740 4228 19796
rect 4060 19346 4116 19358
rect 4060 19294 4062 19346
rect 4114 19294 4116 19346
rect 4060 19236 4116 19294
rect 4060 19170 4116 19180
rect 3724 18452 3780 18462
rect 3724 18358 3780 18396
rect 4060 18450 4116 18462
rect 4060 18398 4062 18450
rect 4114 18398 4116 18450
rect 3948 17778 4004 17790
rect 3948 17726 3950 17778
rect 4002 17726 4004 17778
rect 3948 17668 4004 17726
rect 3948 17602 4004 17612
rect 3500 16818 3556 16828
rect 3948 16210 4004 16222
rect 3948 16158 3950 16210
rect 4002 16158 4004 16210
rect 3948 16100 4004 16158
rect 3948 16034 4004 16044
rect 4060 14642 4116 18398
rect 4060 14590 4062 14642
rect 4114 14590 4116 14642
rect 4060 14578 4116 14590
rect 3276 12338 3332 12348
rect 3724 14532 3780 14542
rect 3724 11508 3780 14476
rect 3836 13076 3892 13086
rect 3836 12982 3892 13020
rect 4060 12516 4116 12526
rect 3948 12460 4060 12516
rect 3836 11508 3892 11518
rect 3724 11506 3892 11508
rect 3724 11454 3838 11506
rect 3890 11454 3892 11506
rect 3724 11452 3892 11454
rect 3836 11442 3892 11452
rect 3052 11230 3054 11282
rect 3106 11230 3108 11282
rect 3052 11218 3108 11230
rect 3052 10388 3108 10398
rect 3052 9714 3108 10332
rect 3948 9938 4004 12460
rect 4060 12450 4116 12460
rect 4172 11396 4228 19740
rect 4284 12180 4340 24892
rect 4396 15148 4452 27356
rect 4508 27188 4564 28364
rect 4508 27094 4564 27132
rect 4732 26180 4788 26190
rect 4620 26178 4788 26180
rect 4620 26126 4734 26178
rect 4786 26126 4788 26178
rect 4620 26124 4788 26126
rect 4620 25284 4676 26124
rect 4732 26114 4788 26124
rect 4732 25620 4788 25630
rect 4732 25526 4788 25564
rect 4956 25394 5012 28364
rect 5180 27972 5236 27982
rect 5180 27970 5572 27972
rect 5180 27918 5182 27970
rect 5234 27918 5572 27970
rect 5180 27916 5572 27918
rect 5180 27906 5236 27916
rect 5118 27468 5382 27478
rect 5174 27412 5222 27468
rect 5278 27412 5326 27468
rect 5118 27402 5382 27412
rect 5068 26180 5124 26190
rect 5068 26086 5124 26124
rect 5118 25900 5382 25910
rect 5174 25844 5222 25900
rect 5278 25844 5326 25900
rect 5118 25834 5382 25844
rect 5516 25732 5572 27916
rect 5628 26290 5684 28588
rect 5740 28530 5796 29708
rect 5740 28478 5742 28530
rect 5794 28478 5796 28530
rect 5740 28466 5796 28478
rect 5740 28308 5796 28318
rect 5740 26850 5796 28252
rect 5740 26798 5742 26850
rect 5794 26798 5796 26850
rect 5740 26786 5796 26798
rect 5628 26238 5630 26290
rect 5682 26238 5684 26290
rect 5628 26226 5684 26238
rect 5852 25732 5908 31892
rect 5964 30098 6020 30110
rect 5964 30046 5966 30098
rect 6018 30046 6020 30098
rect 5964 28084 6020 30046
rect 5964 28018 6020 28028
rect 6076 27748 6132 33200
rect 6636 30436 6692 30446
rect 6412 29986 6468 29998
rect 6412 29934 6414 29986
rect 6466 29934 6468 29986
rect 6412 29876 6468 29934
rect 6188 29204 6244 29214
rect 6244 29148 6356 29204
rect 6188 29138 6244 29148
rect 6188 28644 6244 28654
rect 6188 28550 6244 28588
rect 6076 27682 6132 27692
rect 5964 26292 6020 26302
rect 5964 26198 6020 26236
rect 6076 25732 6132 25742
rect 5852 25730 6132 25732
rect 5852 25678 6078 25730
rect 6130 25678 6132 25730
rect 5852 25676 6132 25678
rect 5516 25666 5572 25676
rect 6076 25666 6132 25676
rect 4956 25342 4958 25394
rect 5010 25342 5012 25394
rect 4956 25330 5012 25342
rect 4620 25218 4676 25228
rect 5740 25284 5796 25294
rect 5740 25190 5796 25228
rect 6300 25060 6356 29148
rect 6300 24994 6356 25004
rect 6412 25284 6468 29820
rect 6524 26964 6580 26974
rect 6524 26870 6580 26908
rect 4956 24836 5012 24846
rect 4956 24742 5012 24780
rect 5964 24836 6020 24846
rect 5118 24332 5382 24342
rect 5174 24276 5222 24332
rect 5278 24276 5326 24332
rect 5118 24266 5382 24276
rect 4508 24052 4564 24062
rect 4508 23958 4564 23996
rect 5964 24050 6020 24780
rect 5964 23998 5966 24050
rect 6018 23998 6020 24050
rect 5964 23986 6020 23998
rect 6300 24052 6356 24062
rect 6412 24052 6468 25228
rect 6300 24050 6468 24052
rect 6300 23998 6302 24050
rect 6354 23998 6468 24050
rect 6300 23996 6468 23998
rect 5068 23940 5124 23950
rect 5068 23846 5124 23884
rect 6300 23940 6356 23996
rect 6300 23874 6356 23884
rect 4620 23154 4676 23166
rect 4620 23102 4622 23154
rect 4674 23102 4676 23154
rect 4620 22484 4676 23102
rect 4956 23156 5012 23166
rect 4956 23062 5012 23100
rect 5118 22764 5382 22774
rect 5174 22708 5222 22764
rect 5278 22708 5326 22764
rect 5118 22698 5382 22708
rect 4620 22418 4676 22428
rect 5068 22484 5124 22494
rect 5068 22390 5124 22428
rect 5628 22484 5684 22494
rect 4620 22148 4676 22158
rect 4620 22054 4676 22092
rect 4956 22148 5012 22158
rect 4620 21700 4676 21710
rect 4620 21606 4676 21644
rect 4620 21028 4676 21038
rect 4620 20578 4676 20972
rect 4620 20526 4622 20578
rect 4674 20526 4676 20578
rect 4508 19348 4564 19358
rect 4508 19254 4564 19292
rect 4508 17892 4564 17902
rect 4508 17778 4564 17836
rect 4508 17726 4510 17778
rect 4562 17726 4564 17778
rect 4508 17714 4564 17726
rect 4620 15652 4676 20526
rect 4732 20916 4788 20926
rect 4732 20018 4788 20860
rect 4956 20244 5012 22092
rect 5628 21586 5684 22428
rect 5628 21534 5630 21586
rect 5682 21534 5684 21586
rect 5118 21196 5382 21206
rect 5174 21140 5222 21196
rect 5278 21140 5326 21196
rect 5118 21130 5382 21140
rect 4956 20178 5012 20188
rect 5628 20916 5684 21534
rect 5852 22258 5908 22270
rect 5852 22206 5854 22258
rect 5906 22206 5908 22258
rect 5740 20916 5796 20926
rect 5628 20914 5796 20916
rect 5628 20862 5742 20914
rect 5794 20862 5796 20914
rect 5628 20860 5796 20862
rect 4732 19966 4734 20018
rect 4786 19966 4788 20018
rect 4732 19954 4788 19966
rect 5292 20020 5348 20030
rect 5628 20020 5684 20860
rect 5740 20850 5796 20860
rect 5852 20132 5908 22206
rect 6188 22258 6244 22270
rect 6188 22206 6190 22258
rect 6242 22206 6244 22258
rect 5964 21588 6020 21598
rect 5964 21494 6020 21532
rect 6188 20580 6244 22206
rect 6524 22148 6580 22158
rect 6524 22054 6580 22092
rect 6412 20580 6468 20590
rect 6188 20578 6468 20580
rect 6188 20526 6414 20578
rect 6466 20526 6468 20578
rect 6188 20524 6468 20526
rect 5852 20066 5908 20076
rect 5292 20018 5684 20020
rect 5292 19966 5294 20018
rect 5346 19966 5630 20018
rect 5682 19966 5684 20018
rect 5292 19964 5684 19966
rect 5292 19954 5348 19964
rect 5118 19628 5382 19638
rect 5174 19572 5222 19628
rect 5278 19572 5326 19628
rect 5118 19562 5382 19572
rect 5628 19234 5684 19964
rect 5964 20020 6020 20030
rect 5964 19926 6020 19964
rect 6412 19348 6468 20524
rect 6412 19282 6468 19292
rect 5628 19182 5630 19234
rect 5682 19182 5684 19234
rect 5628 18452 5684 19182
rect 6076 19236 6132 19246
rect 6076 19142 6132 19180
rect 6412 18564 6468 18574
rect 4956 18340 5012 18350
rect 4956 18116 5012 18284
rect 4956 18050 5012 18060
rect 5118 18060 5382 18070
rect 5174 18004 5222 18060
rect 5278 18004 5326 18060
rect 5118 17994 5382 18004
rect 5068 17780 5124 17790
rect 5628 17780 5684 18396
rect 6300 18562 6468 18564
rect 6300 18510 6414 18562
rect 6466 18510 6468 18562
rect 6300 18508 6468 18510
rect 5740 17780 5796 17790
rect 5068 17778 5796 17780
rect 5068 17726 5070 17778
rect 5122 17726 5742 17778
rect 5794 17726 5796 17778
rect 5068 17724 5796 17726
rect 5068 17714 5124 17724
rect 4732 16884 4788 16894
rect 4732 16882 4900 16884
rect 4732 16830 4734 16882
rect 4786 16830 4900 16882
rect 4732 16828 4900 16830
rect 4732 16818 4788 16828
rect 4732 16212 4788 16222
rect 4732 16118 4788 16156
rect 4620 15596 4788 15652
rect 4620 15316 4676 15326
rect 4620 15222 4676 15260
rect 4396 15092 4564 15148
rect 4396 14644 4452 14654
rect 4396 14084 4452 14588
rect 4396 14018 4452 14028
rect 4508 13860 4564 15092
rect 4732 14644 4788 15596
rect 4732 14578 4788 14588
rect 4620 14308 4676 14318
rect 4620 14214 4676 14252
rect 4396 13804 4564 13860
rect 4396 12404 4452 13804
rect 4620 13748 4676 13758
rect 4508 13746 4676 13748
rect 4508 13694 4622 13746
rect 4674 13694 4676 13746
rect 4508 13692 4676 13694
rect 4508 13076 4564 13692
rect 4620 13682 4676 13692
rect 4508 13010 4564 13020
rect 4732 13636 4788 13646
rect 4396 12338 4452 12348
rect 4284 12124 4564 12180
rect 4172 11330 4228 11340
rect 4508 11506 4564 12124
rect 4508 11454 4510 11506
rect 4562 11454 4564 11506
rect 4508 11284 4564 11454
rect 4508 11218 4564 11228
rect 4620 12178 4676 12190
rect 4620 12126 4622 12178
rect 4674 12126 4676 12178
rect 4620 10724 4676 12126
rect 4732 10834 4788 13580
rect 4844 13076 4900 16828
rect 5292 16882 5348 17724
rect 5740 17714 5796 17724
rect 5404 17556 5460 17566
rect 5404 17106 5460 17500
rect 5404 17054 5406 17106
rect 5458 17054 5460 17106
rect 5404 17042 5460 17054
rect 6188 16996 6244 17006
rect 6188 16902 6244 16940
rect 5292 16830 5294 16882
rect 5346 16830 5348 16882
rect 5292 16818 5348 16830
rect 6076 16772 6132 16782
rect 5118 16492 5382 16502
rect 5174 16436 5222 16492
rect 5278 16436 5326 16492
rect 5118 16426 5382 16436
rect 5068 16212 5124 16222
rect 5068 16118 5124 16156
rect 5964 16212 6020 16222
rect 5964 16098 6020 16156
rect 5964 16046 5966 16098
rect 6018 16046 6020 16098
rect 5964 16034 6020 16046
rect 5740 15874 5796 15886
rect 5740 15822 5742 15874
rect 5794 15822 5796 15874
rect 5068 15314 5124 15326
rect 5068 15262 5070 15314
rect 5122 15262 5124 15314
rect 5068 15148 5124 15262
rect 5628 15316 5684 15326
rect 5628 15148 5684 15260
rect 4956 15092 5124 15148
rect 5516 15092 5684 15148
rect 4956 14308 5012 15092
rect 5118 14924 5382 14934
rect 5174 14868 5222 14924
rect 5278 14868 5326 14924
rect 5118 14858 5382 14868
rect 5516 14756 5572 15092
rect 5180 14700 5572 14756
rect 5628 14756 5684 14766
rect 5180 14642 5236 14700
rect 5180 14590 5182 14642
rect 5234 14590 5236 14642
rect 5180 14578 5236 14590
rect 5516 14532 5572 14542
rect 5628 14532 5684 14700
rect 5516 14530 5684 14532
rect 5516 14478 5518 14530
rect 5570 14478 5684 14530
rect 5516 14476 5684 14478
rect 5516 14466 5572 14476
rect 4956 13748 5012 14252
rect 5740 13972 5796 15822
rect 5964 15316 6020 15326
rect 5964 15222 6020 15260
rect 5740 13906 5796 13916
rect 5404 13860 5460 13870
rect 5404 13766 5460 13804
rect 5292 13748 5348 13758
rect 4956 13746 5348 13748
rect 4956 13694 5294 13746
rect 5346 13694 5348 13746
rect 4956 13692 5348 13694
rect 4956 13188 5012 13692
rect 5292 13524 5348 13692
rect 5292 13458 5348 13468
rect 5118 13356 5382 13366
rect 5174 13300 5222 13356
rect 5278 13300 5326 13356
rect 5118 13290 5382 13300
rect 4956 13132 5124 13188
rect 4844 13010 4900 13020
rect 4956 12852 5012 12862
rect 4956 12758 5012 12796
rect 5068 12178 5124 13132
rect 5964 12962 6020 12974
rect 5964 12910 5966 12962
rect 6018 12910 6020 12962
rect 5516 12404 5572 12414
rect 5516 12310 5572 12348
rect 5068 12126 5070 12178
rect 5122 12126 5124 12178
rect 5068 11956 5124 12126
rect 5740 12180 5796 12190
rect 5740 12178 5908 12180
rect 5740 12126 5742 12178
rect 5794 12126 5908 12178
rect 5740 12124 5908 12126
rect 5740 12114 5796 12124
rect 4956 11900 5124 11956
rect 4956 11620 5012 11900
rect 5118 11788 5382 11798
rect 5174 11732 5222 11788
rect 5278 11732 5326 11788
rect 5118 11722 5382 11732
rect 5740 11620 5796 11630
rect 4956 11564 5124 11620
rect 4732 10782 4734 10834
rect 4786 10782 4788 10834
rect 4732 10770 4788 10782
rect 5068 11506 5124 11564
rect 5740 11526 5796 11564
rect 5068 11454 5070 11506
rect 5122 11454 5124 11506
rect 3948 9886 3950 9938
rect 4002 9886 4004 9938
rect 3948 9874 4004 9886
rect 4060 10668 4676 10724
rect 3052 9662 3054 9714
rect 3106 9662 3108 9714
rect 3052 9650 3108 9662
rect 3836 9716 3892 9726
rect 2828 8754 2884 8764
rect 2716 8094 2718 8146
rect 2770 8094 2772 8146
rect 2716 8082 2772 8094
rect 3276 8372 3332 8382
rect 2716 7364 2772 7374
rect 2380 7362 2772 7364
rect 2380 7310 2718 7362
rect 2770 7310 2772 7362
rect 2380 7308 2772 7310
rect 2716 7298 2772 7308
rect 3052 6578 3108 6590
rect 3052 6526 3054 6578
rect 3106 6526 3108 6578
rect 3052 6356 3108 6526
rect 3052 6290 3108 6300
rect 2268 5842 2324 5852
rect 2940 5906 2996 5918
rect 2940 5854 2942 5906
rect 2994 5854 2996 5906
rect 2940 5348 2996 5854
rect 2940 5282 2996 5292
rect 2156 5182 2158 5234
rect 2210 5182 2212 5234
rect 2156 5170 2212 5182
rect 3276 5010 3332 8316
rect 3500 7364 3556 7374
rect 3388 6692 3444 6702
rect 3388 5906 3444 6636
rect 3388 5854 3390 5906
rect 3442 5854 3444 5906
rect 3388 5796 3444 5854
rect 3388 5730 3444 5740
rect 3276 4958 3278 5010
rect 3330 4958 3332 5010
rect 3276 4946 3332 4958
rect 2380 4450 2436 4462
rect 2380 4398 2382 4450
rect 2434 4398 2436 4450
rect 2380 3780 2436 4398
rect 2380 3714 2436 3724
rect 2044 3390 2046 3442
rect 2098 3390 2100 3442
rect 2044 3378 2100 3390
rect 2604 3444 2660 3482
rect 2604 3378 2660 3388
rect 3500 2100 3556 7308
rect 3836 6804 3892 9660
rect 3948 9268 4004 9278
rect 3948 7586 4004 9212
rect 4060 8370 4116 10668
rect 4508 10500 4564 10510
rect 4508 9266 4564 10444
rect 5068 10388 5124 11454
rect 4956 10332 5124 10388
rect 5292 10388 5348 10426
rect 4956 10052 5012 10332
rect 5292 10322 5348 10332
rect 5404 10388 5460 10398
rect 5404 10386 5572 10388
rect 5404 10334 5406 10386
rect 5458 10334 5572 10386
rect 5404 10332 5572 10334
rect 5404 10322 5460 10332
rect 5118 10220 5382 10230
rect 5174 10164 5222 10220
rect 5278 10164 5326 10220
rect 5118 10154 5382 10164
rect 4620 9996 5460 10052
rect 4620 9938 4676 9996
rect 4620 9886 4622 9938
rect 4674 9886 4676 9938
rect 4620 9604 4676 9886
rect 4620 9538 4676 9548
rect 4508 9214 4510 9266
rect 4562 9214 4564 9266
rect 4508 9202 4564 9214
rect 4956 8372 5012 9996
rect 5068 9604 5124 9614
rect 5068 9510 5124 9548
rect 5404 9042 5460 9996
rect 5516 9268 5572 10332
rect 5852 9380 5908 12124
rect 5964 11394 6020 12910
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 10724 6020 11342
rect 5964 9604 6020 10668
rect 5964 9538 6020 9548
rect 5852 9314 5908 9324
rect 6076 9268 6132 16716
rect 6188 15428 6244 15438
rect 6300 15428 6356 18508
rect 6412 18498 6468 18508
rect 6636 18340 6692 30380
rect 6748 29988 6804 33200
rect 7420 31948 7476 33200
rect 8092 31948 8148 33200
rect 7420 31892 7700 31948
rect 7420 30322 7476 30334
rect 7420 30270 7422 30322
rect 7474 30270 7476 30322
rect 6748 29922 6804 29932
rect 6972 30100 7028 30110
rect 6972 29988 7028 30044
rect 6972 29986 7252 29988
rect 6972 29934 6974 29986
rect 7026 29934 7252 29986
rect 6972 29932 7252 29934
rect 6972 29922 7028 29932
rect 6860 29316 6916 29326
rect 6860 28754 6916 29260
rect 6860 28702 6862 28754
rect 6914 28702 6916 28754
rect 6860 28690 6916 28702
rect 7196 26908 7252 29932
rect 7420 29426 7476 30270
rect 7644 29652 7700 31892
rect 7644 29586 7700 29596
rect 7980 31892 8148 31948
rect 7420 29374 7422 29426
rect 7474 29374 7476 29426
rect 7420 29362 7476 29374
rect 7308 28980 7364 28990
rect 7308 28642 7364 28924
rect 7308 28590 7310 28642
rect 7362 28590 7364 28642
rect 7308 28578 7364 28590
rect 7420 28756 7476 28766
rect 7420 27858 7476 28700
rect 7420 27806 7422 27858
rect 7474 27806 7476 27858
rect 7420 27794 7476 27806
rect 7756 28530 7812 28542
rect 7756 28478 7758 28530
rect 7810 28478 7812 28530
rect 7532 27188 7588 27198
rect 7532 27094 7588 27132
rect 7196 26852 7588 26908
rect 6860 25620 6916 25630
rect 6860 25282 6916 25564
rect 6860 25230 6862 25282
rect 6914 25230 6916 25282
rect 6860 21812 6916 25230
rect 7420 25394 7476 25406
rect 7420 25342 7422 25394
rect 7474 25342 7476 25394
rect 7308 24836 7364 24846
rect 7308 24722 7364 24780
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 24658 7364 24670
rect 7084 23826 7140 23838
rect 7084 23774 7086 23826
rect 7138 23774 7140 23826
rect 7084 22148 7140 23774
rect 7420 23378 7476 25342
rect 7420 23326 7422 23378
rect 7474 23326 7476 23378
rect 7420 23314 7476 23326
rect 7084 22082 7140 22092
rect 6860 21756 7140 21812
rect 6860 20916 6916 20926
rect 6860 20822 6916 20860
rect 6412 18284 6692 18340
rect 6412 17778 6468 18284
rect 6412 17726 6414 17778
rect 6466 17726 6468 17778
rect 6412 17714 6468 17726
rect 6972 17780 7028 17790
rect 6860 17444 6916 17454
rect 6748 17442 6916 17444
rect 6748 17390 6862 17442
rect 6914 17390 6916 17442
rect 6748 17388 6916 17390
rect 6188 15426 6356 15428
rect 6188 15374 6190 15426
rect 6242 15374 6356 15426
rect 6188 15372 6356 15374
rect 6412 15876 6468 15886
rect 6188 15362 6244 15372
rect 6412 15148 6468 15820
rect 6636 15428 6692 15438
rect 6636 15334 6692 15372
rect 6300 15092 6468 15148
rect 6300 14418 6356 15092
rect 6300 14366 6302 14418
rect 6354 14366 6356 14418
rect 6300 14354 6356 14366
rect 6188 13858 6244 13870
rect 6188 13806 6190 13858
rect 6242 13806 6244 13858
rect 6188 13074 6244 13806
rect 6188 13022 6190 13074
rect 6242 13022 6244 13074
rect 6188 13010 6244 13022
rect 6748 12964 6804 17388
rect 6860 17378 6916 17388
rect 6972 16210 7028 17724
rect 7084 16884 7140 21756
rect 7420 18450 7476 18462
rect 7420 18398 7422 18450
rect 7474 18398 7476 18450
rect 7084 16818 7140 16828
rect 7196 18226 7252 18238
rect 7196 18174 7198 18226
rect 7250 18174 7252 18226
rect 7196 16324 7252 18174
rect 7420 18004 7476 18398
rect 7420 17938 7476 17948
rect 7420 17780 7476 17818
rect 7420 17714 7476 17724
rect 6972 16158 6974 16210
rect 7026 16158 7028 16210
rect 6972 16146 7028 16158
rect 7084 16268 7252 16324
rect 7084 15988 7140 16268
rect 7420 16212 7476 16222
rect 7420 16100 7476 16156
rect 6748 12898 6804 12908
rect 6860 15932 7140 15988
rect 7196 16098 7476 16100
rect 7196 16046 7422 16098
rect 7474 16046 7476 16098
rect 7196 16044 7476 16046
rect 6860 12290 6916 15932
rect 7196 15148 7252 16044
rect 7420 16034 7476 16044
rect 7308 15876 7364 15886
rect 7308 15782 7364 15820
rect 6972 15092 7252 15148
rect 6972 13074 7028 15092
rect 6972 13022 6974 13074
rect 7026 13022 7028 13074
rect 6972 13010 7028 13022
rect 7420 13412 7476 13422
rect 7420 12738 7476 13356
rect 7420 12686 7422 12738
rect 7474 12686 7476 12738
rect 7420 12404 7476 12686
rect 7420 12338 7476 12348
rect 6860 12238 6862 12290
rect 6914 12238 6916 12290
rect 6860 12226 6916 12238
rect 7532 12292 7588 26852
rect 7756 25620 7812 28478
rect 7980 28308 8036 31892
rect 8652 30436 8708 30446
rect 8540 30380 8652 30436
rect 7980 28242 8036 28252
rect 8092 29426 8148 29438
rect 8092 29374 8094 29426
rect 8146 29374 8148 29426
rect 8092 28644 8148 29374
rect 8092 27858 8148 28588
rect 8540 27972 8596 30380
rect 8652 30370 8708 30380
rect 8652 30098 8708 30110
rect 8652 30046 8654 30098
rect 8706 30046 8708 30098
rect 8652 29988 8708 30046
rect 8652 29922 8708 29932
rect 8764 29764 8820 33200
rect 9436 31948 9492 33200
rect 9324 31892 9492 31948
rect 9324 30212 9380 31892
rect 9324 30146 9380 30156
rect 9436 30324 9492 30334
rect 9436 30098 9492 30268
rect 9436 30046 9438 30098
rect 9490 30046 9492 30098
rect 9436 30034 9492 30046
rect 9772 30100 9828 30110
rect 9772 30006 9828 30044
rect 9996 29876 10052 29886
rect 9024 29820 9288 29830
rect 9080 29764 9128 29820
rect 9184 29764 9232 29820
rect 9024 29754 9288 29764
rect 8764 29698 8820 29708
rect 9548 29652 9604 29662
rect 9548 29558 9604 29596
rect 8764 29540 8820 29550
rect 8764 29426 8820 29484
rect 8764 29374 8766 29426
rect 8818 29374 8820 29426
rect 8764 29362 8820 29374
rect 8988 29538 9044 29550
rect 8988 29486 8990 29538
rect 9042 29486 9044 29538
rect 8988 29092 9044 29486
rect 9996 29540 10052 29820
rect 10108 29652 10164 33200
rect 10780 31948 10836 33200
rect 11452 31948 11508 33200
rect 10668 31892 10836 31948
rect 11228 31892 11508 31948
rect 10556 30098 10612 30110
rect 10556 30046 10558 30098
rect 10610 30046 10612 30098
rect 10108 29596 10276 29652
rect 9548 29316 9604 29326
rect 8988 29036 9492 29092
rect 9324 28868 9380 28878
rect 9100 28866 9380 28868
rect 9100 28814 9326 28866
rect 9378 28814 9380 28866
rect 9100 28812 9380 28814
rect 9100 28754 9156 28812
rect 9324 28802 9380 28812
rect 9100 28702 9102 28754
rect 9154 28702 9156 28754
rect 9100 28690 9156 28702
rect 8988 28532 9044 28542
rect 8876 28476 8988 28532
rect 8876 28084 8932 28476
rect 8988 28466 9044 28476
rect 9024 28252 9288 28262
rect 9080 28196 9128 28252
rect 9184 28196 9232 28252
rect 9024 28186 9288 28196
rect 8988 28084 9044 28094
rect 8876 28082 9044 28084
rect 8876 28030 8990 28082
rect 9042 28030 9044 28082
rect 8876 28028 9044 28030
rect 8988 28018 9044 28028
rect 8652 27972 8708 27982
rect 8540 27970 8708 27972
rect 8540 27918 8654 27970
rect 8706 27918 8708 27970
rect 8540 27916 8708 27918
rect 8652 27906 8708 27916
rect 8764 27972 8820 27982
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 7980 27188 8036 27198
rect 8092 27188 8148 27806
rect 8764 27298 8820 27916
rect 8764 27246 8766 27298
rect 8818 27246 8820 27298
rect 8764 27234 8820 27246
rect 7980 27186 8148 27188
rect 7980 27134 7982 27186
rect 8034 27134 8148 27186
rect 7980 27132 8148 27134
rect 7980 25956 8036 27132
rect 8540 26850 8596 26862
rect 8540 26798 8542 26850
rect 8594 26798 8596 26850
rect 8316 26402 8372 26414
rect 8316 26350 8318 26402
rect 8370 26350 8372 26402
rect 7980 25900 8260 25956
rect 8092 25620 8148 25630
rect 7756 25618 8148 25620
rect 7756 25566 8094 25618
rect 8146 25566 8148 25618
rect 7756 25564 8148 25566
rect 8092 25554 8148 25564
rect 7756 25394 7812 25406
rect 7756 25342 7758 25394
rect 7810 25342 7812 25394
rect 7756 25284 7812 25342
rect 7756 25218 7812 25228
rect 8092 25172 8148 25182
rect 7756 24948 7812 24958
rect 7756 24722 7812 24892
rect 8092 24946 8148 25116
rect 8092 24894 8094 24946
rect 8146 24894 8148 24946
rect 8092 24882 8148 24894
rect 8204 24948 8260 25900
rect 8204 24882 8260 24892
rect 7756 24670 7758 24722
rect 7810 24670 7812 24722
rect 7756 24658 7812 24670
rect 8092 24050 8148 24062
rect 8092 23998 8094 24050
rect 8146 23998 8148 24050
rect 8092 23156 8148 23998
rect 8316 23716 8372 26350
rect 8540 25172 8596 26798
rect 9024 26684 9288 26694
rect 9080 26628 9128 26684
rect 9184 26628 9232 26684
rect 9024 26618 9288 26628
rect 9100 26404 9156 26414
rect 9100 26310 9156 26348
rect 8540 24724 8596 25116
rect 8876 25282 8932 25294
rect 8876 25230 8878 25282
rect 8930 25230 8932 25282
rect 8540 24658 8596 24668
rect 8652 24948 8708 24958
rect 8652 24052 8708 24892
rect 8876 24946 8932 25230
rect 9024 25116 9288 25126
rect 9080 25060 9128 25116
rect 9184 25060 9232 25116
rect 9024 25050 9288 25060
rect 8876 24894 8878 24946
rect 8930 24894 8932 24946
rect 8876 24882 8932 24894
rect 8988 24724 9044 24734
rect 8988 24630 9044 24668
rect 8316 23650 8372 23660
rect 8540 24050 8708 24052
rect 8540 23998 8654 24050
rect 8706 23998 8708 24050
rect 8540 23996 8708 23998
rect 8092 23090 8148 23100
rect 8428 23042 8484 23054
rect 8428 22990 8430 23042
rect 8482 22990 8484 23042
rect 8092 22930 8148 22942
rect 8092 22878 8094 22930
rect 8146 22878 8148 22930
rect 8092 20692 8148 22878
rect 8092 20626 8148 20636
rect 8204 20690 8260 20702
rect 8204 20638 8206 20690
rect 8258 20638 8260 20690
rect 8204 19796 8260 20638
rect 8428 20242 8484 22990
rect 8540 22484 8596 23996
rect 8652 23986 8708 23996
rect 9100 23828 9156 23838
rect 9100 23716 9156 23772
rect 8652 23714 9156 23716
rect 8652 23662 9102 23714
rect 9154 23662 9156 23714
rect 8652 23660 9156 23662
rect 8652 23266 8708 23660
rect 9100 23650 9156 23660
rect 9024 23548 9288 23558
rect 9080 23492 9128 23548
rect 9184 23492 9232 23548
rect 9024 23482 9288 23492
rect 9436 23492 9492 29036
rect 9548 28756 9604 29260
rect 9996 29204 10052 29484
rect 10108 29428 10164 29438
rect 10108 29334 10164 29372
rect 10220 29204 10276 29596
rect 9996 29148 10164 29204
rect 9548 28662 9604 28700
rect 9996 28866 10052 28878
rect 9996 28814 9998 28866
rect 10050 28814 10052 28866
rect 9548 28084 9604 28094
rect 9548 26962 9604 28028
rect 9548 26910 9550 26962
rect 9602 26910 9604 26962
rect 9548 26898 9604 26910
rect 9660 27858 9716 27870
rect 9660 27806 9662 27858
rect 9714 27806 9716 27858
rect 9660 24164 9716 27806
rect 9772 27076 9828 27086
rect 9772 26908 9828 27020
rect 9772 26852 9940 26908
rect 9884 26402 9940 26852
rect 9884 26350 9886 26402
rect 9938 26350 9940 26402
rect 9884 26338 9940 26350
rect 9884 24724 9940 24734
rect 9772 24612 9828 24622
rect 9772 24518 9828 24556
rect 9548 23940 9604 23950
rect 9660 23940 9716 24108
rect 9548 23938 9716 23940
rect 9548 23886 9550 23938
rect 9602 23886 9716 23938
rect 9548 23884 9716 23886
rect 9548 23874 9604 23884
rect 9436 23426 9492 23436
rect 9548 23716 9604 23726
rect 8652 23214 8654 23266
rect 8706 23214 8708 23266
rect 8652 23202 8708 23214
rect 9548 23266 9604 23660
rect 9660 23604 9716 23614
rect 9716 23548 9828 23604
rect 9660 23538 9716 23548
rect 9548 23214 9550 23266
rect 9602 23214 9604 23266
rect 9548 23202 9604 23214
rect 8540 22390 8596 22428
rect 9024 21980 9288 21990
rect 9080 21924 9128 21980
rect 9184 21924 9232 21980
rect 9024 21914 9288 21924
rect 8540 21810 8596 21822
rect 8540 21758 8542 21810
rect 8594 21758 8596 21810
rect 8540 21588 8596 21758
rect 8540 21522 8596 21532
rect 8764 21700 8820 21710
rect 8764 20802 8820 21644
rect 9100 21586 9156 21598
rect 9100 21534 9102 21586
rect 9154 21534 9156 21586
rect 9100 21476 9156 21534
rect 9548 21588 9604 21598
rect 9548 21494 9604 21532
rect 9100 21410 9156 21420
rect 8764 20750 8766 20802
rect 8818 20750 8820 20802
rect 8764 20738 8820 20750
rect 9100 20804 9156 20814
rect 9100 20710 9156 20748
rect 9024 20412 9288 20422
rect 9080 20356 9128 20412
rect 9184 20356 9232 20412
rect 9024 20346 9288 20356
rect 8428 20190 8430 20242
rect 8482 20190 8484 20242
rect 8428 20178 8484 20190
rect 9660 20132 9716 20142
rect 9436 20130 9716 20132
rect 9436 20078 9662 20130
rect 9714 20078 9716 20130
rect 9436 20076 9716 20078
rect 9100 19908 9156 19918
rect 9100 19814 9156 19852
rect 8204 19730 8260 19740
rect 8652 19010 8708 19022
rect 9212 19012 9268 19022
rect 8652 18958 8654 19010
rect 8706 18958 8708 19010
rect 7644 18452 7700 18462
rect 7644 17780 7700 18396
rect 7868 18340 7924 18350
rect 7868 18246 7924 18284
rect 7644 17666 7700 17724
rect 7644 17614 7646 17666
rect 7698 17614 7700 17666
rect 7644 17602 7700 17614
rect 7756 18004 7812 18014
rect 7756 16772 7812 17948
rect 8204 17668 8260 17678
rect 8204 17574 8260 17612
rect 8652 17108 8708 18958
rect 8652 17042 8708 17052
rect 8764 19010 9268 19012
rect 8764 18958 9214 19010
rect 9266 18958 9268 19010
rect 8764 18956 9268 18958
rect 7756 16706 7812 16716
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 8204 15874 8260 15886
rect 8204 15822 8206 15874
rect 8258 15822 8260 15874
rect 8204 15428 8260 15822
rect 8204 15362 8260 15372
rect 7980 15202 8036 15214
rect 7980 15150 7982 15202
rect 8034 15150 8036 15202
rect 7980 14868 8036 15150
rect 8428 15148 8484 16830
rect 8540 15316 8596 15326
rect 8540 15222 8596 15260
rect 7980 14802 8036 14812
rect 8204 15092 8484 15148
rect 8092 13076 8148 13086
rect 8092 12982 8148 13020
rect 7532 12226 7588 12236
rect 7980 12068 8036 12078
rect 8204 12068 8260 15092
rect 8652 14980 8708 14990
rect 8540 14532 8596 14542
rect 8540 14438 8596 14476
rect 8428 13746 8484 13758
rect 8428 13694 8430 13746
rect 8482 13694 8484 13746
rect 8428 12516 8484 13694
rect 8652 13636 8708 14924
rect 8652 13570 8708 13580
rect 8764 12852 8820 18956
rect 9212 18946 9268 18956
rect 9024 18844 9288 18854
rect 9080 18788 9128 18844
rect 9184 18788 9232 18844
rect 9024 18778 9288 18788
rect 9436 18674 9492 20076
rect 9660 20066 9716 20076
rect 9772 19908 9828 23548
rect 9884 23266 9940 24668
rect 9996 23938 10052 28814
rect 10108 28754 10164 29148
rect 10220 29138 10276 29148
rect 10108 28702 10110 28754
rect 10162 28702 10164 28754
rect 10108 28690 10164 28702
rect 10332 28980 10388 28990
rect 10108 27860 10164 27870
rect 10108 27766 10164 27804
rect 10220 26964 10276 26974
rect 10220 26514 10276 26908
rect 10332 26908 10388 28924
rect 10556 28868 10612 30046
rect 10556 28802 10612 28812
rect 10332 26852 10500 26908
rect 10220 26462 10222 26514
rect 10274 26462 10276 26514
rect 10220 26450 10276 26462
rect 10220 24724 10276 24734
rect 10220 24722 10388 24724
rect 10220 24670 10222 24722
rect 10274 24670 10388 24722
rect 10220 24668 10388 24670
rect 10220 24658 10276 24668
rect 9996 23886 9998 23938
rect 10050 23886 10052 23938
rect 9996 23874 10052 23886
rect 10220 24164 10276 24174
rect 10108 23828 10164 23838
rect 10108 23604 10164 23772
rect 9884 23214 9886 23266
rect 9938 23214 9940 23266
rect 9884 23202 9940 23214
rect 9996 23548 10164 23604
rect 9884 21700 9940 21710
rect 9996 21700 10052 23548
rect 10220 23154 10276 24108
rect 10332 23604 10388 24668
rect 10332 23538 10388 23548
rect 10220 23102 10222 23154
rect 10274 23102 10276 23154
rect 10220 23090 10276 23102
rect 10332 21812 10388 21822
rect 10444 21812 10500 26852
rect 10668 24052 10724 31892
rect 10780 29652 10836 29662
rect 10780 29558 10836 29596
rect 11004 26402 11060 26414
rect 11004 26350 11006 26402
rect 11058 26350 11060 26402
rect 10780 25060 10836 25070
rect 10780 24946 10836 25004
rect 10780 24894 10782 24946
rect 10834 24894 10836 24946
rect 10780 24724 10836 24894
rect 10780 24658 10836 24668
rect 11004 24612 11060 26350
rect 11116 25508 11172 25518
rect 11116 25414 11172 25452
rect 11004 24546 11060 24556
rect 10668 23986 10724 23996
rect 10780 23156 10836 23166
rect 10780 23062 10836 23100
rect 10332 21810 10500 21812
rect 10332 21758 10334 21810
rect 10386 21758 10500 21810
rect 10332 21756 10500 21758
rect 10332 21746 10388 21756
rect 9884 21698 10052 21700
rect 9884 21646 9886 21698
rect 9938 21646 10052 21698
rect 9884 21644 10052 21646
rect 9884 21634 9940 21644
rect 10556 21588 10612 21598
rect 10556 21494 10612 21532
rect 9436 18622 9438 18674
rect 9490 18622 9492 18674
rect 9436 18610 9492 18622
rect 9548 19852 9828 19908
rect 10892 21028 10948 21038
rect 8988 18452 9044 18462
rect 8876 18396 8988 18452
rect 8876 16882 8932 18396
rect 8988 18358 9044 18396
rect 9024 17276 9288 17286
rect 9080 17220 9128 17276
rect 9184 17220 9232 17276
rect 9024 17210 9288 17220
rect 9548 17108 9604 19852
rect 9772 19348 9828 19358
rect 9772 19254 9828 19292
rect 10892 19122 10948 20972
rect 10892 19070 10894 19122
rect 10946 19070 10948 19122
rect 10892 19058 10948 19070
rect 11004 19906 11060 19918
rect 11004 19854 11006 19906
rect 11058 19854 11060 19906
rect 9884 19010 9940 19022
rect 9884 18958 9886 19010
rect 9938 18958 9940 19010
rect 9884 17556 9940 18958
rect 10220 18562 10276 18574
rect 10220 18510 10222 18562
rect 10274 18510 10276 18562
rect 10220 17780 10276 18510
rect 11004 18228 11060 19854
rect 11228 19348 11284 31892
rect 11564 30322 11620 30334
rect 11564 30270 11566 30322
rect 11618 30270 11620 30322
rect 11340 29316 11396 29326
rect 11340 29222 11396 29260
rect 11340 28756 11396 28766
rect 11340 25284 11396 28700
rect 11564 28644 11620 30270
rect 11900 30324 11956 30334
rect 11564 28578 11620 28588
rect 11676 28754 11732 28766
rect 11676 28702 11678 28754
rect 11730 28702 11732 28754
rect 11676 25732 11732 28702
rect 11788 27636 11844 27646
rect 11788 27076 11844 27580
rect 11788 27010 11844 27020
rect 11900 27074 11956 30268
rect 12012 30100 12068 30110
rect 12012 30006 12068 30044
rect 12012 29540 12068 29550
rect 12012 29446 12068 29484
rect 12124 28196 12180 33200
rect 12796 31948 12852 33200
rect 12684 31892 12852 31948
rect 12684 28420 12740 31892
rect 12930 30604 13194 30614
rect 12986 30548 13034 30604
rect 13090 30548 13138 30604
rect 12930 30538 13194 30548
rect 13244 30436 13300 30446
rect 13244 30098 13300 30380
rect 13244 30046 13246 30098
rect 13298 30046 13300 30098
rect 13244 30034 13300 30046
rect 13468 29876 13524 33200
rect 14140 31948 14196 33200
rect 14140 31892 14756 31948
rect 13580 30212 13636 30222
rect 13580 30118 13636 30156
rect 14028 30212 14084 30222
rect 14028 30118 14084 30156
rect 13468 29810 13524 29820
rect 13020 29316 13076 29326
rect 13020 29222 13076 29260
rect 12930 29036 13194 29046
rect 12986 28980 13034 29036
rect 13090 28980 13138 29036
rect 12930 28970 13194 28980
rect 13468 28644 13524 28654
rect 13356 28642 13524 28644
rect 13356 28590 13470 28642
rect 13522 28590 13524 28642
rect 13356 28588 13524 28590
rect 12684 28354 12740 28364
rect 12796 28530 12852 28542
rect 12796 28478 12798 28530
rect 12850 28478 12852 28530
rect 12124 28130 12180 28140
rect 12572 28084 12628 28094
rect 12572 27990 12628 28028
rect 12236 27748 12292 27758
rect 12292 27692 12404 27748
rect 12236 27682 12292 27692
rect 11900 27022 11902 27074
rect 11954 27022 11956 27074
rect 11900 27010 11956 27022
rect 12348 26908 12404 27692
rect 12460 27076 12516 27086
rect 12460 26982 12516 27020
rect 12348 26852 12740 26908
rect 12684 26850 12740 26852
rect 12684 26798 12686 26850
rect 12738 26798 12740 26850
rect 12684 26786 12740 26798
rect 11788 26516 11844 26526
rect 11788 25844 11844 26460
rect 11900 26178 11956 26190
rect 11900 26126 11902 26178
rect 11954 26126 11956 26178
rect 11900 25956 11956 26126
rect 12460 26178 12516 26190
rect 12460 26126 12462 26178
rect 12514 26126 12516 26178
rect 11900 25900 12292 25956
rect 11788 25788 12068 25844
rect 11676 25676 11956 25732
rect 11788 25508 11844 25518
rect 11788 25284 11844 25452
rect 11340 25218 11396 25228
rect 11676 25228 11844 25284
rect 11676 24948 11732 25228
rect 11676 24882 11732 24892
rect 11564 24724 11620 24734
rect 11900 24724 11956 25676
rect 12012 25394 12068 25788
rect 12012 25342 12014 25394
rect 12066 25342 12068 25394
rect 12012 25330 12068 25342
rect 12124 24724 12180 24734
rect 11900 24722 12180 24724
rect 11900 24670 12126 24722
rect 12178 24670 12180 24722
rect 11900 24668 12180 24670
rect 11340 24610 11396 24622
rect 11340 24558 11342 24610
rect 11394 24558 11396 24610
rect 11340 23828 11396 24558
rect 11564 24164 11620 24668
rect 12124 24658 12180 24668
rect 11620 24108 11732 24164
rect 11564 24098 11620 24108
rect 11340 23762 11396 23772
rect 11564 22370 11620 22382
rect 11564 22318 11566 22370
rect 11618 22318 11620 22370
rect 11452 22260 11508 22270
rect 11452 20690 11508 22204
rect 11564 21812 11620 22318
rect 11564 21746 11620 21756
rect 11676 21700 11732 24108
rect 12236 23940 12292 25900
rect 12460 25508 12516 26126
rect 12460 25442 12516 25452
rect 12572 25618 12628 25630
rect 12796 25620 12852 28478
rect 13356 27858 13412 28588
rect 13468 28578 13524 28588
rect 13916 28644 13972 28654
rect 13916 28550 13972 28588
rect 13356 27806 13358 27858
rect 13410 27806 13412 27858
rect 13132 27636 13188 27674
rect 13132 27570 13188 27580
rect 12930 27468 13194 27478
rect 12986 27412 13034 27468
rect 13090 27412 13138 27468
rect 12930 27402 13194 27412
rect 13356 27076 13412 27806
rect 13692 28084 13748 28094
rect 13692 27186 13748 28028
rect 13692 27134 13694 27186
rect 13746 27134 13748 27186
rect 13692 27122 13748 27134
rect 13804 27858 13860 27870
rect 13804 27806 13806 27858
rect 13858 27806 13860 27858
rect 13804 27188 13860 27806
rect 13804 27122 13860 27132
rect 13916 27748 13972 27758
rect 13020 26292 13076 26302
rect 13020 26198 13076 26236
rect 13356 26290 13412 27020
rect 13356 26238 13358 26290
rect 13410 26238 13412 26290
rect 12930 25900 13194 25910
rect 12986 25844 13034 25900
rect 13090 25844 13138 25900
rect 12930 25834 13194 25844
rect 12572 25566 12574 25618
rect 12626 25566 12628 25618
rect 12236 23874 12292 23884
rect 12460 23716 12516 23726
rect 12572 23716 12628 25566
rect 12684 25564 12852 25620
rect 12908 25732 12964 25742
rect 12684 24388 12740 25564
rect 12796 25396 12852 25406
rect 12908 25396 12964 25676
rect 12796 25394 12964 25396
rect 12796 25342 12798 25394
rect 12850 25342 12964 25394
rect 12796 25340 12964 25342
rect 12796 25060 12852 25340
rect 12796 24994 12852 25004
rect 13244 24724 13300 24734
rect 13356 24724 13412 26238
rect 13916 26290 13972 27692
rect 14700 27188 14756 31892
rect 14812 29652 14868 33200
rect 14924 30324 14980 30334
rect 14924 30230 14980 30268
rect 15484 30100 15540 33200
rect 16156 30212 16212 33200
rect 16156 30146 16212 30156
rect 15484 30034 15540 30044
rect 16268 30098 16324 30110
rect 16268 30046 16270 30098
rect 16322 30046 16324 30098
rect 14812 29586 14868 29596
rect 15372 29314 15428 29326
rect 15372 29262 15374 29314
rect 15426 29262 15428 29314
rect 14812 27188 14868 27198
rect 14700 27186 14868 27188
rect 14700 27134 14814 27186
rect 14866 27134 14868 27186
rect 14700 27132 14868 27134
rect 14812 27122 14868 27132
rect 13916 26238 13918 26290
rect 13970 26238 13972 26290
rect 13916 26226 13972 26238
rect 14028 27076 14084 27086
rect 14028 26962 14084 27020
rect 14028 26910 14030 26962
rect 14082 26910 14084 26962
rect 14028 26292 14084 26910
rect 14364 26964 14420 26974
rect 15372 26908 15428 29262
rect 16268 29204 16324 30046
rect 16828 30100 16884 33200
rect 16828 30044 17444 30100
rect 16836 29820 17100 29830
rect 16892 29764 16940 29820
rect 16996 29764 17044 29820
rect 16836 29754 17100 29764
rect 17388 29652 17444 30044
rect 17500 29876 17556 33200
rect 17500 29810 17556 29820
rect 17948 30322 18004 30334
rect 17948 30270 17950 30322
rect 18002 30270 18004 30322
rect 17388 29596 17892 29652
rect 16604 29540 16660 29550
rect 17052 29540 17108 29550
rect 16604 29538 16772 29540
rect 16604 29486 16606 29538
rect 16658 29486 16772 29538
rect 16604 29484 16772 29486
rect 16604 29474 16660 29484
rect 16268 29138 16324 29148
rect 16604 28644 16660 28654
rect 16492 28420 16548 28430
rect 16492 28326 16548 28364
rect 15932 28196 15988 28206
rect 15596 27076 15652 27086
rect 15596 26982 15652 27020
rect 14364 26870 14420 26908
rect 13692 26180 13748 26190
rect 13300 24668 13524 24724
rect 13244 24658 13300 24668
rect 12684 24332 12852 24388
rect 12796 24164 12852 24332
rect 12930 24332 13194 24342
rect 12986 24276 13034 24332
rect 13090 24276 13138 24332
rect 12930 24266 13194 24276
rect 13020 24164 13076 24174
rect 12796 24162 13076 24164
rect 12796 24110 13022 24162
rect 13074 24110 13076 24162
rect 12796 24108 13076 24110
rect 13020 24098 13076 24108
rect 13468 23938 13524 24668
rect 13468 23886 13470 23938
rect 13522 23886 13524 23938
rect 13468 23874 13524 23886
rect 12460 23714 12628 23716
rect 12460 23662 12462 23714
rect 12514 23662 12628 23714
rect 12460 23660 12628 23662
rect 12796 23828 12852 23838
rect 12460 23650 12516 23660
rect 12796 22372 12852 23772
rect 13356 23378 13412 23390
rect 13356 23326 13358 23378
rect 13410 23326 13412 23378
rect 12930 22764 13194 22774
rect 12986 22708 13034 22764
rect 13090 22708 13138 22764
rect 12930 22698 13194 22708
rect 12796 22278 12852 22316
rect 12572 22260 12628 22270
rect 12572 22166 12628 22204
rect 12236 22148 12292 22158
rect 11788 21700 11844 21710
rect 11732 21698 12180 21700
rect 11732 21646 11790 21698
rect 11842 21646 12180 21698
rect 11732 21644 12180 21646
rect 11676 21606 11732 21644
rect 11788 21634 11844 21644
rect 11452 20638 11454 20690
rect 11506 20638 11508 20690
rect 11452 20626 11508 20638
rect 12012 20804 12068 20814
rect 12012 20130 12068 20748
rect 12012 20078 12014 20130
rect 12066 20078 12068 20130
rect 12012 20066 12068 20078
rect 12124 20020 12180 21644
rect 12236 21026 12292 22092
rect 12460 21812 12516 21822
rect 12236 20974 12238 21026
rect 12290 20974 12292 21026
rect 12236 20962 12292 20974
rect 12348 21756 12460 21812
rect 12236 20020 12292 20030
rect 12124 20018 12292 20020
rect 12124 19966 12238 20018
rect 12290 19966 12292 20018
rect 12124 19964 12292 19966
rect 11228 19282 11284 19292
rect 11452 19906 11508 19918
rect 11452 19854 11454 19906
rect 11506 19854 11508 19906
rect 11452 19236 11508 19854
rect 12236 19458 12292 19964
rect 12236 19406 12238 19458
rect 12290 19406 12292 19458
rect 12236 19394 12292 19406
rect 11900 19346 11956 19358
rect 11900 19294 11902 19346
rect 11954 19294 11956 19346
rect 11508 19180 11620 19236
rect 11452 19170 11508 19180
rect 11004 18162 11060 18172
rect 11452 18452 11508 18462
rect 10220 17714 10276 17724
rect 10556 17556 10612 17566
rect 9884 17554 10612 17556
rect 9884 17502 10558 17554
rect 10610 17502 10612 17554
rect 9884 17500 10612 17502
rect 10556 17490 10612 17500
rect 11340 17444 11396 17454
rect 10780 17442 11396 17444
rect 10780 17390 11342 17442
rect 11394 17390 11396 17442
rect 10780 17388 11396 17390
rect 8876 16830 8878 16882
rect 8930 16830 8932 16882
rect 8876 16818 8932 16830
rect 9436 17052 9604 17108
rect 10668 17108 10724 17118
rect 8988 15876 9044 15914
rect 8988 15810 9044 15820
rect 9024 15708 9288 15718
rect 9080 15652 9128 15708
rect 9184 15652 9232 15708
rect 9024 15642 9288 15652
rect 8988 15540 9044 15550
rect 8988 15446 9044 15484
rect 9436 15148 9492 17052
rect 10668 16994 10724 17052
rect 10668 16942 10670 16994
rect 10722 16942 10724 16994
rect 10668 16930 10724 16942
rect 9772 16882 9828 16894
rect 9772 16830 9774 16882
rect 9826 16830 9828 16882
rect 9660 16658 9716 16670
rect 9660 16606 9662 16658
rect 9714 16606 9716 16658
rect 9436 15092 9604 15148
rect 9436 14756 9492 14766
rect 9548 14756 9604 15092
rect 9660 14980 9716 16606
rect 9772 16212 9828 16830
rect 9772 15540 9828 16156
rect 10332 16884 10388 16894
rect 9772 15314 9828 15484
rect 9884 15876 9940 15886
rect 9884 15538 9940 15820
rect 9884 15486 9886 15538
rect 9938 15486 9940 15538
rect 9884 15474 9940 15486
rect 9772 15262 9774 15314
rect 9826 15262 9828 15314
rect 9772 15148 9828 15262
rect 9772 15092 10164 15148
rect 9660 14914 9716 14924
rect 9884 14868 9940 14878
rect 9548 14700 9828 14756
rect 9212 14532 9268 14542
rect 8876 14476 9212 14532
rect 8876 13746 8932 14476
rect 9212 14438 9268 14476
rect 9024 14140 9288 14150
rect 9080 14084 9128 14140
rect 9184 14084 9232 14140
rect 9024 14074 9288 14084
rect 9436 13860 9492 14700
rect 9548 14532 9604 14542
rect 9548 14530 9716 14532
rect 9548 14478 9550 14530
rect 9602 14478 9716 14530
rect 9548 14476 9716 14478
rect 9548 14466 9604 14476
rect 9548 13860 9604 13870
rect 9436 13858 9604 13860
rect 9436 13806 9550 13858
rect 9602 13806 9604 13858
rect 9436 13804 9604 13806
rect 9548 13794 9604 13804
rect 8876 13694 8878 13746
rect 8930 13694 8932 13746
rect 8876 13682 8932 13694
rect 9100 12852 9156 12862
rect 8764 12850 9156 12852
rect 8764 12798 9102 12850
rect 9154 12798 9156 12850
rect 8764 12796 9156 12798
rect 9100 12786 9156 12796
rect 9024 12572 9288 12582
rect 9080 12516 9128 12572
rect 9184 12516 9232 12572
rect 9024 12506 9288 12516
rect 8428 12450 8484 12460
rect 8988 12404 9044 12414
rect 7980 12066 8260 12068
rect 7980 12014 7982 12066
rect 8034 12014 8260 12066
rect 7980 12012 8260 12014
rect 8876 12348 8988 12404
rect 7980 12002 8036 12012
rect 6188 11956 6244 11966
rect 6188 10834 6244 11900
rect 6188 10782 6190 10834
rect 6242 10782 6244 10834
rect 6188 10770 6244 10782
rect 6748 11170 6804 11182
rect 6748 11118 6750 11170
rect 6802 11118 6804 11170
rect 6636 10724 6692 10734
rect 6636 9826 6692 10668
rect 6636 9774 6638 9826
rect 6690 9774 6692 9826
rect 6636 9762 6692 9774
rect 6636 9604 6692 9614
rect 6636 9510 6692 9548
rect 5516 9202 5572 9212
rect 5964 9212 6132 9268
rect 5404 8990 5406 9042
rect 5458 8990 5460 9042
rect 5404 8978 5460 8990
rect 5292 8820 5348 8830
rect 5292 8818 5796 8820
rect 5292 8766 5294 8818
rect 5346 8766 5796 8818
rect 5292 8764 5796 8766
rect 5292 8754 5348 8764
rect 5118 8652 5382 8662
rect 5174 8596 5222 8652
rect 5278 8596 5326 8652
rect 5118 8586 5382 8596
rect 5068 8372 5124 8382
rect 4060 8318 4062 8370
rect 4114 8318 4116 8370
rect 4060 8306 4116 8318
rect 4620 8370 5572 8372
rect 4620 8318 5070 8370
rect 5122 8318 5572 8370
rect 4620 8316 5572 8318
rect 3948 7534 3950 7586
rect 4002 7534 4004 7586
rect 3948 7522 4004 7534
rect 4620 7474 4676 8316
rect 4620 7422 4622 7474
rect 4674 7422 4676 7474
rect 4620 7410 4676 7422
rect 4620 6916 4676 6926
rect 3836 6738 3892 6748
rect 4060 6802 4116 6814
rect 4060 6750 4062 6802
rect 4114 6750 4116 6802
rect 4060 6692 4116 6750
rect 4060 6626 4116 6636
rect 3612 6580 3668 6590
rect 3612 6130 3668 6524
rect 4508 6466 4564 6478
rect 4508 6414 4510 6466
rect 4562 6414 4564 6466
rect 3612 6078 3614 6130
rect 3666 6078 3668 6130
rect 3612 6066 3668 6078
rect 4060 6356 4116 6366
rect 4060 6130 4116 6300
rect 4508 6244 4564 6414
rect 4508 6178 4564 6188
rect 4060 6078 4062 6130
rect 4114 6078 4116 6130
rect 4060 6066 4116 6078
rect 3948 5796 4004 5806
rect 3836 5684 3892 5694
rect 3836 3666 3892 5628
rect 3948 5234 4004 5740
rect 3948 5182 3950 5234
rect 4002 5182 4004 5234
rect 3948 5170 4004 5182
rect 3836 3614 3838 3666
rect 3890 3614 3892 3666
rect 3836 3602 3892 3614
rect 4172 4116 4228 4126
rect 4172 3332 4228 4060
rect 4620 3892 4676 6860
rect 4956 6804 5012 8316
rect 5068 8306 5124 8316
rect 5516 8258 5572 8316
rect 5516 8206 5518 8258
rect 5570 8206 5572 8258
rect 5516 8194 5572 8206
rect 5068 7474 5124 7486
rect 5068 7422 5070 7474
rect 5122 7422 5124 7474
rect 5068 7252 5124 7422
rect 5404 7252 5460 7262
rect 5068 7196 5404 7252
rect 5404 7186 5460 7196
rect 5118 7084 5382 7094
rect 5174 7028 5222 7084
rect 5278 7028 5326 7084
rect 5118 7018 5382 7028
rect 5068 6804 5124 6814
rect 4956 6748 5068 6804
rect 5068 6710 5124 6748
rect 5404 6804 5460 6814
rect 5460 6748 5572 6804
rect 5404 6738 5460 6748
rect 4844 6018 4900 6030
rect 4844 5966 4846 6018
rect 4898 5966 4900 6018
rect 4844 5796 4900 5966
rect 4732 5740 4844 5796
rect 4732 5234 4788 5740
rect 4844 5730 4900 5740
rect 5118 5516 5382 5526
rect 5174 5460 5222 5516
rect 5278 5460 5326 5516
rect 5118 5450 5382 5460
rect 5516 5348 5572 6748
rect 5628 6580 5684 6590
rect 5628 6486 5684 6524
rect 4732 5182 4734 5234
rect 4786 5182 4788 5234
rect 4732 5170 4788 5182
rect 5292 5292 5572 5348
rect 5628 5908 5684 5918
rect 5068 4900 5124 4910
rect 5068 4806 5124 4844
rect 4732 4564 4788 4574
rect 4732 4338 4788 4508
rect 4732 4286 4734 4338
rect 4786 4286 4788 4338
rect 4732 4274 4788 4286
rect 5292 4340 5348 5292
rect 5516 4564 5572 4574
rect 5628 4564 5684 5852
rect 5740 4788 5796 8764
rect 5964 6578 6020 9212
rect 6076 9042 6132 9054
rect 6076 8990 6078 9042
rect 6130 8990 6132 9042
rect 6076 8820 6132 8990
rect 6076 8764 6580 8820
rect 5964 6526 5966 6578
rect 6018 6526 6020 6578
rect 5964 6514 6020 6526
rect 6076 8258 6132 8270
rect 6076 8206 6078 8258
rect 6130 8206 6132 8258
rect 6076 5684 6132 8206
rect 6300 6804 6356 6814
rect 6300 6690 6356 6748
rect 6300 6638 6302 6690
rect 6354 6638 6356 6690
rect 6300 6626 6356 6638
rect 6076 5618 6132 5628
rect 6412 5460 6468 5470
rect 6412 5122 6468 5404
rect 6412 5070 6414 5122
rect 6466 5070 6468 5122
rect 6300 5012 6356 5022
rect 6300 4918 6356 4956
rect 5740 4722 5796 4732
rect 5516 4562 5684 4564
rect 5516 4510 5518 4562
rect 5570 4510 5684 4562
rect 5516 4508 5684 4510
rect 5516 4498 5572 4508
rect 5740 4452 5796 4462
rect 5796 4396 5908 4452
rect 5740 4386 5796 4396
rect 5292 4338 5684 4340
rect 5292 4286 5294 4338
rect 5346 4286 5684 4338
rect 5292 4284 5684 4286
rect 5292 4274 5348 4284
rect 4508 3836 4676 3892
rect 5118 3948 5382 3958
rect 5174 3892 5222 3948
rect 5278 3892 5326 3948
rect 5118 3882 5382 3892
rect 4508 3556 4564 3836
rect 5068 3780 5124 3790
rect 4620 3668 4676 3678
rect 4620 3574 4676 3612
rect 5068 3666 5124 3724
rect 5068 3614 5070 3666
rect 5122 3614 5124 3666
rect 5068 3602 5124 3614
rect 5628 3668 5684 4284
rect 5852 4338 5908 4396
rect 5852 4286 5854 4338
rect 5906 4286 5908 4338
rect 5852 4274 5908 4286
rect 5740 3668 5796 3678
rect 5628 3666 5796 3668
rect 5628 3614 5742 3666
rect 5794 3614 5796 3666
rect 5628 3612 5796 3614
rect 5740 3602 5796 3612
rect 6300 3668 6356 3678
rect 6412 3668 6468 5070
rect 6524 4226 6580 8764
rect 6748 7364 6804 11118
rect 7308 11170 7364 11182
rect 7308 11118 7310 11170
rect 7362 11118 7364 11170
rect 7308 10724 7364 11118
rect 8428 10836 8484 10846
rect 8316 10724 8372 10734
rect 7308 10658 7364 10668
rect 8204 10668 8316 10724
rect 6748 7298 6804 7308
rect 7420 7698 7476 7710
rect 7420 7646 7422 7698
rect 7474 7646 7476 7698
rect 6524 4174 6526 4226
rect 6578 4174 6580 4226
rect 6524 4162 6580 4174
rect 6636 7252 6692 7262
rect 6300 3666 6468 3668
rect 6300 3614 6302 3666
rect 6354 3614 6468 3666
rect 6300 3612 6468 3614
rect 6636 3666 6692 7196
rect 6860 6692 6916 6702
rect 6860 6598 6916 6636
rect 7420 6132 7476 7646
rect 8092 7252 8148 7262
rect 7756 7250 8148 7252
rect 7756 7198 8094 7250
rect 8146 7198 8148 7250
rect 7756 7196 8148 7198
rect 7420 6066 7476 6076
rect 7532 6692 7588 6702
rect 7196 5908 7252 5918
rect 7196 5814 7252 5852
rect 7532 5908 7588 6636
rect 7532 5814 7588 5852
rect 7196 5572 7252 5582
rect 6972 5516 7196 5572
rect 6972 5234 7028 5516
rect 7196 5506 7252 5516
rect 6972 5182 6974 5234
rect 7026 5182 7028 5234
rect 6972 5170 7028 5182
rect 6636 3614 6638 3666
rect 6690 3614 6692 3666
rect 6300 3602 6356 3612
rect 6636 3602 6692 3614
rect 6748 4900 6804 4910
rect 4508 3490 4564 3500
rect 6076 3556 6132 3566
rect 4172 3266 4228 3276
rect 3500 2034 3556 2044
rect 6076 800 6132 3500
rect 6748 800 6804 4844
rect 7196 4898 7252 4910
rect 7196 4846 7198 4898
rect 7250 4846 7252 4898
rect 7196 3388 7252 4846
rect 7532 4788 7588 4798
rect 7532 3442 7588 4732
rect 7756 4450 7812 7196
rect 8092 7186 8148 7196
rect 8092 6132 8148 6142
rect 8092 6038 8148 6076
rect 8092 5908 8148 5918
rect 8204 5908 8260 10668
rect 8316 10658 8372 10668
rect 8316 9828 8372 9838
rect 8316 9734 8372 9772
rect 8316 9604 8372 9614
rect 8316 9266 8372 9548
rect 8316 9214 8318 9266
rect 8370 9214 8372 9266
rect 8316 9202 8372 9214
rect 8428 7474 8484 10780
rect 8540 10610 8596 10622
rect 8540 10558 8542 10610
rect 8594 10558 8596 10610
rect 8540 9044 8596 10558
rect 8876 10052 8932 12348
rect 8988 12310 9044 12348
rect 9436 11396 9492 11406
rect 9436 11302 9492 11340
rect 9024 11004 9288 11014
rect 9080 10948 9128 11004
rect 9184 10948 9232 11004
rect 9024 10938 9288 10948
rect 9660 10836 9716 14476
rect 9772 13972 9828 14700
rect 9884 14530 9940 14812
rect 9884 14478 9886 14530
rect 9938 14478 9940 14530
rect 9884 14466 9940 14478
rect 9996 14532 10052 14542
rect 9884 13972 9940 13982
rect 9772 13970 9940 13972
rect 9772 13918 9886 13970
rect 9938 13918 9940 13970
rect 9772 13916 9940 13918
rect 9884 13906 9940 13916
rect 9996 13074 10052 14476
rect 10108 13636 10164 15092
rect 10108 13570 10164 13580
rect 9996 13022 9998 13074
rect 10050 13022 10052 13074
rect 9996 12404 10052 13022
rect 9996 12338 10052 12348
rect 9100 10834 9716 10836
rect 9100 10782 9662 10834
rect 9714 10782 9716 10834
rect 9100 10780 9716 10782
rect 9100 10610 9156 10780
rect 9100 10558 9102 10610
rect 9154 10558 9156 10610
rect 9100 10546 9156 10558
rect 9660 10386 9716 10780
rect 10108 10836 10164 10846
rect 10108 10742 10164 10780
rect 9660 10334 9662 10386
rect 9714 10334 9716 10386
rect 9660 10322 9716 10334
rect 8876 9996 9156 10052
rect 9100 9940 9156 9996
rect 9100 9938 9492 9940
rect 9100 9886 9102 9938
rect 9154 9886 9492 9938
rect 9100 9884 9492 9886
rect 9100 9874 9156 9884
rect 9024 9436 9288 9446
rect 9080 9380 9128 9436
rect 9184 9380 9232 9436
rect 9024 9370 9288 9380
rect 8540 8978 8596 8988
rect 9100 8818 9156 8830
rect 9100 8766 9102 8818
rect 9154 8766 9156 8818
rect 8764 8260 8820 8270
rect 8652 8036 8708 8046
rect 8652 7942 8708 7980
rect 8652 7700 8708 7710
rect 8764 7700 8820 8204
rect 9100 8148 9156 8766
rect 9436 8260 9492 9884
rect 9548 9156 9604 9166
rect 9548 9062 9604 9100
rect 9772 9042 9828 9054
rect 9772 8990 9774 9042
rect 9826 8990 9828 9042
rect 9436 8258 9716 8260
rect 9436 8206 9438 8258
rect 9490 8206 9716 8258
rect 9436 8204 9716 8206
rect 9436 8194 9492 8204
rect 9100 8082 9156 8092
rect 9212 8036 9268 8046
rect 9212 8034 9604 8036
rect 9212 7982 9214 8034
rect 9266 7982 9604 8034
rect 9212 7980 9604 7982
rect 9212 7970 9268 7980
rect 9024 7868 9288 7878
rect 9080 7812 9128 7868
rect 9184 7812 9232 7868
rect 9024 7802 9288 7812
rect 8652 7698 8820 7700
rect 8652 7646 8654 7698
rect 8706 7646 8820 7698
rect 8652 7644 8820 7646
rect 8652 7634 8708 7644
rect 8428 7422 8430 7474
rect 8482 7422 8484 7474
rect 8428 7410 8484 7422
rect 9436 6466 9492 6478
rect 9436 6414 9438 6466
rect 9490 6414 9492 6466
rect 9024 6300 9288 6310
rect 9080 6244 9128 6300
rect 9184 6244 9232 6300
rect 9024 6234 9288 6244
rect 8092 5906 8260 5908
rect 8092 5854 8094 5906
rect 8146 5854 8260 5906
rect 8092 5852 8260 5854
rect 8316 5908 8372 5918
rect 8372 5852 8484 5908
rect 8092 5572 8148 5852
rect 8316 5842 8372 5852
rect 8092 5506 8148 5516
rect 7980 4900 8036 4910
rect 8204 4900 8260 4910
rect 7980 4898 8148 4900
rect 7980 4846 7982 4898
rect 8034 4846 8148 4898
rect 7980 4844 8148 4846
rect 7980 4834 8036 4844
rect 7756 4398 7758 4450
rect 7810 4398 7812 4450
rect 7756 4386 7812 4398
rect 7532 3390 7534 3442
rect 7586 3390 7588 3442
rect 7196 3332 7476 3388
rect 7532 3378 7588 3390
rect 8092 3444 8148 4844
rect 8204 4806 8260 4844
rect 8428 4564 8484 5852
rect 9436 5348 9492 6414
rect 9548 6356 9604 7980
rect 9660 7700 9716 8204
rect 9772 7924 9828 8990
rect 9884 8258 9940 8270
rect 9884 8206 9886 8258
rect 9938 8206 9940 8258
rect 9884 7924 9940 8206
rect 9996 7924 10052 7934
rect 9884 7868 9996 7924
rect 9772 7858 9828 7868
rect 9996 7858 10052 7868
rect 10332 7812 10388 16828
rect 10780 13858 10836 17388
rect 11340 17378 11396 17388
rect 11004 17220 11060 17230
rect 10892 16996 10948 17006
rect 10892 15426 10948 16940
rect 11004 16996 11060 17164
rect 11004 16994 11172 16996
rect 11004 16942 11006 16994
rect 11058 16942 11172 16994
rect 11004 16940 11172 16942
rect 11004 16930 11060 16940
rect 10892 15374 10894 15426
rect 10946 15374 10948 15426
rect 10892 15362 10948 15374
rect 11116 15316 11172 16940
rect 11452 16882 11508 18396
rect 11564 17220 11620 19180
rect 11900 19124 11956 19294
rect 12348 19348 12404 21756
rect 12460 21746 12516 21756
rect 12572 21364 12628 21374
rect 12572 20802 12628 21308
rect 12930 21196 13194 21206
rect 12986 21140 13034 21196
rect 13090 21140 13138 21196
rect 12930 21130 13194 21140
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12572 20738 12628 20750
rect 12796 20692 12852 20702
rect 13356 20692 13412 23326
rect 13580 22372 13636 22382
rect 13580 22278 13636 22316
rect 13468 20692 13524 20702
rect 13356 20690 13524 20692
rect 13356 20638 13470 20690
rect 13522 20638 13524 20690
rect 13356 20636 13524 20638
rect 12796 20598 12852 20636
rect 13468 20626 13524 20636
rect 13692 20580 13748 26124
rect 14028 25732 14084 26236
rect 15148 26852 15428 26908
rect 14028 25666 14084 25676
rect 14588 25732 14644 25742
rect 14588 25638 14644 25676
rect 13804 25508 13860 25518
rect 13804 25414 13860 25452
rect 13916 25284 13972 25294
rect 15148 25284 15204 26852
rect 13972 25228 14084 25284
rect 13916 25218 13972 25228
rect 13916 23940 13972 23950
rect 13916 23846 13972 23884
rect 13916 22932 13972 22942
rect 13804 22930 13972 22932
rect 13804 22878 13918 22930
rect 13970 22878 13972 22930
rect 13804 22876 13972 22878
rect 13804 21028 13860 22876
rect 13916 22866 13972 22876
rect 14028 22482 14084 25228
rect 14924 25228 15204 25284
rect 15260 25508 15316 25518
rect 14700 24946 14756 24958
rect 14700 24894 14702 24946
rect 14754 24894 14756 24946
rect 14700 24612 14756 24894
rect 14812 24836 14868 24846
rect 14924 24836 14980 25228
rect 15260 25060 15316 25452
rect 14868 24780 14980 24836
rect 15148 25004 15316 25060
rect 14812 24770 14868 24780
rect 14700 24546 14756 24556
rect 14140 23492 14196 23502
rect 14140 23154 14196 23436
rect 14140 23102 14142 23154
rect 14194 23102 14196 23154
rect 14140 23090 14196 23102
rect 15148 23378 15204 25004
rect 15484 24948 15540 24958
rect 15484 24854 15540 24892
rect 15260 24836 15316 24846
rect 15260 24742 15316 24780
rect 15932 24610 15988 28140
rect 16380 28082 16436 28094
rect 16380 28030 16382 28082
rect 16434 28030 16436 28082
rect 16268 27074 16324 27086
rect 16268 27022 16270 27074
rect 16322 27022 16324 27074
rect 16268 26964 16324 27022
rect 16268 26898 16324 26908
rect 16380 26852 16436 28030
rect 16604 27074 16660 28588
rect 16604 27022 16606 27074
rect 16658 27022 16660 27074
rect 16604 27010 16660 27022
rect 16716 26908 16772 29484
rect 17052 28866 17108 29484
rect 17500 29426 17556 29438
rect 17500 29374 17502 29426
rect 17554 29374 17556 29426
rect 17052 28814 17054 28866
rect 17106 28814 17108 28866
rect 17052 28802 17108 28814
rect 17164 28868 17220 28878
rect 16836 28252 17100 28262
rect 16892 28196 16940 28252
rect 16996 28196 17044 28252
rect 16836 28186 17100 28196
rect 16940 28084 16996 28094
rect 17164 28084 17220 28812
rect 16940 28082 17220 28084
rect 16940 28030 16942 28082
rect 16994 28030 17220 28082
rect 16940 28028 17220 28030
rect 17276 28642 17332 28654
rect 17276 28590 17278 28642
rect 17330 28590 17332 28642
rect 16940 28018 16996 28028
rect 16380 26786 16436 26796
rect 16604 26852 16772 26908
rect 17164 27860 17220 27870
rect 16380 26514 16436 26526
rect 16380 26462 16382 26514
rect 16434 26462 16436 26514
rect 16380 26404 16436 26462
rect 16380 26338 16436 26348
rect 15932 24558 15934 24610
rect 15986 24558 15988 24610
rect 15932 24546 15988 24558
rect 16492 25618 16548 25630
rect 16492 25566 16494 25618
rect 16546 25566 16548 25618
rect 15148 23326 15150 23378
rect 15202 23326 15204 23378
rect 14028 22430 14030 22482
rect 14082 22430 14084 22482
rect 14028 22418 14084 22430
rect 13804 20962 13860 20972
rect 13916 22372 13972 22382
rect 13916 20916 13972 22316
rect 15036 22372 15092 22382
rect 15036 22278 15092 22316
rect 14700 22146 14756 22158
rect 14700 22094 14702 22146
rect 14754 22094 14756 22146
rect 14252 20916 14308 20926
rect 13916 20914 14308 20916
rect 13916 20862 14254 20914
rect 14306 20862 14308 20914
rect 13916 20860 14308 20862
rect 13804 20804 13860 20814
rect 13916 20804 13972 20860
rect 14252 20850 14308 20860
rect 13860 20748 13972 20804
rect 13804 20710 13860 20748
rect 13580 20524 13748 20580
rect 12796 20020 12852 20030
rect 12572 20018 12852 20020
rect 12572 19966 12798 20018
rect 12850 19966 12852 20018
rect 12572 19964 12852 19966
rect 12460 19348 12516 19358
rect 12348 19346 12516 19348
rect 12348 19294 12462 19346
rect 12514 19294 12516 19346
rect 12348 19292 12516 19294
rect 12460 19282 12516 19292
rect 12572 19124 12628 19964
rect 12796 19954 12852 19964
rect 12930 19628 13194 19638
rect 12986 19572 13034 19628
rect 13090 19572 13138 19628
rect 12930 19562 13194 19572
rect 13020 19458 13076 19470
rect 13020 19406 13022 19458
rect 13074 19406 13076 19458
rect 12908 19348 12964 19358
rect 12908 19254 12964 19292
rect 11900 19068 12628 19124
rect 12460 18452 12516 18462
rect 11900 18450 12516 18452
rect 11900 18398 12462 18450
rect 12514 18398 12516 18450
rect 11900 18396 12516 18398
rect 11676 18340 11732 18350
rect 11676 17778 11732 18284
rect 11676 17726 11678 17778
rect 11730 17726 11732 17778
rect 11676 17714 11732 17726
rect 11788 18228 11844 18238
rect 11564 17154 11620 17164
rect 11452 16830 11454 16882
rect 11506 16830 11508 16882
rect 11452 16818 11508 16830
rect 11788 16882 11844 18172
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 11788 16818 11844 16830
rect 11900 16324 11956 18396
rect 12460 18386 12516 18396
rect 13020 18452 13076 19406
rect 13468 19124 13524 19134
rect 13580 19124 13636 20524
rect 14476 19796 14532 19806
rect 14476 19458 14532 19740
rect 14476 19406 14478 19458
rect 14530 19406 14532 19458
rect 14476 19394 14532 19406
rect 13692 19348 13748 19358
rect 13692 19234 13748 19292
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13692 19170 13748 19182
rect 13468 19122 13636 19124
rect 13468 19070 13470 19122
rect 13522 19070 13636 19122
rect 13468 19068 13636 19070
rect 13468 19058 13524 19068
rect 13244 18452 13300 18462
rect 13076 18450 13300 18452
rect 13076 18398 13246 18450
rect 13298 18398 13300 18450
rect 13076 18396 13300 18398
rect 13020 18358 13076 18396
rect 13244 18386 13300 18396
rect 13916 18452 13972 18462
rect 13916 18358 13972 18396
rect 14364 18228 14420 18238
rect 11788 16268 11956 16324
rect 12012 18116 12068 18126
rect 11228 16100 11284 16110
rect 11228 16006 11284 16044
rect 11788 15316 11844 16268
rect 11900 16098 11956 16110
rect 11900 16046 11902 16098
rect 11954 16046 11956 16098
rect 11900 15540 11956 16046
rect 12012 15988 12068 18060
rect 12930 18060 13194 18070
rect 12986 18004 13034 18060
rect 13090 18004 13138 18060
rect 12930 17994 13194 18004
rect 12124 17780 12180 17790
rect 12124 17686 12180 17724
rect 12348 17666 12404 17678
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12348 17220 12404 17614
rect 14364 17554 14420 18172
rect 14364 17502 14366 17554
rect 14418 17502 14420 17554
rect 14364 17490 14420 17502
rect 12348 17154 12404 17164
rect 12908 17442 12964 17454
rect 12908 17390 12910 17442
rect 12962 17390 12964 17442
rect 12908 17220 12964 17390
rect 12908 17154 12964 17164
rect 13580 17442 13636 17454
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13580 17220 13636 17390
rect 13636 17164 13972 17220
rect 13580 17154 13636 17164
rect 12572 16884 12628 16894
rect 12124 15988 12180 15998
rect 12012 15986 12180 15988
rect 12012 15934 12126 15986
rect 12178 15934 12180 15986
rect 12012 15932 12180 15934
rect 12124 15922 12180 15932
rect 12460 15986 12516 15998
rect 12460 15934 12462 15986
rect 12514 15934 12516 15986
rect 11900 15484 12180 15540
rect 11116 15250 11172 15260
rect 11676 15260 11844 15316
rect 11676 14868 11732 15260
rect 12124 15148 12180 15484
rect 11788 15092 11844 15102
rect 12124 15092 12404 15148
rect 11788 15090 12068 15092
rect 11788 15038 11790 15090
rect 11842 15038 12068 15090
rect 11788 15036 12068 15038
rect 11788 15026 11844 15036
rect 11676 14812 11844 14868
rect 10780 13806 10782 13858
rect 10834 13806 10836 13858
rect 10780 13794 10836 13806
rect 10892 14308 10948 14318
rect 10892 12850 10948 14252
rect 10892 12798 10894 12850
rect 10946 12798 10948 12850
rect 10892 12786 10948 12798
rect 11676 13636 11732 13646
rect 11676 12180 11732 13580
rect 11788 13634 11844 14812
rect 11788 13582 11790 13634
rect 11842 13582 11844 13634
rect 11788 13570 11844 13582
rect 11900 13748 11956 13758
rect 11900 13074 11956 13692
rect 11900 13022 11902 13074
rect 11954 13022 11956 13074
rect 11900 13010 11956 13022
rect 12012 12852 12068 15036
rect 12348 14532 12404 15092
rect 12460 14644 12516 15934
rect 12572 15538 12628 16828
rect 12930 16492 13194 16502
rect 12986 16436 13034 16492
rect 13090 16436 13138 16492
rect 12930 16426 13194 16436
rect 13916 16322 13972 17164
rect 14364 17108 14420 17118
rect 14364 17014 14420 17052
rect 13916 16270 13918 16322
rect 13970 16270 13972 16322
rect 13916 16258 13972 16270
rect 13020 16212 13076 16222
rect 13020 16118 13076 16156
rect 12572 15486 12574 15538
rect 12626 15486 12628 15538
rect 12572 15474 12628 15486
rect 14700 14980 14756 22094
rect 14924 20804 14980 20814
rect 14812 20748 14924 20804
rect 14812 16212 14868 20748
rect 14924 20738 14980 20748
rect 15148 20804 15204 23326
rect 15148 20710 15204 20748
rect 15260 24052 15316 24062
rect 15260 20580 15316 23996
rect 16380 23714 16436 23726
rect 16380 23662 16382 23714
rect 16434 23662 16436 23714
rect 16380 23268 16436 23662
rect 16380 23202 16436 23212
rect 16156 22370 16212 22382
rect 16156 22318 16158 22370
rect 16210 22318 16212 22370
rect 15148 20524 15316 20580
rect 15372 22258 15428 22270
rect 15372 22206 15374 22258
rect 15426 22206 15428 22258
rect 14924 16660 14980 16670
rect 14924 16566 14980 16604
rect 14812 16098 14868 16156
rect 14812 16046 14814 16098
rect 14866 16046 14868 16098
rect 14812 16034 14868 16046
rect 15148 15540 15204 20524
rect 15372 20242 15428 22206
rect 16156 22148 16212 22318
rect 16492 22370 16548 25566
rect 16604 24948 16660 26852
rect 16836 26684 17100 26694
rect 16892 26628 16940 26684
rect 16996 26628 17044 26684
rect 16836 26618 17100 26628
rect 16940 26516 16996 26526
rect 17164 26516 17220 27804
rect 17276 26964 17332 28590
rect 17276 26898 17332 26908
rect 17500 26908 17556 29374
rect 17724 29316 17780 29326
rect 17724 28642 17780 29260
rect 17836 29314 17892 29596
rect 17836 29262 17838 29314
rect 17890 29262 17892 29314
rect 17836 29250 17892 29262
rect 17724 28590 17726 28642
rect 17778 28590 17780 28642
rect 17724 28578 17780 28590
rect 17948 28644 18004 30270
rect 18172 30212 18228 33200
rect 18172 30146 18228 30156
rect 18844 29652 18900 33200
rect 20742 30604 21006 30614
rect 20798 30548 20846 30604
rect 20902 30548 20950 30604
rect 20742 30538 21006 30548
rect 21756 30322 21812 30334
rect 21756 30270 21758 30322
rect 21810 30270 21812 30322
rect 19964 30212 20020 30222
rect 19964 30118 20020 30156
rect 21420 30212 21476 30222
rect 21420 30118 21476 30156
rect 19180 30098 19236 30110
rect 19180 30046 19182 30098
rect 19234 30046 19236 30098
rect 19068 29652 19124 29662
rect 18844 29650 19124 29652
rect 18844 29598 19070 29650
rect 19122 29598 19124 29650
rect 18844 29596 19124 29598
rect 19068 29586 19124 29596
rect 17948 28578 18004 28588
rect 18844 28308 18900 28318
rect 18732 27748 18788 27758
rect 18732 27654 18788 27692
rect 17500 26852 18004 26908
rect 16940 26514 17220 26516
rect 16940 26462 16942 26514
rect 16994 26462 17220 26514
rect 16940 26460 17220 26462
rect 16940 26450 16996 26460
rect 17388 26404 17444 26414
rect 17388 26310 17444 26348
rect 17724 26178 17780 26190
rect 17724 26126 17726 26178
rect 17778 26126 17780 26178
rect 16828 25732 16884 25742
rect 16828 25284 16884 25676
rect 17612 25732 17668 25742
rect 17500 25396 17556 25406
rect 16716 25228 16884 25284
rect 17164 25394 17556 25396
rect 17164 25342 17502 25394
rect 17554 25342 17556 25394
rect 17164 25340 17556 25342
rect 16716 24948 16772 25228
rect 16836 25116 17100 25126
rect 16892 25060 16940 25116
rect 16996 25060 17044 25116
rect 16836 25050 17100 25060
rect 16828 24948 16884 24958
rect 16716 24946 16884 24948
rect 16716 24894 16830 24946
rect 16882 24894 16884 24946
rect 16716 24892 16884 24894
rect 16604 24882 16660 24892
rect 16828 24882 16884 24892
rect 17052 24164 17108 24174
rect 17164 24164 17220 25340
rect 17500 25330 17556 25340
rect 17612 24836 17668 25676
rect 17500 24780 17668 24836
rect 17500 24722 17556 24780
rect 17500 24670 17502 24722
rect 17554 24670 17556 24722
rect 17500 24658 17556 24670
rect 17724 24724 17780 26126
rect 17724 24658 17780 24668
rect 17836 25620 17892 25630
rect 17612 24612 17668 24622
rect 17612 24518 17668 24556
rect 17052 24162 17220 24164
rect 17052 24110 17054 24162
rect 17106 24110 17220 24162
rect 17052 24108 17220 24110
rect 17052 24098 17108 24108
rect 17164 23938 17220 23950
rect 17164 23886 17166 23938
rect 17218 23886 17220 23938
rect 16836 23548 17100 23558
rect 16892 23492 16940 23548
rect 16996 23492 17044 23548
rect 16836 23482 17100 23492
rect 16492 22318 16494 22370
rect 16546 22318 16548 22370
rect 16492 22306 16548 22318
rect 16716 23156 16772 23166
rect 16156 22082 16212 22092
rect 16268 21812 16324 21822
rect 16716 21812 16772 23100
rect 17164 22148 17220 23886
rect 17836 23938 17892 25564
rect 17836 23886 17838 23938
rect 17890 23886 17892 23938
rect 17836 23874 17892 23886
rect 17724 23380 17780 23390
rect 17724 23286 17780 23324
rect 17500 23156 17556 23166
rect 17500 23154 17780 23156
rect 17500 23102 17502 23154
rect 17554 23102 17780 23154
rect 17500 23100 17780 23102
rect 17500 23090 17556 23100
rect 17164 22082 17220 22092
rect 16836 21980 17100 21990
rect 16892 21924 16940 21980
rect 16996 21924 17044 21980
rect 16836 21914 17100 21924
rect 16324 21810 16772 21812
rect 16324 21758 16718 21810
rect 16770 21758 16772 21810
rect 16324 21756 16772 21758
rect 16268 21586 16324 21756
rect 16716 21746 16772 21756
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21522 16324 21534
rect 17500 20916 17556 20926
rect 17500 20578 17556 20860
rect 17500 20526 17502 20578
rect 17554 20526 17556 20578
rect 16836 20412 17100 20422
rect 16892 20356 16940 20412
rect 16996 20356 17044 20412
rect 16836 20346 17100 20356
rect 15372 20190 15374 20242
rect 15426 20190 15428 20242
rect 15372 20178 15428 20190
rect 15932 20132 15988 20142
rect 15932 20038 15988 20076
rect 16492 19908 16548 19918
rect 16044 19906 16548 19908
rect 16044 19854 16494 19906
rect 16546 19854 16548 19906
rect 16044 19852 16548 19854
rect 16044 19460 16100 19852
rect 16492 19842 16548 19852
rect 16828 19908 16884 19918
rect 17500 19908 17556 20526
rect 16828 19906 17556 19908
rect 16828 19854 16830 19906
rect 16882 19854 17502 19906
rect 17554 19854 17556 19906
rect 16828 19852 17556 19854
rect 16828 19842 16884 19852
rect 15260 19404 16100 19460
rect 16716 19460 16772 19470
rect 15260 19122 15316 19404
rect 15260 19070 15262 19122
rect 15314 19070 15316 19122
rect 15260 19058 15316 19070
rect 16380 18674 16436 18686
rect 16380 18622 16382 18674
rect 16434 18622 16436 18674
rect 15372 17778 15428 17790
rect 15372 17726 15374 17778
rect 15426 17726 15428 17778
rect 15372 17668 15428 17726
rect 15372 17602 15428 17612
rect 15820 17442 15876 17454
rect 15820 17390 15822 17442
rect 15874 17390 15876 17442
rect 15484 17220 15540 17230
rect 15820 17220 15876 17390
rect 16268 17442 16324 17454
rect 16268 17390 16270 17442
rect 16322 17390 16324 17442
rect 16268 17220 16324 17390
rect 15540 17164 16324 17220
rect 15260 16996 15316 17006
rect 15260 16902 15316 16940
rect 15484 16882 15540 17164
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16818 15540 16830
rect 15932 16884 15988 16894
rect 15932 16790 15988 16828
rect 16156 16882 16212 17164
rect 16380 17108 16436 18622
rect 16604 18564 16660 18574
rect 16604 17666 16660 18508
rect 16604 17614 16606 17666
rect 16658 17614 16660 17666
rect 16604 17602 16660 17614
rect 16716 17108 16772 19404
rect 16836 18844 17100 18854
rect 16892 18788 16940 18844
rect 16996 18788 17044 18844
rect 16836 18778 17100 18788
rect 17388 18562 17444 18574
rect 17388 18510 17390 18562
rect 17442 18510 17444 18562
rect 16940 18228 16996 18238
rect 16940 18134 16996 18172
rect 17164 17668 17220 17678
rect 17164 17574 17220 17612
rect 16836 17276 17100 17286
rect 16892 17220 16940 17276
rect 16996 17220 17044 17276
rect 16836 17210 17100 17220
rect 16828 17108 16884 17118
rect 16716 17106 16884 17108
rect 16716 17054 16830 17106
rect 16882 17054 16884 17106
rect 16716 17052 16884 17054
rect 16380 17042 16436 17052
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 16156 16818 16212 16830
rect 16828 16884 16884 17052
rect 16828 16818 16884 16828
rect 15820 16660 15876 16670
rect 15148 15474 15204 15484
rect 15484 16098 15540 16110
rect 15484 16046 15486 16098
rect 15538 16046 15540 16098
rect 12930 14924 13194 14934
rect 12986 14868 13034 14924
rect 13090 14868 13138 14924
rect 14700 14914 14756 14924
rect 14812 15314 14868 15326
rect 14812 15262 14814 15314
rect 14866 15262 14868 15314
rect 12930 14858 13194 14868
rect 12460 14578 12516 14588
rect 14812 14642 14868 15262
rect 15484 15314 15540 16046
rect 15484 15262 15486 15314
rect 15538 15262 15540 15314
rect 15484 15148 15540 15262
rect 14812 14590 14814 14642
rect 14866 14590 14868 14642
rect 14812 14578 14868 14590
rect 15260 15092 15540 15148
rect 12348 13970 12404 14476
rect 12348 13918 12350 13970
rect 12402 13918 12404 13970
rect 12348 13906 12404 13918
rect 12460 14306 12516 14318
rect 12460 14254 12462 14306
rect 12514 14254 12516 14306
rect 12460 13076 12516 14254
rect 13020 14308 13076 14318
rect 13580 14308 13636 14318
rect 14028 14308 14084 14318
rect 14476 14308 14532 14318
rect 13020 14214 13076 14252
rect 13356 14306 14532 14308
rect 13356 14254 13582 14306
rect 13634 14254 14030 14306
rect 14082 14254 14478 14306
rect 14530 14254 14532 14306
rect 13356 14252 14532 14254
rect 13356 13746 13412 14252
rect 13580 14242 13636 14252
rect 14028 14242 14084 14252
rect 13356 13694 13358 13746
rect 13410 13694 13412 13746
rect 13356 13682 13412 13694
rect 13692 13748 13748 13758
rect 13692 13654 13748 13692
rect 14476 13748 14532 14252
rect 14476 13682 14532 13692
rect 15260 13748 15316 15092
rect 15820 14418 15876 16604
rect 16156 16100 16212 16110
rect 16156 16098 16772 16100
rect 16156 16046 16158 16098
rect 16210 16046 16772 16098
rect 16156 16044 16772 16046
rect 16156 16034 16212 16044
rect 16492 15314 16548 15326
rect 16492 15262 16494 15314
rect 16546 15262 16548 15314
rect 15820 14366 15822 14418
rect 15874 14366 15876 14418
rect 15820 14354 15876 14366
rect 16044 15202 16100 15214
rect 16044 15150 16046 15202
rect 16098 15150 16100 15202
rect 16044 13970 16100 15150
rect 16044 13918 16046 13970
rect 16098 13918 16100 13970
rect 16044 13906 16100 13918
rect 16380 14644 16436 14654
rect 15260 13682 15316 13692
rect 16156 13748 16212 13758
rect 12796 13636 12852 13646
rect 12796 13542 12852 13580
rect 12930 13356 13194 13366
rect 12986 13300 13034 13356
rect 13090 13300 13138 13356
rect 12930 13290 13194 13300
rect 13692 13300 13748 13310
rect 12460 13010 12516 13020
rect 13580 13076 13636 13086
rect 13580 12982 13636 13020
rect 12012 12786 12068 12796
rect 13692 12962 13748 13244
rect 15372 13300 15428 13310
rect 15372 13074 15428 13244
rect 15372 13022 15374 13074
rect 15426 13022 15428 13074
rect 15372 13010 15428 13022
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 12460 12738 12516 12750
rect 12460 12686 12462 12738
rect 12514 12686 12516 12738
rect 12460 12180 12516 12686
rect 12908 12740 12964 12750
rect 12908 12646 12964 12684
rect 13692 12740 13748 12910
rect 14588 12964 14644 12974
rect 14812 12964 14868 12974
rect 14588 12850 14644 12908
rect 14588 12798 14590 12850
rect 14642 12798 14644 12850
rect 14588 12786 14644 12798
rect 14700 12962 14868 12964
rect 14700 12910 14814 12962
rect 14866 12910 14868 12962
rect 14700 12908 14868 12910
rect 12796 12180 12852 12190
rect 12460 12178 12852 12180
rect 12460 12126 12798 12178
rect 12850 12126 12852 12178
rect 12460 12124 12852 12126
rect 10444 12066 10500 12078
rect 10444 12014 10446 12066
rect 10498 12014 10500 12066
rect 10444 9268 10500 12014
rect 11676 11506 11732 12124
rect 11676 11454 11678 11506
rect 11730 11454 11732 11506
rect 10892 11396 10948 11406
rect 10556 10836 10612 10846
rect 10556 10742 10612 10780
rect 10892 10610 10948 11340
rect 11676 10836 11732 11454
rect 12796 11396 12852 12124
rect 12930 11788 13194 11798
rect 12986 11732 13034 11788
rect 13090 11732 13138 11788
rect 12930 11722 13194 11732
rect 12908 11396 12964 11406
rect 12796 11340 12908 11396
rect 12908 11302 12964 11340
rect 13468 11394 13524 11406
rect 13468 11342 13470 11394
rect 13522 11342 13524 11394
rect 11676 10770 11732 10780
rect 13468 11172 13524 11342
rect 10892 10558 10894 10610
rect 10946 10558 10948 10610
rect 10892 10546 10948 10558
rect 10444 9174 10500 9212
rect 10668 10386 10724 10398
rect 10668 10334 10670 10386
rect 10722 10334 10724 10386
rect 10668 8932 10724 10334
rect 10892 10388 10948 10398
rect 10892 9828 10948 10332
rect 13468 10388 13524 11116
rect 13468 10322 13524 10332
rect 13692 10386 13748 12684
rect 14364 12180 14420 12190
rect 14364 12086 14420 12124
rect 13692 10334 13694 10386
rect 13746 10334 13748 10386
rect 12930 10220 13194 10230
rect 12986 10164 13034 10220
rect 13090 10164 13138 10220
rect 12930 10154 13194 10164
rect 10332 7756 10500 7812
rect 9660 7698 10388 7700
rect 9660 7646 9662 7698
rect 9714 7646 10388 7698
rect 9660 7644 10388 7646
rect 9660 7634 9716 7644
rect 10108 7362 10164 7374
rect 10108 7310 10110 7362
rect 10162 7310 10164 7362
rect 9772 6468 9828 6478
rect 9548 6300 9716 6356
rect 9548 6132 9604 6142
rect 9548 6038 9604 6076
rect 9436 5282 9492 5292
rect 8764 5012 8820 5022
rect 8764 4898 8820 4956
rect 8764 4846 8766 4898
rect 8818 4846 8820 4898
rect 8764 4834 8820 4846
rect 9024 4732 9288 4742
rect 9080 4676 9128 4732
rect 9184 4676 9232 4732
rect 9024 4666 9288 4676
rect 8988 4564 9044 4574
rect 8428 4562 9044 4564
rect 8428 4510 8430 4562
rect 8482 4510 8990 4562
rect 9042 4510 9044 4562
rect 8428 4508 9044 4510
rect 8428 4498 8484 4508
rect 8988 4498 9044 4508
rect 9660 4564 9716 6300
rect 9772 5906 9828 6412
rect 9772 5854 9774 5906
rect 9826 5854 9828 5906
rect 9772 5842 9828 5854
rect 9996 6466 10052 6478
rect 9996 6414 9998 6466
rect 10050 6414 10052 6466
rect 9660 4498 9716 4508
rect 8316 3444 8372 3454
rect 8092 3442 8372 3444
rect 8092 3390 8318 3442
rect 8370 3390 8372 3442
rect 8092 3388 8372 3390
rect 8316 3378 8372 3388
rect 8652 3444 8708 3482
rect 8652 3378 8708 3388
rect 9996 3442 10052 6414
rect 10108 5124 10164 7310
rect 10332 6692 10388 7644
rect 10332 6598 10388 6636
rect 10444 6132 10500 7756
rect 10444 6066 10500 6076
rect 10668 7476 10724 8876
rect 10780 9380 10836 9390
rect 10780 7698 10836 9324
rect 10892 9266 10948 9772
rect 11340 9828 11396 9838
rect 10892 9214 10894 9266
rect 10946 9214 10948 9266
rect 10892 9202 10948 9214
rect 11228 9268 11284 9278
rect 11228 9174 11284 9212
rect 10780 7646 10782 7698
rect 10834 7646 10836 7698
rect 10780 7634 10836 7646
rect 11228 7924 11284 7934
rect 11116 7476 11172 7486
rect 10668 7474 11172 7476
rect 10668 7422 11118 7474
rect 11170 7422 11172 7474
rect 10668 7420 11172 7422
rect 10668 6580 10724 7420
rect 11116 7410 11172 7420
rect 11228 6802 11284 7868
rect 11340 6916 11396 9772
rect 13468 9826 13524 9838
rect 13468 9774 13470 9826
rect 13522 9774 13524 9826
rect 12460 9604 12516 9614
rect 11676 8930 11732 8942
rect 11676 8878 11678 8930
rect 11730 8878 11732 8930
rect 11676 7474 11732 8878
rect 11676 7422 11678 7474
rect 11730 7422 11732 7474
rect 11676 7410 11732 7422
rect 12236 8148 12292 8158
rect 11340 6850 11396 6860
rect 11228 6750 11230 6802
rect 11282 6750 11284 6802
rect 11228 6738 11284 6750
rect 10780 6692 10836 6702
rect 10780 6598 10836 6636
rect 11676 6692 11732 6702
rect 10668 5906 10724 6524
rect 10668 5854 10670 5906
rect 10722 5854 10724 5906
rect 10668 5842 10724 5854
rect 11116 5906 11172 5918
rect 11116 5854 11118 5906
rect 11170 5854 11172 5906
rect 10108 5058 10164 5068
rect 10108 4900 10164 4910
rect 10108 4450 10164 4844
rect 10108 4398 10110 4450
rect 10162 4398 10164 4450
rect 10108 4386 10164 4398
rect 11116 4226 11172 5854
rect 11116 4174 11118 4226
rect 11170 4174 11172 4226
rect 11116 4162 11172 4174
rect 11228 5122 11284 5134
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 11004 3668 11060 3678
rect 11228 3668 11284 5070
rect 11676 5124 11732 6636
rect 12236 6578 12292 8092
rect 12460 8034 12516 9548
rect 12460 7982 12462 8034
rect 12514 7982 12516 8034
rect 12460 7970 12516 7982
rect 12684 9602 12740 9614
rect 12684 9550 12686 9602
rect 12738 9550 12740 9602
rect 12236 6526 12238 6578
rect 12290 6526 12292 6578
rect 12236 6514 12292 6526
rect 12684 5684 12740 9550
rect 13468 9268 13524 9774
rect 13580 9604 13636 9614
rect 13580 9510 13636 9548
rect 13468 9202 13524 9212
rect 12796 9154 12852 9166
rect 12796 9102 12798 9154
rect 12850 9102 12852 9154
rect 12796 8484 12852 9102
rect 13244 9042 13300 9054
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 13244 8932 13300 8990
rect 13244 8866 13300 8876
rect 12930 8652 13194 8662
rect 12986 8596 13034 8652
rect 13090 8596 13138 8652
rect 12930 8586 13194 8596
rect 13020 8484 13076 8494
rect 12796 8482 13076 8484
rect 12796 8430 13022 8482
rect 13074 8430 13076 8482
rect 12796 8428 13076 8430
rect 13020 8418 13076 8428
rect 12930 7084 13194 7094
rect 12986 7028 13034 7084
rect 13090 7028 13138 7084
rect 12930 7018 13194 7028
rect 13468 6578 13524 6590
rect 13468 6526 13470 6578
rect 13522 6526 13524 6578
rect 13356 6020 13412 6030
rect 12236 5628 12740 5684
rect 12796 6018 13412 6020
rect 12796 5966 13358 6018
rect 13410 5966 13412 6018
rect 12796 5964 13412 5966
rect 11676 5122 11956 5124
rect 11676 5070 11678 5122
rect 11730 5070 11956 5122
rect 11676 5068 11956 5070
rect 11676 5058 11732 5068
rect 11900 4562 11956 5068
rect 11900 4510 11902 4562
rect 11954 4510 11956 4562
rect 11900 4498 11956 4510
rect 11004 3666 11284 3668
rect 11004 3614 11006 3666
rect 11058 3614 11284 3666
rect 11004 3612 11284 3614
rect 11004 3602 11060 3612
rect 12124 3556 12180 3566
rect 12124 3462 12180 3500
rect 9996 3390 9998 3442
rect 10050 3390 10052 3442
rect 9996 3378 10052 3390
rect 7420 800 7476 3332
rect 9024 3164 9288 3174
rect 9080 3108 9128 3164
rect 9184 3108 9232 3164
rect 9024 3098 9288 3108
rect 12236 2772 12292 5628
rect 12572 5460 12628 5470
rect 12572 5124 12628 5404
rect 12796 5346 12852 5964
rect 13356 5954 13412 5964
rect 13468 6020 13524 6526
rect 13468 5954 13524 5964
rect 13692 5908 13748 10334
rect 14028 12066 14084 12078
rect 14028 12014 14030 12066
rect 14082 12014 14084 12066
rect 14028 9716 14084 12014
rect 14700 11508 14756 12908
rect 14812 12898 14868 12908
rect 16156 12738 16212 13692
rect 16156 12686 16158 12738
rect 16210 12686 16212 12738
rect 15148 12180 15204 12190
rect 14924 12068 14980 12078
rect 14924 11974 14980 12012
rect 14700 11442 14756 11452
rect 15148 10610 15204 12124
rect 15260 11956 15316 11966
rect 15260 11862 15316 11900
rect 15148 10558 15150 10610
rect 15202 10558 15204 10610
rect 15148 10546 15204 10558
rect 15372 11732 15428 11742
rect 15260 10500 15316 10510
rect 15260 10406 15316 10444
rect 14028 9650 14084 9660
rect 14812 9826 14868 9838
rect 14812 9774 14814 9826
rect 14866 9774 14868 9826
rect 14812 9716 14868 9774
rect 14812 9650 14868 9660
rect 15260 9826 15316 9838
rect 15260 9774 15262 9826
rect 15314 9774 15316 9826
rect 14588 9602 14644 9614
rect 14588 9550 14590 9602
rect 14642 9550 14644 9602
rect 14252 9268 14308 9278
rect 13916 9044 13972 9054
rect 13916 9042 14084 9044
rect 13916 8990 13918 9042
rect 13970 8990 14084 9042
rect 13916 8988 14084 8990
rect 13916 8978 13972 8988
rect 13804 8932 13860 8942
rect 13804 6578 13860 8876
rect 14028 7140 14084 8988
rect 14252 8372 14308 9212
rect 14252 8258 14308 8316
rect 14252 8206 14254 8258
rect 14306 8206 14308 8258
rect 14140 8034 14196 8046
rect 14140 7982 14142 8034
rect 14194 7982 14196 8034
rect 14140 7698 14196 7982
rect 14140 7646 14142 7698
rect 14194 7646 14196 7698
rect 14140 7634 14196 7646
rect 14028 7074 14084 7084
rect 14252 6802 14308 8206
rect 14252 6750 14254 6802
rect 14306 6750 14308 6802
rect 14252 6738 14308 6750
rect 13804 6526 13806 6578
rect 13858 6526 13860 6578
rect 13804 6514 13860 6526
rect 14476 6020 14532 6030
rect 14476 5926 14532 5964
rect 13916 5908 13972 5918
rect 13692 5852 13916 5908
rect 12930 5516 13194 5526
rect 12986 5460 13034 5516
rect 13090 5460 13138 5516
rect 12930 5450 13194 5460
rect 12796 5294 12798 5346
rect 12850 5294 12852 5346
rect 12796 5282 12852 5294
rect 12348 5068 12572 5124
rect 12348 4562 12404 5068
rect 12572 5030 12628 5068
rect 13916 5124 13972 5852
rect 14140 5684 14196 5694
rect 14140 5682 14308 5684
rect 14140 5630 14142 5682
rect 14194 5630 14308 5682
rect 14140 5628 14308 5630
rect 14140 5618 14196 5628
rect 12348 4510 12350 4562
rect 12402 4510 12404 4562
rect 12348 4498 12404 4510
rect 12796 4340 12852 4350
rect 12796 4246 12852 4284
rect 13244 4338 13300 4350
rect 13244 4286 13246 4338
rect 13298 4286 13300 4338
rect 13244 4116 13300 4286
rect 13244 4050 13300 4060
rect 12930 3948 13194 3958
rect 12986 3892 13034 3948
rect 13090 3892 13138 3948
rect 12930 3882 13194 3892
rect 13916 3668 13972 5068
rect 14140 4900 14196 4910
rect 14140 4806 14196 4844
rect 14028 3668 14084 3678
rect 13916 3666 14084 3668
rect 13916 3614 14030 3666
rect 14082 3614 14084 3666
rect 13916 3612 14084 3614
rect 14028 3602 14084 3612
rect 13356 3556 13412 3566
rect 13132 3444 13188 3482
rect 13356 3462 13412 3500
rect 13132 3378 13188 3388
rect 14252 3444 14308 5628
rect 14588 4676 14644 9550
rect 14812 9156 14868 9166
rect 14812 8370 14868 9100
rect 15260 8484 15316 9774
rect 15260 8418 15316 8428
rect 14812 8318 14814 8370
rect 14866 8318 14868 8370
rect 14812 8306 14868 8318
rect 15036 8372 15092 8382
rect 15036 8258 15092 8316
rect 15036 8206 15038 8258
rect 15090 8206 15092 8258
rect 15036 7476 15092 8206
rect 15260 7700 15316 7710
rect 15372 7700 15428 11676
rect 15820 11284 15876 11294
rect 16156 11284 16212 12686
rect 16268 12404 16324 12414
rect 16380 12404 16436 14588
rect 16492 13300 16548 15262
rect 16604 15204 16660 15214
rect 16604 14530 16660 15148
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 13748 16660 14478
rect 16604 13682 16660 13692
rect 16492 13234 16548 13244
rect 16716 13074 16772 16044
rect 16836 15708 17100 15718
rect 16892 15652 16940 15708
rect 16996 15652 17044 15708
rect 16836 15642 17100 15652
rect 17052 15092 17108 15102
rect 17052 14308 17108 15036
rect 17388 14756 17444 18510
rect 17500 17444 17556 19852
rect 17612 19908 17668 19918
rect 17612 19234 17668 19852
rect 17612 19182 17614 19234
rect 17666 19182 17668 19234
rect 17612 19170 17668 19182
rect 17612 18450 17668 18462
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18116 17668 18398
rect 17612 18050 17668 18060
rect 17612 17444 17668 17454
rect 17500 17388 17612 17444
rect 17612 17378 17668 17388
rect 17500 16884 17556 16894
rect 17500 16790 17556 16828
rect 17724 15652 17780 23100
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 17836 16772 17892 21534
rect 17948 20692 18004 26852
rect 18060 26852 18116 26862
rect 18060 24834 18116 26796
rect 18060 24782 18062 24834
rect 18114 24782 18116 24834
rect 18060 24770 18116 24782
rect 18284 26852 18340 26862
rect 18284 26290 18340 26796
rect 18284 26238 18286 26290
rect 18338 26238 18340 26290
rect 18060 23268 18116 23278
rect 18060 23174 18116 23212
rect 18284 22148 18340 26238
rect 18844 26290 18900 28252
rect 19180 27860 19236 30046
rect 20188 30100 20244 30110
rect 19404 29988 19460 29998
rect 19740 29988 19796 29998
rect 19404 29650 19460 29932
rect 19404 29598 19406 29650
rect 19458 29598 19460 29650
rect 19404 29586 19460 29598
rect 19516 29986 19796 29988
rect 19516 29934 19742 29986
rect 19794 29934 19796 29986
rect 19516 29932 19796 29934
rect 19180 27794 19236 27804
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 26226 18900 26238
rect 18956 26850 19012 26862
rect 18956 26798 18958 26850
rect 19010 26798 19012 26850
rect 18956 24946 19012 26798
rect 19292 25620 19348 25630
rect 19292 25526 19348 25564
rect 18956 24894 18958 24946
rect 19010 24894 19012 24946
rect 18956 24882 19012 24894
rect 18396 24724 18452 24734
rect 18396 24630 18452 24668
rect 18956 24724 19012 24734
rect 18956 24630 19012 24668
rect 18396 23268 18452 23278
rect 18732 23268 18788 23278
rect 18396 23266 18732 23268
rect 18396 23214 18398 23266
rect 18450 23214 18732 23266
rect 18396 23212 18732 23214
rect 18396 23202 18452 23212
rect 18732 23174 18788 23212
rect 18956 23042 19012 23054
rect 18956 22990 18958 23042
rect 19010 22990 19012 23042
rect 18396 22148 18452 22158
rect 18284 22092 18396 22148
rect 18060 21812 18116 21822
rect 18060 21718 18116 21756
rect 17948 20626 18004 20636
rect 18396 21586 18452 22092
rect 18956 22146 19012 22990
rect 18956 22094 18958 22146
rect 19010 22094 19012 22146
rect 18956 22082 19012 22094
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18396 20188 18452 21534
rect 18956 21588 19012 21598
rect 18956 21494 19012 21532
rect 19516 21364 19572 29932
rect 19740 29922 19796 29932
rect 20188 29650 20244 30044
rect 20188 29598 20190 29650
rect 20242 29598 20244 29650
rect 20188 29586 20244 29598
rect 21084 29986 21140 29998
rect 21084 29934 21086 29986
rect 21138 29934 21140 29986
rect 20742 29036 21006 29046
rect 20798 28980 20846 29036
rect 20902 28980 20950 29036
rect 20742 28970 21006 28980
rect 20860 28868 20916 28878
rect 20860 28774 20916 28812
rect 19740 28644 19796 28654
rect 19740 27298 19796 28588
rect 19740 27246 19742 27298
rect 19794 27246 19796 27298
rect 19740 27234 19796 27246
rect 19964 28420 20020 28430
rect 19964 27186 20020 28364
rect 20076 28418 20132 28430
rect 20076 28366 20078 28418
rect 20130 28366 20132 28418
rect 20076 28196 20132 28366
rect 20076 28130 20132 28140
rect 21084 28084 21140 29934
rect 21308 29540 21364 29550
rect 21308 28868 21364 29484
rect 21308 28802 21364 28812
rect 21308 28532 21364 28542
rect 21308 28438 21364 28476
rect 21756 28308 21812 30270
rect 22764 30098 22820 30110
rect 22764 30046 22766 30098
rect 22818 30046 22820 30098
rect 21868 29876 21924 29886
rect 21868 28754 21924 29820
rect 22540 29426 22596 29438
rect 22540 29374 22542 29426
rect 22594 29374 22596 29426
rect 22540 29316 22596 29374
rect 22540 29250 22596 29260
rect 22652 29428 22708 29438
rect 21868 28702 21870 28754
rect 21922 28702 21924 28754
rect 21868 28690 21924 28702
rect 21756 28242 21812 28252
rect 22540 28642 22596 28654
rect 22540 28590 22542 28642
rect 22594 28590 22596 28642
rect 20636 28028 21140 28084
rect 19964 27134 19966 27186
rect 20018 27134 20020 27186
rect 19964 27122 20020 27134
rect 20076 27970 20132 27982
rect 20076 27918 20078 27970
rect 20130 27918 20132 27970
rect 20076 25732 20132 27918
rect 20636 27860 20692 28028
rect 20524 27858 20692 27860
rect 20524 27806 20638 27858
rect 20690 27806 20692 27858
rect 20524 27804 20692 27806
rect 20524 27300 20580 27804
rect 20636 27794 20692 27804
rect 21084 27858 21140 27870
rect 21084 27806 21086 27858
rect 21138 27806 21140 27858
rect 20742 27468 21006 27478
rect 20798 27412 20846 27468
rect 20902 27412 20950 27468
rect 20742 27402 21006 27412
rect 20524 27244 20804 27300
rect 20748 27186 20804 27244
rect 20748 27134 20750 27186
rect 20802 27134 20804 27186
rect 20300 26964 20356 27002
rect 20300 26898 20356 26908
rect 20748 26852 20804 27134
rect 20748 26786 20804 26796
rect 21084 26180 21140 27806
rect 21644 27860 21700 27870
rect 21644 27186 21700 27804
rect 22204 27300 22260 27310
rect 22204 27206 22260 27244
rect 21644 27134 21646 27186
rect 21698 27134 21700 27186
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 26514 21364 26910
rect 21308 26462 21310 26514
rect 21362 26462 21364 26514
rect 21308 26450 21364 26462
rect 21532 26964 21588 26974
rect 21644 26908 21700 27134
rect 21532 26852 21700 26908
rect 21756 26964 21812 26974
rect 22540 26908 22596 28590
rect 21084 26114 21140 26124
rect 20742 25900 21006 25910
rect 20798 25844 20846 25900
rect 20902 25844 20950 25900
rect 20742 25834 21006 25844
rect 20076 25666 20132 25676
rect 21532 25506 21588 26852
rect 21756 25618 21812 26908
rect 22204 26852 22596 26908
rect 21980 26404 22036 26414
rect 21980 26310 22036 26348
rect 21756 25566 21758 25618
rect 21810 25566 21812 25618
rect 21756 25554 21812 25566
rect 22092 25618 22148 25630
rect 22092 25566 22094 25618
rect 22146 25566 22148 25618
rect 21532 25454 21534 25506
rect 21586 25454 21588 25506
rect 20300 25396 20356 25406
rect 20188 25394 20356 25396
rect 20188 25342 20302 25394
rect 20354 25342 20356 25394
rect 20188 25340 20356 25342
rect 19740 24948 19796 24958
rect 19740 24854 19796 24892
rect 20188 23716 20244 25340
rect 20300 25330 20356 25340
rect 21084 25284 21140 25294
rect 20524 24836 20580 24846
rect 20524 24742 20580 24780
rect 20742 24332 21006 24342
rect 20798 24276 20846 24332
rect 20902 24276 20950 24332
rect 20742 24266 21006 24276
rect 20524 24164 20580 24174
rect 19628 23660 20244 23716
rect 20300 23828 20356 23838
rect 20300 23714 20356 23772
rect 20300 23662 20302 23714
rect 20354 23662 20356 23714
rect 19628 22594 19684 23660
rect 20300 23650 20356 23662
rect 19628 22542 19630 22594
rect 19682 22542 19684 22594
rect 19628 22530 19684 22542
rect 20524 23268 20580 24108
rect 20860 24164 20916 24174
rect 21084 24164 21140 25228
rect 21532 24724 21588 25454
rect 21532 24658 21588 24668
rect 20860 24162 21140 24164
rect 20860 24110 20862 24162
rect 20914 24110 21140 24162
rect 20860 24108 21140 24110
rect 21196 24276 21252 24286
rect 20860 24098 20916 24108
rect 20524 22370 20580 23212
rect 20860 23156 20916 23166
rect 20860 23062 20916 23100
rect 20742 22764 21006 22774
rect 20798 22708 20846 22764
rect 20902 22708 20950 22764
rect 20742 22698 21006 22708
rect 21196 22594 21252 24220
rect 21644 24164 21700 24174
rect 21644 24052 21700 24108
rect 21644 24050 21924 24052
rect 21644 23998 21646 24050
rect 21698 23998 21924 24050
rect 21644 23996 21924 23998
rect 21644 23986 21700 23996
rect 21308 23828 21364 23838
rect 21308 23734 21364 23772
rect 21196 22542 21198 22594
rect 21250 22542 21252 22594
rect 21196 22530 21252 22542
rect 20524 22318 20526 22370
rect 20578 22318 20580 22370
rect 20524 22306 20580 22318
rect 20748 22260 20804 22270
rect 20748 22258 21140 22260
rect 20748 22206 20750 22258
rect 20802 22206 21140 22258
rect 20748 22204 21140 22206
rect 20748 22194 20804 22204
rect 19964 22148 20020 22158
rect 20636 22148 20692 22158
rect 19964 22054 20020 22092
rect 20524 22092 20636 22148
rect 19516 21298 19572 21308
rect 20524 20914 20580 22092
rect 20636 22082 20692 22092
rect 21084 21812 21140 22204
rect 21196 21812 21252 21822
rect 21084 21810 21252 21812
rect 21084 21758 21198 21810
rect 21250 21758 21252 21810
rect 21084 21756 21252 21758
rect 21196 21746 21252 21756
rect 20742 21196 21006 21206
rect 20798 21140 20846 21196
rect 20902 21140 20950 21196
rect 20742 21130 21006 21140
rect 20524 20862 20526 20914
rect 20578 20862 20580 20914
rect 20524 20850 20580 20862
rect 21868 20916 21924 23996
rect 22092 23938 22148 25566
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 22484 22148 23886
rect 22204 25282 22260 26796
rect 22204 25230 22206 25282
rect 22258 25230 22260 25282
rect 22204 24724 22260 25230
rect 22316 26402 22372 26414
rect 22316 26350 22318 26402
rect 22370 26350 22372 26402
rect 22316 25284 22372 26350
rect 22652 25730 22708 29372
rect 22764 28644 22820 30046
rect 23548 30100 23604 30110
rect 23548 30006 23604 30044
rect 23884 30100 23940 30110
rect 24780 30100 24836 30110
rect 23884 30098 24052 30100
rect 23884 30046 23886 30098
rect 23938 30046 24052 30098
rect 23884 30044 24052 30046
rect 23884 30034 23940 30044
rect 23996 29652 24052 30044
rect 24780 30006 24836 30044
rect 24892 29988 24948 33200
rect 25228 30212 25284 30222
rect 25228 30118 25284 30156
rect 24892 29922 24948 29932
rect 24648 29820 24912 29830
rect 24704 29764 24752 29820
rect 24808 29764 24856 29820
rect 24648 29754 24912 29764
rect 24556 29652 24612 29662
rect 23996 29558 24052 29596
rect 24444 29596 24556 29652
rect 23100 29428 23156 29438
rect 24332 29428 24388 29438
rect 23100 29426 23492 29428
rect 23100 29374 23102 29426
rect 23154 29374 23492 29426
rect 23100 29372 23492 29374
rect 23100 29362 23156 29372
rect 22764 28578 22820 28588
rect 22876 29204 22932 29214
rect 22764 28420 22820 28430
rect 22876 28420 22932 29148
rect 22764 28418 22932 28420
rect 22764 28366 22766 28418
rect 22818 28366 22932 28418
rect 22764 28364 22932 28366
rect 23324 28980 23380 28990
rect 22764 28354 22820 28364
rect 23324 28082 23380 28924
rect 23324 28030 23326 28082
rect 23378 28030 23380 28082
rect 23324 28018 23380 28030
rect 23436 28644 23492 29372
rect 24332 29334 24388 29372
rect 22988 26964 23044 27002
rect 22988 26898 23044 26908
rect 23436 26908 23492 28588
rect 23660 29204 23716 29214
rect 23548 28532 23604 28542
rect 23660 28532 23716 29148
rect 23548 28530 23716 28532
rect 23548 28478 23550 28530
rect 23602 28478 23716 28530
rect 23548 28476 23716 28478
rect 23548 28466 23604 28476
rect 24332 28196 24388 28206
rect 24108 27972 24164 27982
rect 24108 27878 24164 27916
rect 24332 27970 24388 28140
rect 24332 27918 24334 27970
rect 24386 27918 24388 27970
rect 24332 27906 24388 27918
rect 24444 27860 24500 29596
rect 24556 29586 24612 29596
rect 25340 29428 25396 29438
rect 25340 29334 25396 29372
rect 24648 28252 24912 28262
rect 24704 28196 24752 28252
rect 24808 28196 24856 28252
rect 24648 28186 24912 28196
rect 24556 27860 24612 27870
rect 24500 27858 24612 27860
rect 24500 27806 24558 27858
rect 24610 27806 24612 27858
rect 24500 27804 24612 27806
rect 24444 27766 24500 27804
rect 24556 27794 24612 27804
rect 25228 27748 25284 27758
rect 25004 27076 25060 27086
rect 23436 26852 23604 26908
rect 23436 26180 23492 26190
rect 22652 25678 22654 25730
rect 22706 25678 22708 25730
rect 22652 25618 22708 25678
rect 22652 25566 22654 25618
rect 22706 25566 22708 25618
rect 22652 25554 22708 25566
rect 22876 26178 23492 26180
rect 22876 26126 23438 26178
rect 23490 26126 23492 26178
rect 22876 26124 23492 26126
rect 22316 25218 22372 25228
rect 22204 23044 22260 24668
rect 22876 24722 22932 26124
rect 23436 26114 23492 26124
rect 23212 25396 23268 25406
rect 22876 24670 22878 24722
rect 22930 24670 22932 24722
rect 22876 24658 22932 24670
rect 23100 25394 23268 25396
rect 23100 25342 23214 25394
rect 23266 25342 23268 25394
rect 23100 25340 23268 25342
rect 22988 24164 23044 24174
rect 22988 24070 23044 24108
rect 22316 23044 22372 23054
rect 22204 23042 22372 23044
rect 22204 22990 22318 23042
rect 22370 22990 22372 23042
rect 22204 22988 22372 22990
rect 22092 22428 22260 22484
rect 21980 22148 22036 22158
rect 21980 22146 22148 22148
rect 21980 22094 21982 22146
rect 22034 22094 22148 22146
rect 21980 22092 22148 22094
rect 21980 22082 22036 22092
rect 21980 21924 22036 21934
rect 21980 21810 22036 21868
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 21868 20822 21924 20860
rect 22092 20914 22148 22092
rect 22092 20862 22094 20914
rect 22146 20862 22148 20914
rect 22092 20850 22148 20862
rect 22204 21476 22260 22428
rect 19068 20804 19124 20814
rect 19068 20710 19124 20748
rect 22204 20804 22260 21420
rect 22316 22372 22372 22988
rect 22316 21476 22372 22316
rect 22988 22708 23044 22718
rect 22764 21476 22820 21486
rect 22316 21474 22484 21476
rect 22316 21422 22318 21474
rect 22370 21422 22484 21474
rect 22316 21420 22484 21422
rect 22316 21410 22372 21420
rect 22204 20738 22260 20748
rect 20748 20692 20804 20702
rect 21420 20692 21476 20702
rect 20748 20690 21476 20692
rect 20748 20638 20750 20690
rect 20802 20638 21422 20690
rect 21474 20638 21476 20690
rect 20748 20636 21476 20638
rect 20748 20626 20804 20636
rect 18396 20132 18564 20188
rect 18396 19908 18452 19918
rect 18396 19814 18452 19852
rect 18060 19234 18116 19246
rect 18060 19182 18062 19234
rect 18114 19182 18116 19234
rect 18060 18564 18116 19182
rect 18508 19010 18564 20132
rect 19404 20132 19460 20142
rect 19404 20038 19460 20076
rect 20300 20132 20356 20142
rect 19068 19908 19124 19918
rect 18508 18958 18510 19010
rect 18562 18958 18564 19010
rect 18060 18498 18116 18508
rect 18396 18564 18452 18574
rect 18508 18564 18564 18958
rect 18452 18508 18564 18564
rect 18396 18498 18452 18508
rect 18508 18450 18564 18508
rect 18508 18398 18510 18450
rect 18562 18398 18564 18450
rect 18172 18338 18228 18350
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 18172 18116 18228 18286
rect 18172 18050 18228 18060
rect 18508 17780 18564 18398
rect 18508 17714 18564 17724
rect 18956 19234 19012 19246
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 17836 16706 17892 16716
rect 18732 17444 18788 17454
rect 18620 16100 18676 16110
rect 18396 15876 18452 15886
rect 17724 15586 17780 15596
rect 18060 15874 18452 15876
rect 18060 15822 18398 15874
rect 18450 15822 18452 15874
rect 18060 15820 18452 15822
rect 18060 15538 18116 15820
rect 18396 15810 18452 15820
rect 18060 15486 18062 15538
rect 18114 15486 18116 15538
rect 18060 15474 18116 15486
rect 18284 15540 18340 15550
rect 18172 15428 18228 15438
rect 18172 15334 18228 15372
rect 17500 15204 17556 15242
rect 17500 15138 17556 15148
rect 17388 14690 17444 14700
rect 17164 14532 17220 14542
rect 17164 14530 17668 14532
rect 17164 14478 17166 14530
rect 17218 14478 17668 14530
rect 17164 14476 17668 14478
rect 17164 14466 17220 14476
rect 17052 14252 17444 14308
rect 16836 14140 17100 14150
rect 16892 14084 16940 14140
rect 16996 14084 17044 14140
rect 16836 14074 17100 14084
rect 17388 13970 17444 14252
rect 17388 13918 17390 13970
rect 17442 13918 17444 13970
rect 17388 13906 17444 13918
rect 16828 13524 16884 13534
rect 16828 13522 17556 13524
rect 16828 13470 16830 13522
rect 16882 13470 17556 13522
rect 16828 13468 17556 13470
rect 16828 13458 16884 13468
rect 16716 13022 16718 13074
rect 16770 13022 16772 13074
rect 16716 13010 16772 13022
rect 17500 12850 17556 13468
rect 17612 13076 17668 14476
rect 18060 13972 18116 13982
rect 18060 13878 18116 13916
rect 17724 13746 17780 13758
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13188 17780 13694
rect 18284 13746 18340 15484
rect 18620 15314 18676 16044
rect 18620 15262 18622 15314
rect 18674 15262 18676 15314
rect 18620 15148 18676 15262
rect 18284 13694 18286 13746
rect 18338 13694 18340 13746
rect 18284 13636 18340 13694
rect 18284 13570 18340 13580
rect 18508 15092 18676 15148
rect 18508 13412 18564 15092
rect 18732 13748 18788 17388
rect 18956 17220 19012 19182
rect 19068 18450 19124 19852
rect 19180 19460 19236 19470
rect 19180 19122 19236 19404
rect 19740 19234 19796 19246
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19180 19070 19182 19122
rect 19234 19070 19236 19122
rect 19180 19058 19236 19070
rect 19516 19122 19572 19134
rect 19516 19070 19518 19122
rect 19570 19070 19572 19122
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18386 19124 18398
rect 19516 17554 19572 19070
rect 19516 17502 19518 17554
rect 19570 17502 19572 17554
rect 19516 17490 19572 17502
rect 18956 17154 19012 17164
rect 19404 17108 19460 17118
rect 19404 16210 19460 17052
rect 19404 16158 19406 16210
rect 19458 16158 19460 16210
rect 19404 16146 19460 16158
rect 19628 16100 19684 16110
rect 19740 16100 19796 19182
rect 20300 17890 20356 20076
rect 20972 19906 21028 19918
rect 20972 19854 20974 19906
rect 21026 19854 21028 19906
rect 20972 19796 21028 19854
rect 21196 19908 21252 19918
rect 21196 19814 21252 19852
rect 21420 19908 21476 20636
rect 22204 20132 22260 20142
rect 22204 20038 22260 20076
rect 21420 19842 21476 19852
rect 20300 17838 20302 17890
rect 20354 17838 20356 17890
rect 20300 17826 20356 17838
rect 20524 19740 21028 19796
rect 20524 19234 20580 19740
rect 20742 19628 21006 19638
rect 20798 19572 20846 19628
rect 20902 19572 20950 19628
rect 20742 19562 21006 19572
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 19628 16098 19796 16100
rect 19628 16046 19630 16098
rect 19682 16046 19796 16098
rect 19628 16044 19796 16046
rect 20300 16098 20356 16110
rect 20300 16046 20302 16098
rect 20354 16046 20356 16098
rect 19628 15988 19684 16044
rect 19180 15874 19236 15886
rect 19180 15822 19182 15874
rect 19234 15822 19236 15874
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 18844 13748 18900 13758
rect 17724 13122 17780 13132
rect 18172 13356 18564 13412
rect 18620 13746 18900 13748
rect 18620 13694 18846 13746
rect 18898 13694 18900 13746
rect 18620 13692 18900 13694
rect 17612 13010 17668 13020
rect 17500 12798 17502 12850
rect 17554 12798 17556 12850
rect 17500 12786 17556 12798
rect 16836 12572 17100 12582
rect 16892 12516 16940 12572
rect 16996 12516 17044 12572
rect 16836 12506 17100 12516
rect 16268 12402 16436 12404
rect 16268 12350 16270 12402
rect 16322 12350 16436 12402
rect 16268 12348 16436 12350
rect 16268 12338 16324 12348
rect 17388 12292 17444 12302
rect 17388 12198 17444 12236
rect 16492 12178 16548 12190
rect 17612 12180 17668 12190
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16492 12068 16548 12126
rect 16492 12002 16548 12012
rect 17500 12178 17668 12180
rect 17500 12126 17614 12178
rect 17666 12126 17668 12178
rect 17500 12124 17668 12126
rect 15820 11282 16212 11284
rect 15820 11230 15822 11282
rect 15874 11230 16212 11282
rect 15820 11228 16212 11230
rect 15260 7698 15428 7700
rect 15260 7646 15262 7698
rect 15314 7646 15428 7698
rect 15260 7644 15428 7646
rect 15484 9044 15540 9054
rect 15260 7634 15316 7644
rect 15036 7410 15092 7420
rect 14812 7252 14868 7262
rect 14812 7250 15092 7252
rect 14812 7198 14814 7250
rect 14866 7198 15092 7250
rect 14812 7196 15092 7198
rect 14812 7186 14868 7196
rect 14588 4610 14644 4620
rect 14700 6580 14756 6590
rect 15036 6580 15092 7196
rect 14756 6524 14980 6580
rect 14700 5122 14756 6524
rect 14924 6130 14980 6524
rect 15036 6514 15092 6524
rect 15372 7140 15428 7150
rect 14924 6078 14926 6130
rect 14978 6078 14980 6130
rect 14924 6066 14980 6078
rect 15148 6468 15204 6478
rect 15148 5908 15204 6412
rect 15148 5842 15204 5852
rect 15372 5794 15428 7084
rect 15484 6802 15540 8988
rect 15820 8484 15876 11228
rect 16836 11004 17100 11014
rect 16892 10948 16940 11004
rect 16996 10948 17044 11004
rect 16836 10938 17100 10948
rect 16268 10722 16324 10734
rect 16268 10670 16270 10722
rect 16322 10670 16324 10722
rect 15820 8258 15876 8428
rect 15820 8206 15822 8258
rect 15874 8206 15876 8258
rect 15820 7700 15876 8206
rect 15820 7634 15876 7644
rect 15932 9826 15988 9838
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 15932 7588 15988 9774
rect 16268 9380 16324 10670
rect 16268 9314 16324 9324
rect 16492 10610 16548 10622
rect 16492 10558 16494 10610
rect 16546 10558 16548 10610
rect 16156 9156 16212 9166
rect 16156 9062 16212 9100
rect 16492 8932 16548 10558
rect 16836 9436 17100 9446
rect 16892 9380 16940 9436
rect 16996 9380 17044 9436
rect 16836 9370 17100 9380
rect 16492 8866 16548 8876
rect 17388 9154 17444 9166
rect 17388 9102 17390 9154
rect 17442 9102 17444 9154
rect 16940 8818 16996 8830
rect 16940 8766 16942 8818
rect 16994 8766 16996 8818
rect 15932 7522 15988 7532
rect 16268 8258 16324 8270
rect 16268 8206 16270 8258
rect 16322 8206 16324 8258
rect 15484 6750 15486 6802
rect 15538 6750 15540 6802
rect 15484 6738 15540 6750
rect 16044 7474 16100 7486
rect 16044 7422 16046 7474
rect 16098 7422 16100 7474
rect 16044 6692 16100 7422
rect 16044 6468 16100 6636
rect 16044 6402 16100 6412
rect 16156 7362 16212 7374
rect 16156 7310 16158 7362
rect 16210 7310 16212 7362
rect 16156 6020 16212 7310
rect 16268 7364 16324 8206
rect 16940 8148 16996 8766
rect 17388 8428 17444 9102
rect 16940 8082 16996 8092
rect 17164 8372 17444 8428
rect 16836 7868 17100 7878
rect 16892 7812 16940 7868
rect 16996 7812 17044 7868
rect 16836 7802 17100 7812
rect 16828 7700 16884 7710
rect 16828 7606 16884 7644
rect 16268 7298 16324 7308
rect 16716 7252 16772 7262
rect 16156 5954 16212 5964
rect 16380 6580 16436 6590
rect 16380 6018 16436 6524
rect 16716 6578 16772 7196
rect 16716 6526 16718 6578
rect 16770 6526 16772 6578
rect 16716 6514 16772 6526
rect 16836 6300 17100 6310
rect 16892 6244 16940 6300
rect 16996 6244 17044 6300
rect 16836 6234 17100 6244
rect 16380 5966 16382 6018
rect 16434 5966 16436 6018
rect 16380 5954 16436 5966
rect 15372 5742 15374 5794
rect 15426 5742 15428 5794
rect 15372 5730 15428 5742
rect 17164 5236 17220 8372
rect 17500 8260 17556 12124
rect 17612 12114 17668 12124
rect 18172 12178 18228 13356
rect 18172 12126 18174 12178
rect 18226 12126 18228 12178
rect 18172 11396 18228 12126
rect 18508 13076 18564 13086
rect 18620 13076 18676 13692
rect 18844 13682 18900 13692
rect 19068 13748 19124 15262
rect 19180 14308 19236 15822
rect 19628 15428 19684 15932
rect 19628 15362 19684 15372
rect 20076 15986 20132 15998
rect 20076 15934 20078 15986
rect 20130 15934 20132 15986
rect 19180 14242 19236 14252
rect 19628 14308 19684 14318
rect 20076 14308 20132 15934
rect 20300 15988 20356 16046
rect 20300 15922 20356 15932
rect 20524 15148 20580 19182
rect 21196 19234 21252 19246
rect 21196 19182 21198 19234
rect 21250 19182 21252 19234
rect 20748 19124 20804 19134
rect 20748 19030 20804 19068
rect 21196 18452 21252 19182
rect 21868 19236 21924 19246
rect 21868 19142 21924 19180
rect 20742 18060 21006 18070
rect 20798 18004 20846 18060
rect 20902 18004 20950 18060
rect 20742 17994 21006 18004
rect 20748 17780 20804 17790
rect 21196 17780 21252 18396
rect 20804 17724 21252 17780
rect 21308 18562 21364 18574
rect 21308 18510 21310 18562
rect 21362 18510 21364 18562
rect 21308 17778 21364 18510
rect 22428 18452 22484 21420
rect 22820 21420 22932 21476
rect 22764 21382 22820 21420
rect 22652 21364 22708 21374
rect 22540 21308 22652 21364
rect 22540 20804 22596 21308
rect 22652 21298 22708 21308
rect 22540 20802 22708 20804
rect 22540 20750 22542 20802
rect 22594 20750 22708 20802
rect 22540 20748 22708 20750
rect 22540 20738 22596 20748
rect 22428 18358 22484 18396
rect 22092 18228 22148 18238
rect 22092 18134 22148 18172
rect 21308 17726 21310 17778
rect 21362 17726 21364 17778
rect 20748 17686 20804 17724
rect 21308 17714 21364 17726
rect 21532 17724 22260 17780
rect 21532 17666 21588 17724
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 21532 17108 21588 17614
rect 22204 17666 22260 17724
rect 22204 17614 22206 17666
rect 22258 17614 22260 17666
rect 22204 17602 22260 17614
rect 22652 17666 22708 20748
rect 22876 20580 22932 21420
rect 22988 20802 23044 22652
rect 23100 21924 23156 25340
rect 23212 25330 23268 25340
rect 23212 24724 23268 24734
rect 23212 24630 23268 24668
rect 23100 21858 23156 21868
rect 23548 23938 23604 26852
rect 24108 26852 24164 26862
rect 24108 26516 24164 26796
rect 24648 26684 24912 26694
rect 24704 26628 24752 26684
rect 24808 26628 24856 26684
rect 24648 26618 24912 26628
rect 24556 26516 24612 26526
rect 24108 26514 24612 26516
rect 24108 26462 24110 26514
rect 24162 26462 24558 26514
rect 24610 26462 24612 26514
rect 24108 26460 24612 26462
rect 24108 26450 24164 26460
rect 24556 26450 24612 26460
rect 24892 25732 24948 25742
rect 24892 25638 24948 25676
rect 24332 25620 24388 25630
rect 24220 25618 24388 25620
rect 24220 25566 24334 25618
rect 24386 25566 24388 25618
rect 24220 25564 24388 25566
rect 23660 24836 23716 24846
rect 23660 24742 23716 24780
rect 23996 24836 24052 24846
rect 23996 24164 24052 24780
rect 23996 24098 24052 24108
rect 23548 23886 23550 23938
rect 23602 23886 23604 23938
rect 22988 20750 22990 20802
rect 23042 20750 23044 20802
rect 22988 20738 23044 20750
rect 23212 21474 23268 21486
rect 23212 21422 23214 21474
rect 23266 21422 23268 21474
rect 22876 20524 23156 20580
rect 22876 18450 22932 20524
rect 23100 20244 23156 20524
rect 23100 20150 23156 20188
rect 22876 18398 22878 18450
rect 22930 18398 22932 18450
rect 22876 18386 22932 18398
rect 23212 18340 23268 21422
rect 23548 21364 23604 23886
rect 23436 20244 23492 20254
rect 23436 20130 23492 20188
rect 23436 20078 23438 20130
rect 23490 20078 23492 20130
rect 23436 20066 23492 20078
rect 23548 20020 23604 21308
rect 23548 19954 23604 19964
rect 24108 23938 24164 23950
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 18340 24164 23886
rect 24220 22370 24276 25564
rect 24332 25554 24388 25564
rect 24648 25116 24912 25126
rect 24704 25060 24752 25116
rect 24808 25060 24856 25116
rect 24648 25050 24912 25060
rect 24444 24946 24500 24958
rect 24444 24894 24446 24946
rect 24498 24894 24500 24946
rect 24332 24836 24388 24846
rect 24332 24742 24388 24780
rect 24444 23044 24500 24894
rect 24648 23548 24912 23558
rect 24704 23492 24752 23548
rect 24808 23492 24856 23548
rect 24648 23482 24912 23492
rect 24444 22978 24500 22988
rect 25004 22594 25060 27020
rect 25228 27074 25284 27692
rect 25228 27022 25230 27074
rect 25282 27022 25284 27074
rect 25228 27010 25284 27022
rect 25340 27746 25396 27758
rect 25340 27694 25342 27746
rect 25394 27694 25396 27746
rect 25340 27076 25396 27694
rect 25564 27636 25620 33200
rect 25900 29988 25956 29998
rect 25900 29894 25956 29932
rect 26236 29540 26292 33200
rect 26908 31948 26964 33200
rect 26908 31892 27188 31948
rect 26348 30212 26404 30222
rect 26796 30212 26852 30222
rect 26404 30156 26516 30212
rect 26348 30146 26404 30156
rect 26236 29484 26404 29540
rect 26236 29316 26292 29326
rect 26236 29222 26292 29260
rect 25900 28868 25956 28878
rect 25900 28642 25956 28812
rect 25900 28590 25902 28642
rect 25954 28590 25956 28642
rect 25900 28578 25956 28590
rect 26236 28644 26292 28654
rect 26236 28550 26292 28588
rect 26236 27748 26292 27758
rect 26236 27654 26292 27692
rect 25564 27580 25956 27636
rect 25676 27076 25732 27086
rect 25340 27074 25732 27076
rect 25340 27022 25678 27074
rect 25730 27022 25732 27074
rect 25340 27020 25732 27022
rect 25004 22542 25006 22594
rect 25058 22542 25060 22594
rect 25004 22530 25060 22542
rect 25340 24610 25396 27020
rect 25676 27010 25732 27020
rect 25788 26964 25844 26974
rect 25340 24558 25342 24610
rect 25394 24558 25396 24610
rect 24220 22318 24222 22370
rect 24274 22318 24276 22370
rect 24220 22306 24276 22318
rect 24668 22372 24724 22382
rect 24668 22278 24724 22316
rect 25116 22372 25172 22382
rect 25340 22372 25396 24558
rect 25452 26178 25508 26190
rect 25452 26126 25454 26178
rect 25506 26126 25508 26178
rect 25452 24612 25508 26126
rect 25676 25396 25732 25406
rect 25788 25396 25844 26908
rect 25676 25394 25844 25396
rect 25676 25342 25678 25394
rect 25730 25342 25844 25394
rect 25676 25340 25844 25342
rect 25676 25330 25732 25340
rect 25788 24612 25844 24622
rect 25452 24610 25844 24612
rect 25452 24558 25790 24610
rect 25842 24558 25844 24610
rect 25452 24556 25844 24558
rect 25788 23156 25844 24556
rect 25788 23090 25844 23100
rect 25172 22316 25396 22372
rect 25676 23044 25732 23054
rect 25116 22306 25172 22316
rect 24648 21980 24912 21990
rect 24704 21924 24752 21980
rect 24808 21924 24856 21980
rect 24648 21914 24912 21924
rect 25116 21924 25172 21934
rect 25116 21810 25172 21868
rect 25116 21758 25118 21810
rect 25170 21758 25172 21810
rect 25116 21746 25172 21758
rect 24444 21698 24500 21710
rect 24444 21646 24446 21698
rect 24498 21646 24500 21698
rect 24332 19906 24388 19918
rect 24332 19854 24334 19906
rect 24386 19854 24388 19906
rect 24332 19796 24388 19854
rect 24332 19730 24388 19740
rect 24332 19010 24388 19022
rect 24332 18958 24334 19010
rect 24386 18958 24388 19010
rect 24332 18562 24388 18958
rect 24444 18676 24500 21646
rect 24648 20412 24912 20422
rect 24704 20356 24752 20412
rect 24808 20356 24856 20412
rect 24648 20346 24912 20356
rect 25228 20132 25284 22316
rect 25564 22148 25620 22158
rect 25564 22054 25620 22092
rect 25676 21810 25732 22988
rect 25676 21758 25678 21810
rect 25730 21758 25732 21810
rect 25676 21746 25732 21758
rect 25788 20692 25844 20702
rect 25564 20580 25620 20590
rect 25788 20580 25844 20636
rect 25564 20578 25844 20580
rect 25564 20526 25566 20578
rect 25618 20526 25844 20578
rect 25564 20524 25844 20526
rect 25564 20514 25620 20524
rect 25340 20132 25396 20142
rect 25228 20130 25396 20132
rect 25228 20078 25342 20130
rect 25394 20078 25396 20130
rect 25228 20076 25396 20078
rect 25340 20066 25396 20076
rect 25004 20020 25060 20030
rect 24892 19460 24948 19470
rect 24892 19366 24948 19404
rect 25004 19234 25060 19964
rect 25564 20020 25620 20030
rect 25564 19926 25620 19964
rect 25004 19182 25006 19234
rect 25058 19182 25060 19234
rect 25004 19170 25060 19182
rect 25564 19796 25620 19806
rect 24648 18844 24912 18854
rect 24704 18788 24752 18844
rect 24808 18788 24856 18844
rect 24648 18778 24912 18788
rect 24444 18620 25060 18676
rect 24332 18510 24334 18562
rect 24386 18510 24388 18562
rect 24332 18498 24388 18510
rect 24556 18450 24612 18462
rect 24556 18398 24558 18450
rect 24610 18398 24612 18450
rect 24108 18284 24500 18340
rect 23212 18274 23268 18284
rect 23324 18226 23380 18238
rect 23324 18174 23326 18226
rect 23378 18174 23380 18226
rect 23324 18116 23380 18174
rect 23324 17892 23380 18060
rect 22652 17614 22654 17666
rect 22706 17614 22708 17666
rect 22652 17602 22708 17614
rect 23212 17836 23380 17892
rect 21980 17556 22036 17566
rect 21308 17052 21588 17108
rect 21756 17554 22036 17556
rect 21756 17502 21982 17554
rect 22034 17502 22036 17554
rect 21756 17500 22036 17502
rect 20742 16492 21006 16502
rect 20798 16436 20846 16492
rect 20902 16436 20950 16492
rect 20742 16426 21006 16436
rect 21308 15988 21364 17052
rect 21756 16996 21812 17500
rect 21980 17490 22036 17500
rect 21532 16940 21812 16996
rect 22540 17220 22596 17230
rect 21420 16100 21476 16110
rect 21420 16006 21476 16044
rect 21308 15922 21364 15932
rect 21532 15538 21588 16940
rect 21532 15486 21534 15538
rect 21586 15486 21588 15538
rect 21532 15474 21588 15486
rect 21644 16770 21700 16782
rect 21644 16718 21646 16770
rect 21698 16718 21700 16770
rect 20524 15092 21140 15148
rect 20412 14980 20468 14990
rect 20412 14418 20468 14924
rect 20742 14924 21006 14934
rect 20798 14868 20846 14924
rect 20902 14868 20950 14924
rect 20742 14858 21006 14868
rect 20412 14366 20414 14418
rect 20466 14366 20468 14418
rect 20412 14354 20468 14366
rect 20748 14420 20804 14430
rect 19628 14306 20132 14308
rect 19628 14254 19630 14306
rect 19682 14254 20132 14306
rect 19628 14252 20132 14254
rect 20188 14306 20244 14318
rect 20188 14254 20190 14306
rect 20242 14254 20244 14306
rect 19628 14242 19684 14252
rect 19068 13682 19124 13692
rect 18508 13074 18676 13076
rect 18508 13022 18510 13074
rect 18562 13022 18676 13074
rect 18508 13020 18676 13022
rect 18956 13636 19012 13646
rect 18956 13074 19012 13580
rect 18956 13022 18958 13074
rect 19010 13022 19012 13074
rect 18508 11732 18564 13020
rect 18956 13010 19012 13022
rect 19292 13076 19348 13086
rect 19292 12982 19348 13020
rect 20188 12292 20244 14254
rect 20524 14308 20580 14318
rect 20524 12850 20580 14252
rect 20748 13860 20804 14364
rect 20748 13794 20804 13804
rect 20742 13356 21006 13366
rect 20798 13300 20846 13356
rect 20902 13300 20950 13356
rect 20742 13290 21006 13300
rect 20524 12798 20526 12850
rect 20578 12798 20580 12850
rect 20524 12786 20580 12798
rect 20860 12292 20916 12302
rect 20188 12226 20244 12236
rect 20412 12290 20916 12292
rect 20412 12238 20862 12290
rect 20914 12238 20916 12290
rect 20412 12236 20916 12238
rect 18508 11666 18564 11676
rect 18620 12178 18676 12190
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 11620 18676 12126
rect 18956 11620 19012 11630
rect 18620 11618 19012 11620
rect 18620 11566 18958 11618
rect 19010 11566 19012 11618
rect 18620 11564 19012 11566
rect 18956 11554 19012 11564
rect 20412 11618 20468 12236
rect 20860 12226 20916 12236
rect 20742 11788 21006 11798
rect 20798 11732 20846 11788
rect 20902 11732 20950 11788
rect 20742 11722 21006 11732
rect 20412 11566 20414 11618
rect 20466 11566 20468 11618
rect 20412 11554 20468 11566
rect 19180 11508 19236 11518
rect 18228 11340 18340 11396
rect 18172 11330 18228 11340
rect 18172 10612 18228 10622
rect 18172 10518 18228 10556
rect 18060 10386 18116 10398
rect 18060 10334 18062 10386
rect 18114 10334 18116 10386
rect 18060 9716 18116 10334
rect 18172 9716 18228 9726
rect 18060 9714 18228 9716
rect 18060 9662 18174 9714
rect 18226 9662 18228 9714
rect 18060 9660 18228 9662
rect 18172 9650 18228 9660
rect 17724 9604 17780 9614
rect 17724 9154 17780 9548
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17724 9090 17780 9102
rect 18284 9044 18340 11340
rect 19180 11172 19236 11452
rect 19180 11078 19236 11116
rect 19740 11394 19796 11406
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19068 10724 19124 10734
rect 18956 10498 19012 10510
rect 18956 10446 18958 10498
rect 19010 10446 19012 10498
rect 18956 10276 19012 10446
rect 18844 10220 19012 10276
rect 18844 9828 18900 10220
rect 18956 10052 19012 10062
rect 19068 10052 19124 10668
rect 19404 10612 19460 10622
rect 19404 10518 19460 10556
rect 19740 10500 19796 11342
rect 20524 11394 20580 11406
rect 20524 11342 20526 11394
rect 20578 11342 20580 11394
rect 19964 10500 20020 10510
rect 19740 10498 20020 10500
rect 19740 10446 19966 10498
rect 20018 10446 20020 10498
rect 19740 10444 20020 10446
rect 19964 10434 20020 10444
rect 20524 10500 20580 11342
rect 21084 11284 21140 15092
rect 21532 14530 21588 14542
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21420 13860 21476 13870
rect 21420 13074 21476 13804
rect 21420 13022 21422 13074
rect 21474 13022 21476 13074
rect 21420 13010 21476 13022
rect 21196 11396 21252 11406
rect 21196 11302 21252 11340
rect 21084 11218 21140 11228
rect 20972 10724 21028 10734
rect 20972 10630 21028 10668
rect 20524 10434 20580 10444
rect 20742 10220 21006 10230
rect 20798 10164 20846 10220
rect 20902 10164 20950 10220
rect 20742 10154 21006 10164
rect 18956 10050 19124 10052
rect 18956 9998 18958 10050
rect 19010 9998 19124 10050
rect 18956 9996 19124 9998
rect 21532 10052 21588 14478
rect 21644 13188 21700 16718
rect 21868 16098 21924 16110
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21868 14980 21924 16046
rect 21868 14914 21924 14924
rect 21980 16100 22036 16110
rect 21980 14530 22036 16044
rect 22540 15538 22596 17164
rect 22988 16994 23044 17006
rect 22988 16942 22990 16994
rect 23042 16942 23044 16994
rect 22988 16772 23044 16942
rect 22988 16706 23044 16716
rect 23100 16660 23156 16670
rect 22540 15486 22542 15538
rect 22594 15486 22596 15538
rect 22540 15474 22596 15486
rect 22652 16212 22708 16222
rect 22092 15092 22148 15102
rect 22092 14998 22148 15036
rect 21980 14478 21982 14530
rect 22034 14478 22036 14530
rect 21980 14466 22036 14478
rect 22652 14530 22708 16156
rect 22876 15428 22932 15438
rect 23100 15428 23156 16604
rect 22876 15426 23156 15428
rect 22876 15374 22878 15426
rect 22930 15374 23156 15426
rect 22876 15372 23156 15374
rect 22876 15362 22932 15372
rect 22652 14478 22654 14530
rect 22706 14478 22708 14530
rect 22652 14466 22708 14478
rect 21756 14420 21812 14430
rect 21756 14326 21812 14364
rect 23100 13972 23156 15372
rect 23212 15988 23268 17836
rect 23324 17668 23380 17678
rect 23324 17574 23380 17612
rect 23660 17108 23716 17118
rect 23324 16996 23380 17006
rect 23324 16902 23380 16940
rect 23660 16994 23716 17052
rect 24332 17108 24388 17118
rect 23996 16996 24052 17006
rect 24332 16996 24388 17052
rect 23660 16942 23662 16994
rect 23714 16942 23716 16994
rect 23660 16930 23716 16942
rect 23884 16940 23996 16996
rect 23212 15426 23268 15932
rect 23212 15374 23214 15426
rect 23266 15374 23268 15426
rect 23212 15362 23268 15374
rect 23548 15876 23604 15886
rect 23548 15426 23604 15820
rect 23548 15374 23550 15426
rect 23602 15374 23604 15426
rect 23548 15362 23604 15374
rect 23884 15148 23940 16940
rect 23996 16930 24052 16940
rect 24108 16994 24388 16996
rect 24108 16942 24334 16994
rect 24386 16942 24388 16994
rect 24108 16940 24388 16942
rect 23996 16772 24052 16782
rect 23996 16678 24052 16716
rect 24108 16100 24164 16940
rect 24332 16930 24388 16940
rect 23996 16044 24164 16100
rect 23996 15540 24052 16044
rect 24108 15876 24164 15886
rect 24108 15782 24164 15820
rect 24332 15652 24388 15662
rect 24108 15540 24164 15550
rect 23996 15538 24164 15540
rect 23996 15486 24110 15538
rect 24162 15486 24164 15538
rect 23996 15484 24164 15486
rect 24108 15474 24164 15484
rect 24332 15426 24388 15596
rect 24332 15374 24334 15426
rect 24386 15374 24388 15426
rect 24332 15362 24388 15374
rect 23884 15092 24052 15148
rect 23324 13972 23380 13982
rect 23100 13970 23380 13972
rect 23100 13918 23326 13970
rect 23378 13918 23380 13970
rect 23100 13916 23380 13918
rect 23996 13972 24052 15092
rect 24444 14644 24500 18284
rect 24556 18116 24612 18398
rect 24556 18050 24612 18060
rect 24648 17276 24912 17286
rect 24704 17220 24752 17276
rect 24808 17220 24856 17276
rect 24648 17210 24912 17220
rect 24668 16770 24724 16782
rect 24668 16718 24670 16770
rect 24722 16718 24724 16770
rect 24668 16100 24724 16718
rect 25004 16322 25060 18620
rect 25564 18450 25620 19740
rect 25676 19236 25732 19246
rect 25676 19234 25844 19236
rect 25676 19182 25678 19234
rect 25730 19182 25844 19234
rect 25676 19180 25844 19182
rect 25676 19170 25732 19180
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25564 18340 25620 18398
rect 25564 18274 25620 18284
rect 25676 18338 25732 18350
rect 25676 18286 25678 18338
rect 25730 18286 25732 18338
rect 25452 18116 25508 18126
rect 25340 16884 25396 16894
rect 25340 16790 25396 16828
rect 25004 16270 25006 16322
rect 25058 16270 25060 16322
rect 25004 16258 25060 16270
rect 24668 16034 24724 16044
rect 24892 15988 24948 15998
rect 24892 15894 24948 15932
rect 24648 15708 24912 15718
rect 24704 15652 24752 15708
rect 24808 15652 24856 15708
rect 24648 15642 24912 15652
rect 24668 15428 24724 15438
rect 24668 15334 24724 15372
rect 25452 15314 25508 18060
rect 25676 17442 25732 18286
rect 25788 17780 25844 19180
rect 25788 17714 25844 17724
rect 25676 17390 25678 17442
rect 25730 17390 25732 17442
rect 25676 17378 25732 17390
rect 25900 16996 25956 27580
rect 26348 27524 26404 29484
rect 25900 16930 25956 16940
rect 26012 27468 26404 27524
rect 25788 16882 25844 16894
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 25564 16772 25620 16782
rect 25564 15874 25620 16716
rect 25788 16772 25844 16830
rect 25788 16706 25844 16716
rect 25564 15822 25566 15874
rect 25618 15822 25620 15874
rect 25564 15810 25620 15822
rect 25452 15262 25454 15314
rect 25506 15262 25508 15314
rect 25452 15250 25508 15262
rect 25676 15652 25732 15662
rect 25228 15202 25284 15214
rect 25228 15150 25230 15202
rect 25282 15150 25284 15202
rect 25228 15148 25284 15150
rect 25116 15092 25284 15148
rect 24556 14644 24612 14654
rect 24444 14588 24556 14644
rect 24556 14578 24612 14588
rect 25116 14306 25172 15092
rect 25676 14754 25732 15596
rect 25676 14702 25678 14754
rect 25730 14702 25732 14754
rect 25676 14690 25732 14702
rect 26012 15428 26068 27468
rect 26460 26908 26516 30156
rect 26684 30098 26740 30110
rect 26684 30046 26686 30098
rect 26738 30046 26740 30098
rect 26684 28980 26740 30046
rect 26684 28914 26740 28924
rect 26796 28530 26852 30156
rect 26908 30210 26964 30222
rect 26908 30158 26910 30210
rect 26962 30158 26964 30210
rect 26908 29652 26964 30158
rect 26908 29586 26964 29596
rect 27132 28756 27188 31892
rect 27580 30212 27636 33200
rect 27580 30146 27636 30156
rect 27356 30098 27412 30110
rect 27356 30046 27358 30098
rect 27410 30046 27412 30098
rect 27356 29652 27412 30046
rect 28252 30100 28308 33200
rect 28924 31948 28980 33200
rect 28924 31892 29204 31948
rect 28554 30604 28818 30614
rect 28610 30548 28658 30604
rect 28714 30548 28762 30604
rect 28554 30538 28818 30548
rect 28252 30034 28308 30044
rect 28476 30098 28532 30110
rect 28476 30046 28478 30098
rect 28530 30046 28532 30098
rect 27356 29586 27412 29596
rect 27468 29986 27524 29998
rect 27468 29934 27470 29986
rect 27522 29934 27524 29986
rect 27244 29540 27300 29550
rect 27244 29446 27300 29484
rect 27468 29204 27524 29934
rect 28476 29876 28532 30046
rect 28812 30100 28868 30110
rect 28812 30098 28980 30100
rect 28812 30046 28814 30098
rect 28866 30046 28980 30098
rect 28812 30044 28980 30046
rect 28812 30034 28868 30044
rect 27468 29138 27524 29148
rect 27804 29820 28532 29876
rect 27580 28756 27636 28766
rect 27132 28754 27636 28756
rect 27132 28702 27582 28754
rect 27634 28702 27636 28754
rect 27132 28700 27636 28702
rect 27580 28690 27636 28700
rect 27804 28532 27860 29820
rect 28028 29652 28084 29662
rect 26796 28478 26798 28530
rect 26850 28478 26852 28530
rect 26796 28466 26852 28478
rect 27468 28476 27860 28532
rect 27916 29596 28028 29652
rect 27132 28420 27188 28430
rect 27020 28418 27188 28420
rect 27020 28366 27134 28418
rect 27186 28366 27188 28418
rect 27020 28364 27188 28366
rect 26348 26852 26516 26908
rect 26572 26962 26628 26974
rect 26572 26910 26574 26962
rect 26626 26910 26628 26962
rect 26236 26180 26292 26190
rect 26236 26086 26292 26124
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 22708 26292 24558
rect 26236 22642 26292 22652
rect 26348 21812 26404 26852
rect 26572 25284 26628 26910
rect 26572 25218 26628 25228
rect 26684 25620 26740 25630
rect 26572 24612 26628 24622
rect 26572 23714 26628 24556
rect 26572 23662 26574 23714
rect 26626 23662 26628 23714
rect 26572 23650 26628 23662
rect 26684 23492 26740 25564
rect 26348 21746 26404 21756
rect 26572 23436 26740 23492
rect 26348 20692 26404 20702
rect 26348 20598 26404 20636
rect 26124 20580 26180 20590
rect 26124 20486 26180 20524
rect 26236 20020 26292 20030
rect 26572 20020 26628 23436
rect 27020 23380 27076 28364
rect 27132 28354 27188 28364
rect 27244 27972 27300 27982
rect 27244 27878 27300 27916
rect 27468 26908 27524 28476
rect 27356 26852 27524 26908
rect 27580 27186 27636 27198
rect 27580 27134 27582 27186
rect 27634 27134 27636 27186
rect 27244 26404 27300 26414
rect 27244 26310 27300 26348
rect 27132 25284 27188 25294
rect 27132 24162 27188 25228
rect 27244 24834 27300 24846
rect 27244 24782 27246 24834
rect 27298 24782 27300 24834
rect 27244 24276 27300 24782
rect 27244 24210 27300 24220
rect 27132 24110 27134 24162
rect 27186 24110 27188 24162
rect 27132 24098 27188 24110
rect 27356 23940 27412 26852
rect 27580 25508 27636 27134
rect 27916 26908 27972 29596
rect 28028 29586 28084 29596
rect 28140 29650 28196 29820
rect 28140 29598 28142 29650
rect 28194 29598 28196 29650
rect 28140 29586 28196 29598
rect 28554 29036 28818 29046
rect 28610 28980 28658 29036
rect 28714 28980 28762 29036
rect 28554 28970 28818 28980
rect 28588 28532 28644 28542
rect 28588 27860 28644 28476
rect 28924 28084 28980 30044
rect 29036 29314 29092 29326
rect 29036 29262 29038 29314
rect 29090 29262 29092 29314
rect 29036 28868 29092 29262
rect 29036 28802 29092 28812
rect 28924 28018 28980 28028
rect 29036 28644 29092 28654
rect 28588 27858 28980 27860
rect 28588 27806 28590 27858
rect 28642 27806 28980 27858
rect 28588 27804 28980 27806
rect 28588 27794 28644 27804
rect 28028 27746 28084 27758
rect 28028 27694 28030 27746
rect 28082 27694 28084 27746
rect 28028 27524 28084 27694
rect 28364 27746 28420 27758
rect 28364 27694 28366 27746
rect 28418 27694 28420 27746
rect 28028 27468 28308 27524
rect 27916 26852 28084 26908
rect 27916 25508 27972 25518
rect 27580 25506 27972 25508
rect 27580 25454 27918 25506
rect 27970 25454 27972 25506
rect 27580 25452 27972 25454
rect 27916 25442 27972 25452
rect 27916 25284 27972 25294
rect 27804 25228 27916 25284
rect 27804 24050 27860 25228
rect 27916 25218 27972 25228
rect 28028 24836 28084 26852
rect 27804 23998 27806 24050
rect 27858 23998 27860 24050
rect 27804 23986 27860 23998
rect 27916 24780 28084 24836
rect 28252 24836 28308 27468
rect 28364 26964 28420 27694
rect 28554 27468 28818 27478
rect 28610 27412 28658 27468
rect 28714 27412 28762 27468
rect 28554 27402 28818 27412
rect 28924 26908 28980 27804
rect 28364 26898 28420 26908
rect 28476 26852 28980 26908
rect 28364 26292 28420 26302
rect 28476 26292 28532 26852
rect 28364 26290 28532 26292
rect 28364 26238 28366 26290
rect 28418 26238 28532 26290
rect 28364 26236 28532 26238
rect 28812 26628 28868 26638
rect 28812 26290 28868 26572
rect 28812 26238 28814 26290
rect 28866 26238 28868 26290
rect 28364 25508 28420 26236
rect 28812 26226 28868 26238
rect 28554 25900 28818 25910
rect 28610 25844 28658 25900
rect 28714 25844 28762 25900
rect 28554 25834 28818 25844
rect 28364 25506 28644 25508
rect 28364 25454 28366 25506
rect 28418 25454 28644 25506
rect 28364 25452 28644 25454
rect 28364 25442 28420 25452
rect 27020 23314 27076 23324
rect 27132 23884 27412 23940
rect 26684 23156 26740 23166
rect 26740 23100 26852 23156
rect 26684 23062 26740 23100
rect 26684 20916 26740 20926
rect 26684 20822 26740 20860
rect 26236 20018 26628 20020
rect 26236 19966 26238 20018
rect 26290 19966 26628 20018
rect 26236 19964 26628 19966
rect 26236 19954 26292 19964
rect 26684 18564 26740 18574
rect 26684 18470 26740 18508
rect 26460 18450 26516 18462
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26124 18340 26180 18350
rect 26124 17108 26180 18284
rect 26460 18340 26516 18398
rect 26460 18274 26516 18284
rect 26572 18116 26628 18126
rect 26572 17778 26628 18060
rect 26572 17726 26574 17778
rect 26626 17726 26628 17778
rect 26572 17714 26628 17726
rect 26348 17556 26404 17566
rect 26348 17462 26404 17500
rect 26124 15538 26180 17052
rect 26124 15486 26126 15538
rect 26178 15486 26180 15538
rect 26124 15474 26180 15486
rect 26012 14644 26068 15372
rect 26796 15148 26852 23100
rect 27132 18450 27188 23884
rect 27356 23716 27412 23726
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 27132 18340 27188 18398
rect 27132 17668 27188 18284
rect 27132 17602 27188 17612
rect 27244 23714 27412 23716
rect 27244 23662 27358 23714
rect 27410 23662 27412 23714
rect 27244 23660 27412 23662
rect 26908 17554 26964 17566
rect 26908 17502 26910 17554
rect 26962 17502 26964 17554
rect 26908 17108 26964 17502
rect 26908 17042 26964 17052
rect 26908 16100 26964 16110
rect 26908 15538 26964 16044
rect 26908 15486 26910 15538
rect 26962 15486 26964 15538
rect 26908 15474 26964 15486
rect 26348 15090 26404 15102
rect 26348 15038 26350 15090
rect 26402 15038 26404 15090
rect 26124 14644 26180 14654
rect 26012 14642 26180 14644
rect 26012 14590 26126 14642
rect 26178 14590 26180 14642
rect 26012 14588 26180 14590
rect 26124 14578 26180 14588
rect 25116 14254 25118 14306
rect 25170 14254 25172 14306
rect 25116 14242 25172 14254
rect 24648 14140 24912 14150
rect 24704 14084 24752 14140
rect 24808 14084 24856 14140
rect 24648 14074 24912 14084
rect 24108 13972 24164 13982
rect 23996 13970 24164 13972
rect 23996 13918 24110 13970
rect 24162 13918 24164 13970
rect 23996 13916 24164 13918
rect 23324 13906 23380 13916
rect 24108 13906 24164 13916
rect 22876 13748 22932 13758
rect 22540 13636 22596 13646
rect 21868 13188 21924 13198
rect 21644 13132 21868 13188
rect 21644 11954 21700 11966
rect 21644 11902 21646 11954
rect 21698 11902 21700 11954
rect 21644 10724 21700 11902
rect 21756 11732 21812 13132
rect 21868 13074 21924 13132
rect 21868 13022 21870 13074
rect 21922 13022 21924 13074
rect 21868 13010 21924 13022
rect 21756 11666 21812 11676
rect 21868 11396 21924 11406
rect 21868 11394 22036 11396
rect 21868 11342 21870 11394
rect 21922 11342 22036 11394
rect 21868 11340 22036 11342
rect 21868 11330 21924 11340
rect 21644 10658 21700 10668
rect 18956 9986 19012 9996
rect 21532 9986 21588 9996
rect 21868 10500 21924 10510
rect 21980 10500 22036 11340
rect 22316 10836 22372 10846
rect 22540 10836 22596 13580
rect 22876 12066 22932 13692
rect 25676 13746 25732 13758
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 24668 13636 24724 13646
rect 24668 13542 24724 13580
rect 25676 13636 25732 13694
rect 25676 13570 25732 13580
rect 26348 13636 26404 15038
rect 26348 13570 26404 13580
rect 26460 15092 26852 15148
rect 26460 14642 26516 15092
rect 26460 14590 26462 14642
rect 26514 14590 26516 14642
rect 26460 13746 26516 14590
rect 26796 14980 26852 14990
rect 26796 14644 26852 14924
rect 26908 14644 26964 14654
rect 26796 14642 26964 14644
rect 26796 14590 26910 14642
rect 26962 14590 26964 14642
rect 26796 14588 26964 14590
rect 26908 14578 26964 14588
rect 27244 14420 27300 23660
rect 27356 23650 27412 23660
rect 27916 20914 27972 24780
rect 28252 24724 28308 24780
rect 28028 24668 28308 24724
rect 28588 24724 28644 25452
rect 29036 25284 29092 28588
rect 29148 28532 29204 31892
rect 32284 31668 32340 31678
rect 29932 30996 29988 31006
rect 29820 30940 29932 30996
rect 29148 28466 29204 28476
rect 29260 30770 29316 30782
rect 29260 30718 29262 30770
rect 29314 30718 29316 30770
rect 29036 25218 29092 25228
rect 29148 28308 29204 28318
rect 28588 24722 28980 24724
rect 28588 24670 28590 24722
rect 28642 24670 28980 24722
rect 28588 24668 28980 24670
rect 28028 24610 28084 24668
rect 28588 24658 28644 24668
rect 28028 24558 28030 24610
rect 28082 24558 28084 24610
rect 28028 24546 28084 24558
rect 28364 24612 28420 24622
rect 28364 24518 28420 24556
rect 28554 24332 28818 24342
rect 28610 24276 28658 24332
rect 28714 24276 28762 24332
rect 28554 24266 28818 24276
rect 28924 23266 28980 24668
rect 28924 23214 28926 23266
rect 28978 23214 28980 23266
rect 28554 22764 28818 22774
rect 28610 22708 28658 22764
rect 28714 22708 28762 22764
rect 28554 22698 28818 22708
rect 28140 22484 28196 22494
rect 28140 22370 28196 22428
rect 28140 22318 28142 22370
rect 28194 22318 28196 22370
rect 28140 22306 28196 22318
rect 28700 22372 28756 22382
rect 28924 22372 28980 23214
rect 28700 22370 28980 22372
rect 28700 22318 28702 22370
rect 28754 22318 28980 22370
rect 28700 22316 28980 22318
rect 28252 21586 28308 21598
rect 28252 21534 28254 21586
rect 28306 21534 28308 21586
rect 28252 21476 28308 21534
rect 28700 21586 28756 22316
rect 28700 21534 28702 21586
rect 28754 21534 28756 21586
rect 28700 21522 28756 21534
rect 28252 21410 28308 21420
rect 28554 21196 28818 21206
rect 28610 21140 28658 21196
rect 28714 21140 28762 21196
rect 28554 21130 28818 21140
rect 27916 20862 27918 20914
rect 27970 20862 27972 20914
rect 27916 20850 27972 20862
rect 29148 20692 29204 28252
rect 29260 27858 29316 30718
rect 29260 27806 29262 27858
rect 29314 27806 29316 27858
rect 29260 27794 29316 27806
rect 29372 27636 29428 27646
rect 29372 26850 29428 27580
rect 29708 26964 29764 26974
rect 29372 26798 29374 26850
rect 29426 26798 29428 26850
rect 29372 26786 29428 26798
rect 29596 26908 29708 26964
rect 29260 25844 29316 25854
rect 29260 24722 29316 25788
rect 29260 24670 29262 24722
rect 29314 24670 29316 24722
rect 29260 24658 29316 24670
rect 29596 21140 29652 26908
rect 29708 26898 29764 26908
rect 29820 26908 29876 30940
rect 29932 30930 29988 30940
rect 30156 30770 30212 30782
rect 30156 30718 30158 30770
rect 30210 30718 30212 30770
rect 30156 30322 30212 30718
rect 30156 30270 30158 30322
rect 30210 30270 30212 30322
rect 30156 30258 30212 30270
rect 32060 30324 32116 30334
rect 31276 30098 31332 30110
rect 31276 30046 31278 30098
rect 31330 30046 31332 30098
rect 30268 29538 30324 29550
rect 30268 29486 30270 29538
rect 30322 29486 30324 29538
rect 30156 28754 30212 28766
rect 30156 28702 30158 28754
rect 30210 28702 30212 28754
rect 30156 26908 30212 28702
rect 30268 27300 30324 29486
rect 30268 27234 30324 27244
rect 30940 29426 30996 29438
rect 30940 29374 30942 29426
rect 30994 29374 30996 29426
rect 30940 29316 30996 29374
rect 29820 26852 29988 26908
rect 29708 26180 29764 26190
rect 29708 21364 29764 26124
rect 29708 21308 29876 21364
rect 29148 20626 29204 20636
rect 29372 21084 29652 21140
rect 27356 20578 27412 20590
rect 27356 20526 27358 20578
rect 27410 20526 27412 20578
rect 27356 19572 27412 20526
rect 28476 20244 28532 20254
rect 28476 20130 28532 20188
rect 28476 20078 28478 20130
rect 28530 20078 28532 20130
rect 28476 20066 28532 20078
rect 29260 20132 29316 20142
rect 29372 20132 29428 21084
rect 29820 21028 29876 21308
rect 29932 21252 29988 26852
rect 30044 26852 30212 26908
rect 30716 27186 30772 27198
rect 30716 27134 30718 27186
rect 30770 27134 30772 27186
rect 30044 26628 30100 26852
rect 30044 26562 30100 26572
rect 30716 25844 30772 27134
rect 30716 25778 30772 25788
rect 30156 25620 30212 25630
rect 30156 25526 30212 25564
rect 30156 24052 30212 24062
rect 30044 24050 30212 24052
rect 30044 23998 30158 24050
rect 30210 23998 30212 24050
rect 30044 23996 30212 23998
rect 30044 21812 30100 23996
rect 30156 23986 30212 23996
rect 30156 22484 30212 22494
rect 30156 22390 30212 22428
rect 30044 21746 30100 21756
rect 30044 21476 30100 21486
rect 30044 21382 30100 21420
rect 29932 21196 30100 21252
rect 29820 20972 29988 21028
rect 29260 20130 29428 20132
rect 29260 20078 29262 20130
rect 29314 20078 29428 20130
rect 29260 20076 29428 20078
rect 29484 20690 29540 20702
rect 29484 20638 29486 20690
rect 29538 20638 29540 20690
rect 29260 20066 29316 20076
rect 28554 19628 28818 19638
rect 28610 19572 28658 19628
rect 28714 19572 28762 19628
rect 28554 19562 28818 19572
rect 27356 19506 27412 19516
rect 28700 19236 28756 19246
rect 28700 19142 28756 19180
rect 29484 19236 29540 20638
rect 29484 19170 29540 19180
rect 27916 19012 27972 19022
rect 27356 19010 27972 19012
rect 27356 18958 27918 19010
rect 27970 18958 27972 19010
rect 27356 18956 27972 18958
rect 27356 18562 27412 18956
rect 27916 18946 27972 18956
rect 29260 19010 29316 19022
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 28140 18676 28196 18686
rect 28140 18582 28196 18620
rect 27356 18510 27358 18562
rect 27410 18510 27412 18562
rect 27356 18498 27412 18510
rect 29148 18452 29204 18462
rect 27580 18340 27636 18350
rect 27580 18246 27636 18284
rect 28554 18060 28818 18070
rect 28610 18004 28658 18060
rect 28714 18004 28762 18060
rect 28554 17994 28818 18004
rect 27356 17668 27412 17678
rect 27356 17574 27412 17612
rect 28588 17666 28644 17678
rect 28588 17614 28590 17666
rect 28642 17614 28644 17666
rect 28364 17554 28420 17566
rect 28364 17502 28366 17554
rect 28418 17502 28420 17554
rect 28028 17108 28084 17118
rect 28028 17014 28084 17052
rect 28140 16098 28196 16110
rect 28140 16046 28142 16098
rect 28194 16046 28196 16098
rect 27244 14354 27300 14364
rect 27916 15092 27972 15102
rect 27916 14418 27972 15036
rect 27916 14366 27918 14418
rect 27970 14366 27972 14418
rect 27916 14354 27972 14366
rect 28140 14084 28196 16046
rect 28140 14018 28196 14028
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 25900 13522 25956 13534
rect 25900 13470 25902 13522
rect 25954 13470 25956 13522
rect 22876 12014 22878 12066
rect 22930 12014 22932 12066
rect 22876 12002 22932 12014
rect 23660 12850 23716 12862
rect 23660 12798 23662 12850
rect 23714 12798 23716 12850
rect 23100 11172 23156 11182
rect 22316 10834 23044 10836
rect 22316 10782 22318 10834
rect 22370 10782 23044 10834
rect 22316 10780 23044 10782
rect 22316 10770 22372 10780
rect 22876 10500 22932 10510
rect 21980 10498 22932 10500
rect 21980 10446 22878 10498
rect 22930 10446 22932 10498
rect 21980 10444 22932 10446
rect 18956 9828 19012 9838
rect 18844 9772 18956 9828
rect 18956 9762 19012 9772
rect 19404 9828 19460 9838
rect 19404 9734 19460 9772
rect 20748 9828 20804 9838
rect 20748 9734 20804 9772
rect 21532 9828 21588 9838
rect 21868 9828 21924 10444
rect 22876 10434 22932 10444
rect 21588 9772 21924 9828
rect 22988 9826 23044 10780
rect 23100 10050 23156 11116
rect 23100 9998 23102 10050
rect 23154 9998 23156 10050
rect 23100 9986 23156 9998
rect 22988 9774 22990 9826
rect 23042 9774 23044 9826
rect 19180 9604 19236 9614
rect 19180 9510 19236 9548
rect 20636 9604 20692 9614
rect 20636 9602 21252 9604
rect 20636 9550 20638 9602
rect 20690 9550 21252 9602
rect 20636 9548 21252 9550
rect 20636 9538 20692 9548
rect 21196 9266 21252 9548
rect 21196 9214 21198 9266
rect 21250 9214 21252 9266
rect 21196 9202 21252 9214
rect 21420 9602 21476 9614
rect 21420 9550 21422 9602
rect 21474 9550 21476 9602
rect 18956 9044 19012 9054
rect 18284 9042 18452 9044
rect 18284 8990 18286 9042
rect 18338 8990 18452 9042
rect 18284 8988 18452 8990
rect 18284 8978 18340 8988
rect 18396 8428 18452 8988
rect 18956 8950 19012 8988
rect 19180 9044 19236 9054
rect 19180 8428 19236 8988
rect 21420 9044 21476 9550
rect 21532 9268 21588 9772
rect 21532 9202 21588 9212
rect 21644 9604 21700 9614
rect 21420 8978 21476 8988
rect 17500 8194 17556 8204
rect 17612 8372 18452 8428
rect 17500 7476 17556 7486
rect 17500 7362 17556 7420
rect 17500 7310 17502 7362
rect 17554 7310 17556 7362
rect 17500 7028 17556 7310
rect 17164 5170 17220 5180
rect 17276 6972 17556 7028
rect 14700 5070 14702 5122
rect 14754 5070 14756 5122
rect 14700 4340 14756 5070
rect 14588 4284 14700 4340
rect 14588 3666 14644 4284
rect 14700 4274 14756 4284
rect 15148 5122 15204 5134
rect 15148 5070 15150 5122
rect 15202 5070 15204 5122
rect 15148 4228 15204 5070
rect 17276 5124 17332 6972
rect 17500 6578 17556 6590
rect 17500 6526 17502 6578
rect 17554 6526 17556 6578
rect 17500 6468 17556 6526
rect 17500 6402 17556 6412
rect 17276 5058 17332 5068
rect 17388 6020 17444 6030
rect 16604 5012 16660 5022
rect 15484 4900 15540 4910
rect 15484 4562 15540 4844
rect 15484 4510 15486 4562
rect 15538 4510 15540 4562
rect 15484 4498 15540 4510
rect 16268 4452 16324 4462
rect 16268 4358 16324 4396
rect 16604 4338 16660 4956
rect 17164 5012 17220 5022
rect 16836 4732 17100 4742
rect 16892 4676 16940 4732
rect 16996 4676 17044 4732
rect 16836 4666 17100 4676
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 16828 4450 16884 4462
rect 16828 4398 16830 4450
rect 16882 4398 16884 4450
rect 15148 4162 15204 4172
rect 14588 3614 14590 3666
rect 14642 3614 14644 3666
rect 14588 3602 14644 3614
rect 14812 4116 14868 4126
rect 14812 3666 14868 4060
rect 14812 3614 14814 3666
rect 14866 3614 14868 3666
rect 14812 3602 14868 3614
rect 16828 3556 16884 4398
rect 17164 3666 17220 4956
rect 17388 5010 17444 5964
rect 17500 5908 17556 5918
rect 17612 5908 17668 8372
rect 18396 8260 18452 8372
rect 18396 8194 18452 8204
rect 18732 8372 19236 8428
rect 19292 8820 19348 8830
rect 18732 8034 18788 8372
rect 19292 8370 19348 8764
rect 20742 8652 21006 8662
rect 20798 8596 20846 8652
rect 20902 8596 20950 8652
rect 20742 8586 21006 8596
rect 19292 8318 19294 8370
rect 19346 8318 19348 8370
rect 19292 8306 19348 8318
rect 19516 8258 19572 8270
rect 19516 8206 19518 8258
rect 19570 8206 19572 8258
rect 18732 7982 18734 8034
rect 18786 7982 18788 8034
rect 18732 7970 18788 7982
rect 19404 8148 19460 8158
rect 17948 7700 18004 7710
rect 17836 6804 17892 6814
rect 17500 5906 17668 5908
rect 17500 5854 17502 5906
rect 17554 5854 17668 5906
rect 17500 5852 17668 5854
rect 17724 6748 17836 6804
rect 17724 5908 17780 6748
rect 17836 6738 17892 6748
rect 17836 6466 17892 6478
rect 17836 6414 17838 6466
rect 17890 6414 17892 6466
rect 17836 6356 17892 6414
rect 17836 6290 17892 6300
rect 17836 5908 17892 5918
rect 17724 5906 17892 5908
rect 17724 5854 17838 5906
rect 17890 5854 17892 5906
rect 17724 5852 17892 5854
rect 17500 5842 17556 5852
rect 17836 5842 17892 5852
rect 17388 4958 17390 5010
rect 17442 4958 17444 5010
rect 17388 4946 17444 4958
rect 17724 5124 17780 5134
rect 17724 4562 17780 5068
rect 17724 4510 17726 4562
rect 17778 4510 17780 4562
rect 17724 4498 17780 4510
rect 17948 4564 18004 7644
rect 19404 7586 19460 8092
rect 19404 7534 19406 7586
rect 19458 7534 19460 7586
rect 19404 7522 19460 7534
rect 18732 7476 18788 7486
rect 18396 7364 18452 7374
rect 18396 7270 18452 7308
rect 18172 6580 18228 6590
rect 18060 5796 18116 5806
rect 18060 5124 18116 5740
rect 18172 5346 18228 6524
rect 18284 6468 18340 6478
rect 18284 6374 18340 6412
rect 18172 5294 18174 5346
rect 18226 5294 18228 5346
rect 18172 5282 18228 5294
rect 18620 6356 18676 6366
rect 18060 5068 18228 5124
rect 18060 4564 18116 4574
rect 17948 4562 18116 4564
rect 17948 4510 18062 4562
rect 18114 4510 18116 4562
rect 17948 4508 18116 4510
rect 18060 4498 18116 4508
rect 17164 3614 17166 3666
rect 17218 3614 17220 3666
rect 17164 3602 17220 3614
rect 17724 3668 17780 3678
rect 17724 3574 17780 3612
rect 18172 3666 18228 5068
rect 18508 5122 18564 5134
rect 18508 5070 18510 5122
rect 18562 5070 18564 5122
rect 18508 4340 18564 5070
rect 18396 4228 18452 4238
rect 18396 4134 18452 4172
rect 18172 3614 18174 3666
rect 18226 3614 18228 3666
rect 18172 3602 18228 3614
rect 18396 3668 18452 3678
rect 18508 3668 18564 4284
rect 18620 3780 18676 6300
rect 18732 5010 18788 7420
rect 19180 6804 19236 6814
rect 19180 6710 19236 6748
rect 18844 6692 18900 6702
rect 18844 6598 18900 6636
rect 19516 6692 19572 8206
rect 21196 8260 21252 8270
rect 21196 8166 21252 8204
rect 19516 6626 19572 6636
rect 19628 8034 19684 8046
rect 19628 7982 19630 8034
rect 19682 7982 19684 8034
rect 18732 4958 18734 5010
rect 18786 4958 18788 5010
rect 18732 4946 18788 4958
rect 18620 3714 18676 3724
rect 18956 4564 19012 4574
rect 18452 3612 18564 3668
rect 18396 3602 18452 3612
rect 16828 3490 16884 3500
rect 14252 3378 14308 3388
rect 15820 3444 15876 3454
rect 15820 3350 15876 3388
rect 18956 3442 19012 4508
rect 19404 4452 19460 4462
rect 19404 4358 19460 4396
rect 19628 4004 19684 7982
rect 20524 8036 20580 8046
rect 20076 7252 20132 7262
rect 20076 7158 20132 7196
rect 20300 6692 20356 6702
rect 20188 6580 20244 6590
rect 20188 6486 20244 6524
rect 20188 6020 20244 6030
rect 19740 6018 20244 6020
rect 19740 5966 20190 6018
rect 20242 5966 20244 6018
rect 19740 5964 20244 5966
rect 19740 5346 19796 5964
rect 20188 5954 20244 5964
rect 20300 5572 20356 6636
rect 19740 5294 19742 5346
rect 19794 5294 19796 5346
rect 19740 5282 19796 5294
rect 20188 5516 20356 5572
rect 19852 5124 19908 5134
rect 19852 5030 19908 5068
rect 20188 4338 20244 5516
rect 20300 5348 20356 5358
rect 20300 4562 20356 5292
rect 20412 5236 20468 5246
rect 20412 5122 20468 5180
rect 20412 5070 20414 5122
rect 20466 5070 20468 5122
rect 20412 5058 20468 5070
rect 20300 4510 20302 4562
rect 20354 4510 20356 4562
rect 20300 4498 20356 4510
rect 20188 4286 20190 4338
rect 20242 4286 20244 4338
rect 20188 4228 20244 4286
rect 20188 4162 20244 4172
rect 20300 4340 20356 4350
rect 19628 3938 19684 3948
rect 19852 3556 19908 3566
rect 19852 3462 19908 3500
rect 18956 3390 18958 3442
rect 19010 3390 19012 3442
rect 18956 3378 19012 3390
rect 20188 3444 20244 3454
rect 20300 3444 20356 4284
rect 20524 3780 20580 7980
rect 20748 8034 20804 8046
rect 20748 7982 20750 8034
rect 20802 7982 20804 8034
rect 20748 7700 20804 7982
rect 20748 7634 20804 7644
rect 20860 7586 20916 7598
rect 20860 7534 20862 7586
rect 20914 7534 20916 7586
rect 20860 7252 20916 7534
rect 20860 7196 21140 7252
rect 20742 7084 21006 7094
rect 20798 7028 20846 7084
rect 20902 7028 20950 7084
rect 20742 7018 21006 7028
rect 20972 6020 21028 6030
rect 20972 5926 21028 5964
rect 20742 5516 21006 5526
rect 20798 5460 20846 5516
rect 20902 5460 20950 5516
rect 20742 5450 21006 5460
rect 21084 5348 21140 7196
rect 21532 6690 21588 6702
rect 21532 6638 21534 6690
rect 21586 6638 21588 6690
rect 21532 6580 21588 6638
rect 21532 6514 21588 6524
rect 21644 5906 21700 9548
rect 22316 9268 22372 9278
rect 22876 9268 22932 9278
rect 22372 9212 22596 9268
rect 22316 9174 22372 9212
rect 21980 8818 22036 8830
rect 21980 8766 21982 8818
rect 22034 8766 22036 8818
rect 21868 8258 21924 8270
rect 21868 8206 21870 8258
rect 21922 8206 21924 8258
rect 21868 6804 21924 8206
rect 21980 7364 22036 8766
rect 21980 7298 22036 7308
rect 21980 6804 22036 6814
rect 21868 6748 21980 6804
rect 21980 6738 22036 6748
rect 22316 6580 22372 6590
rect 21644 5854 21646 5906
rect 21698 5854 21700 5906
rect 21644 5842 21700 5854
rect 21756 6466 21812 6478
rect 21756 6414 21758 6466
rect 21810 6414 21812 6466
rect 21308 5684 21364 5694
rect 21196 5348 21252 5358
rect 21084 5292 21196 5348
rect 21196 5282 21252 5292
rect 20748 4900 20804 4910
rect 20748 4806 20804 4844
rect 21308 4564 21364 5628
rect 21756 5460 21812 6414
rect 22316 6468 22372 6524
rect 22316 6466 22484 6468
rect 22316 6414 22318 6466
rect 22370 6414 22484 6466
rect 22316 6412 22484 6414
rect 22316 6402 22372 6412
rect 21868 6020 21924 6030
rect 22316 6020 22372 6030
rect 21868 6018 22260 6020
rect 21868 5966 21870 6018
rect 21922 5966 22260 6018
rect 21868 5964 22260 5966
rect 21868 5954 21924 5964
rect 21756 5394 21812 5404
rect 21980 5348 22036 5358
rect 21980 5254 22036 5292
rect 22092 5124 22148 5134
rect 22092 5030 22148 5068
rect 21420 4900 21476 4910
rect 21420 4898 21588 4900
rect 21420 4846 21422 4898
rect 21474 4846 21588 4898
rect 21420 4844 21588 4846
rect 21420 4834 21476 4844
rect 21420 4564 21476 4574
rect 21308 4562 21476 4564
rect 21308 4510 21422 4562
rect 21474 4510 21476 4562
rect 21308 4508 21476 4510
rect 21420 4498 21476 4508
rect 21308 4340 21364 4350
rect 21532 4340 21588 4844
rect 21308 4338 21588 4340
rect 21308 4286 21310 4338
rect 21362 4286 21588 4338
rect 21308 4284 21588 4286
rect 21308 4228 21364 4284
rect 21084 4172 21308 4228
rect 22204 4228 22260 5964
rect 22316 5926 22372 5964
rect 22428 5684 22484 6412
rect 22428 5618 22484 5628
rect 22540 5124 22596 9212
rect 22876 9174 22932 9212
rect 22988 8708 23044 9774
rect 23660 9826 23716 12798
rect 24648 12572 24912 12582
rect 24704 12516 24752 12572
rect 24808 12516 24856 12572
rect 24648 12506 24912 12516
rect 25900 12402 25956 13470
rect 26460 13188 26516 13694
rect 26460 12962 26516 13132
rect 26460 12910 26462 12962
rect 26514 12910 26516 12962
rect 26460 12898 26516 12910
rect 27804 13412 27860 13422
rect 27804 12962 27860 13356
rect 27804 12910 27806 12962
rect 27858 12910 27860 12962
rect 25900 12350 25902 12402
rect 25954 12350 25956 12402
rect 25900 12338 25956 12350
rect 23884 12292 23940 12302
rect 23884 12198 23940 12236
rect 27804 12180 27860 12910
rect 27804 12114 27860 12124
rect 27916 12738 27972 12750
rect 27916 12686 27918 12738
rect 27970 12686 27972 12738
rect 25116 11954 25172 11966
rect 25116 11902 25118 11954
rect 25170 11902 25172 11954
rect 25116 11284 25172 11902
rect 25228 11508 25284 11518
rect 25228 11394 25284 11452
rect 26348 11508 26404 11518
rect 25228 11342 25230 11394
rect 25282 11342 25284 11394
rect 25228 11330 25284 11342
rect 25676 11394 25732 11406
rect 25676 11342 25678 11394
rect 25730 11342 25732 11394
rect 25116 11218 25172 11228
rect 24108 11172 24164 11182
rect 24108 11078 24164 11116
rect 24892 11172 24948 11182
rect 24892 11170 25060 11172
rect 24892 11118 24894 11170
rect 24946 11118 25060 11170
rect 24892 11116 25060 11118
rect 24892 11106 24948 11116
rect 24648 11004 24912 11014
rect 24704 10948 24752 11004
rect 24808 10948 24856 11004
rect 24648 10938 24912 10948
rect 23884 10724 23940 10734
rect 23884 10630 23940 10668
rect 24444 10612 24500 10622
rect 23660 9774 23662 9826
rect 23714 9774 23716 9826
rect 23212 8932 23268 8942
rect 23212 8838 23268 8876
rect 22988 8642 23044 8652
rect 23660 8428 23716 9774
rect 23548 8372 23716 8428
rect 23996 9826 24052 9838
rect 23996 9774 23998 9826
rect 24050 9774 24052 9826
rect 23548 8260 23604 8372
rect 23212 7474 23268 7486
rect 23212 7422 23214 7474
rect 23266 7422 23268 7474
rect 23100 6804 23156 6814
rect 23100 6710 23156 6748
rect 23212 5796 23268 7422
rect 23548 7474 23604 8204
rect 23548 7422 23550 7474
rect 23602 7422 23604 7474
rect 23548 7410 23604 7422
rect 23996 6804 24052 9774
rect 24220 9156 24276 9166
rect 24220 9062 24276 9100
rect 24332 8820 24388 8830
rect 24332 8034 24388 8764
rect 24332 7982 24334 8034
rect 24386 7982 24388 8034
rect 24332 7970 24388 7982
rect 24444 7700 24500 10556
rect 25004 9716 25060 11116
rect 25004 9650 25060 9660
rect 25564 10722 25620 10734
rect 25564 10670 25566 10722
rect 25618 10670 25620 10722
rect 25564 9604 25620 10670
rect 25676 9940 25732 11342
rect 25676 9874 25732 9884
rect 25900 10610 25956 10622
rect 25900 10558 25902 10610
rect 25954 10558 25956 10610
rect 25564 9538 25620 9548
rect 25788 9604 25844 9614
rect 24648 9436 24912 9446
rect 24704 9380 24752 9436
rect 24808 9380 24856 9436
rect 24648 9370 24912 9380
rect 25228 9268 25284 9278
rect 25228 9042 25284 9212
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 25228 8978 25284 8990
rect 25340 8820 25396 8830
rect 25340 8726 25396 8764
rect 24892 8260 24948 8270
rect 24892 8258 25172 8260
rect 24892 8206 24894 8258
rect 24946 8206 25172 8258
rect 24892 8204 25172 8206
rect 24892 8194 24948 8204
rect 25004 8034 25060 8046
rect 25004 7982 25006 8034
rect 25058 7982 25060 8034
rect 24648 7868 24912 7878
rect 24704 7812 24752 7868
rect 24808 7812 24856 7868
rect 24648 7802 24912 7812
rect 24668 7700 24724 7710
rect 24444 7698 24724 7700
rect 24444 7646 24670 7698
rect 24722 7646 24724 7698
rect 24444 7644 24724 7646
rect 24668 7634 24724 7644
rect 24332 7476 24388 7486
rect 24332 7382 24388 7420
rect 23996 6738 24052 6748
rect 24108 7364 24164 7374
rect 24108 6578 24164 7308
rect 24108 6526 24110 6578
rect 24162 6526 24164 6578
rect 24108 6514 24164 6526
rect 24648 6300 24912 6310
rect 24704 6244 24752 6300
rect 24808 6244 24856 6300
rect 24648 6234 24912 6244
rect 25004 6020 25060 7982
rect 25116 6580 25172 8204
rect 25788 8146 25844 9548
rect 25788 8094 25790 8146
rect 25842 8094 25844 8146
rect 25788 8082 25844 8094
rect 25900 8036 25956 10558
rect 26348 10610 26404 11452
rect 27916 11282 27972 12686
rect 27916 11230 27918 11282
rect 27970 11230 27972 11282
rect 27916 11218 27972 11230
rect 28252 12178 28308 12190
rect 28252 12126 28254 12178
rect 28306 12126 28308 12178
rect 26348 10558 26350 10610
rect 26402 10558 26404 10610
rect 26348 10546 26404 10558
rect 26796 11060 26852 11070
rect 26796 10610 26852 11004
rect 28252 10836 28308 12126
rect 28252 10770 28308 10780
rect 26796 10558 26798 10610
rect 26850 10558 26852 10610
rect 26796 10546 26852 10558
rect 28364 10052 28420 17502
rect 28588 17444 28644 17614
rect 28588 17378 28644 17388
rect 29148 17108 29204 18396
rect 29260 17668 29316 18958
rect 29260 17574 29316 17612
rect 29596 17444 29652 17454
rect 29708 17444 29764 17454
rect 29652 17442 29764 17444
rect 29652 17390 29710 17442
rect 29762 17390 29764 17442
rect 29652 17388 29764 17390
rect 29148 17106 29316 17108
rect 29148 17054 29150 17106
rect 29202 17054 29316 17106
rect 29148 17052 29316 17054
rect 29148 17042 29204 17052
rect 29260 16884 29316 17052
rect 28812 16660 28868 16670
rect 28812 16658 28980 16660
rect 28812 16606 28814 16658
rect 28866 16606 28980 16658
rect 28812 16604 28980 16606
rect 28812 16594 28868 16604
rect 28554 16492 28818 16502
rect 28610 16436 28658 16492
rect 28714 16436 28762 16492
rect 28554 16426 28818 16436
rect 28924 16436 28980 16604
rect 28924 16370 28980 16380
rect 29148 16212 29204 16222
rect 29260 16212 29316 16828
rect 29372 16436 29428 16446
rect 29428 16380 29540 16436
rect 29372 16370 29428 16380
rect 28700 16210 29316 16212
rect 28700 16158 29150 16210
rect 29202 16158 29262 16210
rect 29314 16158 29316 16210
rect 28700 16156 29316 16158
rect 28700 16098 28756 16156
rect 29148 16146 29204 16156
rect 29260 16146 29316 16156
rect 28700 16046 28702 16098
rect 28754 16046 28756 16098
rect 28700 16034 28756 16046
rect 29372 15314 29428 15326
rect 29372 15262 29374 15314
rect 29426 15262 29428 15314
rect 28554 14924 28818 14934
rect 28610 14868 28658 14924
rect 28714 14868 28762 14924
rect 28554 14858 28818 14868
rect 29372 14196 29428 15262
rect 29372 14130 29428 14140
rect 28554 13356 28818 13366
rect 28610 13300 28658 13356
rect 28714 13300 28762 13356
rect 28554 13290 28818 13300
rect 29484 12850 29540 16380
rect 29596 14308 29652 17388
rect 29708 17378 29764 17388
rect 29820 16322 29876 16334
rect 29820 16270 29822 16322
rect 29874 16270 29876 16322
rect 29820 16210 29876 16270
rect 29820 16158 29822 16210
rect 29874 16158 29876 16210
rect 29820 15314 29876 16158
rect 29820 15262 29822 15314
rect 29874 15262 29876 15314
rect 29820 15148 29876 15262
rect 29596 14242 29652 14252
rect 29708 15092 29876 15148
rect 29484 12798 29486 12850
rect 29538 12798 29540 12850
rect 29484 12786 29540 12798
rect 29708 13858 29764 15092
rect 29708 13806 29710 13858
rect 29762 13806 29764 13858
rect 29596 12404 29652 12414
rect 29708 12404 29764 13806
rect 28812 12402 29764 12404
rect 28812 12350 29598 12402
rect 29650 12350 29764 12402
rect 28812 12348 29764 12350
rect 29820 14308 29876 14318
rect 28812 12178 28868 12348
rect 28812 12126 28814 12178
rect 28866 12126 28868 12178
rect 28812 12114 28868 12126
rect 29148 12180 29204 12190
rect 29148 12086 29204 12124
rect 28554 11788 28818 11798
rect 28610 11732 28658 11788
rect 28714 11732 28762 11788
rect 28554 11722 28818 11732
rect 29260 11508 29316 12348
rect 29596 12338 29652 12348
rect 29820 12180 29876 14252
rect 29820 12114 29876 12124
rect 29820 11508 29876 11518
rect 29260 11414 29316 11452
rect 29708 11452 29820 11508
rect 28700 11172 28756 11182
rect 28700 11170 29428 11172
rect 28700 11118 28702 11170
rect 28754 11118 29428 11170
rect 28700 11116 29428 11118
rect 28700 11106 28756 11116
rect 29036 10722 29092 10734
rect 29036 10670 29038 10722
rect 29090 10670 29092 10722
rect 28554 10220 28818 10230
rect 28610 10164 28658 10220
rect 28714 10164 28762 10220
rect 28554 10154 28818 10164
rect 28364 9986 28420 9996
rect 27356 9826 27412 9838
rect 27356 9774 27358 9826
rect 27410 9774 27412 9826
rect 26460 9602 26516 9614
rect 26460 9550 26462 9602
rect 26514 9550 26516 9602
rect 26460 9266 26516 9550
rect 26460 9214 26462 9266
rect 26514 9214 26516 9266
rect 26460 9202 26516 9214
rect 27132 9602 27188 9614
rect 27132 9550 27134 9602
rect 27186 9550 27188 9602
rect 26348 9042 26404 9054
rect 26348 8990 26350 9042
rect 26402 8990 26404 9042
rect 26348 8708 26404 8990
rect 26348 8642 26404 8652
rect 27132 8148 27188 9550
rect 27356 9492 27412 9774
rect 27468 9604 27524 9614
rect 27468 9510 27524 9548
rect 28588 9602 28644 9614
rect 28588 9550 28590 9602
rect 28642 9550 28644 9602
rect 27356 9268 27412 9436
rect 28588 9492 28644 9550
rect 28588 9426 28644 9436
rect 27580 9268 27636 9278
rect 27356 9266 27636 9268
rect 27356 9214 27582 9266
rect 27634 9214 27636 9266
rect 27356 9212 27636 9214
rect 27356 8708 27412 9212
rect 27580 9202 27636 9212
rect 27356 8428 27412 8652
rect 28028 9042 28084 9054
rect 28028 8990 28030 9042
rect 28082 8990 28084 9042
rect 28028 8484 28084 8990
rect 28364 9042 28420 9054
rect 28364 8990 28366 9042
rect 28418 8990 28420 9042
rect 27356 8372 27524 8428
rect 28028 8418 28084 8428
rect 28140 8820 28196 8830
rect 27132 8082 27188 8092
rect 25900 7028 25956 7980
rect 26236 7364 26292 7374
rect 26236 7270 26292 7308
rect 25116 6514 25172 6524
rect 25676 6972 25956 7028
rect 25004 5954 25060 5964
rect 25340 6020 25396 6030
rect 25340 6018 25508 6020
rect 25340 5966 25342 6018
rect 25394 5966 25508 6018
rect 25340 5964 25508 5966
rect 25340 5954 25396 5964
rect 23436 5796 23492 5806
rect 23212 5794 23492 5796
rect 23212 5742 23438 5794
rect 23490 5742 23492 5794
rect 23212 5740 23492 5742
rect 23436 5730 23492 5740
rect 23772 5348 23828 5358
rect 23772 5254 23828 5292
rect 24332 5236 24388 5246
rect 24332 5142 24388 5180
rect 25340 5234 25396 5246
rect 25340 5182 25342 5234
rect 25394 5182 25396 5234
rect 22540 5058 22596 5068
rect 23100 5122 23156 5134
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 22764 4900 22820 4910
rect 22764 4450 22820 4844
rect 23100 4562 23156 5070
rect 24668 5124 24724 5134
rect 24668 5030 24724 5068
rect 25340 4900 25396 5182
rect 25340 4834 25396 4844
rect 24648 4732 24912 4742
rect 24704 4676 24752 4732
rect 24808 4676 24856 4732
rect 24648 4666 24912 4676
rect 23100 4510 23102 4562
rect 23154 4510 23156 4562
rect 23100 4498 23156 4510
rect 22764 4398 22766 4450
rect 22818 4398 22820 4450
rect 22764 4386 22820 4398
rect 23548 4340 23604 4350
rect 23548 4246 23604 4284
rect 25228 4338 25284 4350
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 24108 4228 24164 4238
rect 22204 4172 22820 4228
rect 20742 3948 21006 3958
rect 20798 3892 20846 3948
rect 20902 3892 20950 3948
rect 20742 3882 21006 3892
rect 20860 3780 20916 3790
rect 20524 3778 20916 3780
rect 20524 3726 20862 3778
rect 20914 3726 20916 3778
rect 20524 3724 20916 3726
rect 20860 3714 20916 3724
rect 21084 3554 21140 4172
rect 21308 4162 21364 4172
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 22204 3556 22260 3566
rect 22204 3462 22260 3500
rect 22764 3554 22820 4172
rect 23436 3892 23492 3902
rect 23436 3666 23492 3836
rect 23436 3614 23438 3666
rect 23490 3614 23492 3666
rect 23436 3602 23492 3614
rect 24108 3666 24164 4172
rect 24668 4228 24724 4238
rect 24668 4134 24724 4172
rect 24220 4116 24276 4126
rect 24220 4022 24276 4060
rect 24108 3614 24110 3666
rect 24162 3614 24164 3666
rect 24108 3602 24164 3614
rect 25004 3668 25060 3678
rect 22764 3502 22766 3554
rect 22818 3502 22820 3554
rect 22764 3490 22820 3502
rect 24220 3556 24276 3566
rect 20188 3442 20356 3444
rect 20188 3390 20190 3442
rect 20242 3390 20356 3442
rect 20188 3388 20356 3390
rect 22428 3444 22484 3454
rect 20188 3378 20244 3388
rect 22428 3350 22484 3388
rect 12348 3332 12404 3342
rect 12348 3238 12404 3276
rect 22876 3332 22932 3342
rect 16836 3164 17100 3174
rect 16892 3108 16940 3164
rect 16996 3108 17044 3164
rect 16836 3098 17100 3108
rect 12236 2706 12292 2716
rect 22876 800 22932 3276
rect 24220 800 24276 3500
rect 24556 3332 24612 3370
rect 24556 3266 24612 3276
rect 24648 3164 24912 3174
rect 24704 3108 24752 3164
rect 24808 3108 24856 3164
rect 24648 3098 24912 3108
rect 25004 1652 25060 3612
rect 25116 3556 25172 3566
rect 25116 3462 25172 3500
rect 25228 3444 25284 4286
rect 25228 3378 25284 3388
rect 25452 3444 25508 5964
rect 25564 4450 25620 4462
rect 25564 4398 25566 4450
rect 25618 4398 25620 4450
rect 25564 3554 25620 4398
rect 25564 3502 25566 3554
rect 25618 3502 25620 3554
rect 25564 3490 25620 3502
rect 25452 3378 25508 3388
rect 25676 3332 25732 6972
rect 25900 6804 25956 6814
rect 25900 6710 25956 6748
rect 27468 6692 27524 8372
rect 28140 8258 28196 8764
rect 28140 8206 28142 8258
rect 28194 8206 28196 8258
rect 28140 8194 28196 8206
rect 28364 7812 28420 8990
rect 28554 8652 28818 8662
rect 28610 8596 28658 8652
rect 28714 8596 28762 8652
rect 28554 8586 28818 8596
rect 28700 8484 28756 8494
rect 28700 8260 28756 8428
rect 28364 7746 28420 7756
rect 28476 8258 28756 8260
rect 28476 8206 28702 8258
rect 28754 8206 28756 8258
rect 28476 8204 28756 8206
rect 27580 7588 27636 7598
rect 27580 7586 28420 7588
rect 27580 7534 27582 7586
rect 27634 7534 28420 7586
rect 27580 7532 28420 7534
rect 27580 7522 27636 7532
rect 28252 6692 28308 6702
rect 27468 6690 28308 6692
rect 27468 6638 28254 6690
rect 28306 6638 28308 6690
rect 27468 6636 28308 6638
rect 26908 6580 26964 6590
rect 26908 6486 26964 6524
rect 27356 6132 27412 6142
rect 25788 6020 25844 6030
rect 25788 5926 25844 5964
rect 27132 5794 27188 5806
rect 27132 5742 27134 5794
rect 27186 5742 27188 5794
rect 26236 5460 26292 5470
rect 26124 5012 26180 5022
rect 25788 4900 25844 4910
rect 25788 4898 26068 4900
rect 25788 4846 25790 4898
rect 25842 4846 26068 4898
rect 25788 4844 26068 4846
rect 25788 4834 25844 4844
rect 26012 4562 26068 4844
rect 26012 4510 26014 4562
rect 26066 4510 26068 4562
rect 26012 4498 26068 4510
rect 26012 3668 26068 3678
rect 26012 3574 26068 3612
rect 24892 1596 25060 1652
rect 25564 3276 25732 3332
rect 24892 800 24948 1596
rect 25564 800 25620 3276
rect 26124 2548 26180 4956
rect 26236 4338 26292 5404
rect 26572 5012 26628 5022
rect 26572 4918 26628 4956
rect 27132 4788 27188 5742
rect 27132 4722 27188 4732
rect 26796 4564 26852 4574
rect 26796 4470 26852 4508
rect 26236 4286 26238 4338
rect 26290 4286 26292 4338
rect 26236 4274 26292 4286
rect 27356 4226 27412 6076
rect 27356 4174 27358 4226
rect 27410 4174 27412 4226
rect 27356 4162 27412 4174
rect 27468 6132 27524 6636
rect 28252 6626 28308 6636
rect 27580 6132 27636 6142
rect 27468 6130 27636 6132
rect 27468 6078 27582 6130
rect 27634 6078 27636 6130
rect 27468 6076 27636 6078
rect 27468 4564 27524 6076
rect 27580 6066 27636 6076
rect 28364 6130 28420 7532
rect 28476 7474 28532 8204
rect 28700 8194 28756 8204
rect 28476 7422 28478 7474
rect 28530 7422 28532 7474
rect 28476 7410 28532 7422
rect 28924 7474 28980 7486
rect 28924 7422 28926 7474
rect 28978 7422 28980 7474
rect 28554 7084 28818 7094
rect 28610 7028 28658 7084
rect 28714 7028 28762 7084
rect 28554 7018 28818 7028
rect 28476 6916 28532 6926
rect 28476 6578 28532 6860
rect 28476 6526 28478 6578
rect 28530 6526 28532 6578
rect 28476 6514 28532 6526
rect 28364 6078 28366 6130
rect 28418 6078 28420 6130
rect 28364 6066 28420 6078
rect 28554 5516 28818 5526
rect 28610 5460 28658 5516
rect 28714 5460 28762 5516
rect 28554 5450 28818 5460
rect 27580 5236 27636 5246
rect 27580 5142 27636 5180
rect 28140 5012 28196 5022
rect 27468 3554 27524 4508
rect 27692 4564 27748 4574
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 27468 3490 27524 3502
rect 27580 4116 27636 4126
rect 26908 3444 26964 3454
rect 26124 2492 26292 2548
rect 26236 800 26292 2492
rect 26908 800 26964 3388
rect 27580 800 27636 4060
rect 27692 3778 27748 4508
rect 28140 4562 28196 4956
rect 28140 4510 28142 4562
rect 28194 4510 28196 4562
rect 28140 4498 28196 4510
rect 28700 4564 28756 4574
rect 28700 4470 28756 4508
rect 27916 4340 27972 4350
rect 27916 4338 28420 4340
rect 27916 4286 27918 4338
rect 27970 4286 28420 4338
rect 27916 4284 28420 4286
rect 27916 4274 27972 4284
rect 27692 3726 27694 3778
rect 27746 3726 27748 3778
rect 27692 3714 27748 3726
rect 28252 3892 28308 3902
rect 28252 800 28308 3836
rect 28364 3442 28420 4284
rect 28554 3948 28818 3958
rect 28610 3892 28658 3948
rect 28714 3892 28762 3948
rect 28554 3882 28818 3892
rect 28588 3780 28644 3790
rect 28588 3554 28644 3724
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 28812 3780 28868 3790
rect 28364 3390 28366 3442
rect 28418 3390 28420 3442
rect 28364 3378 28420 3390
rect 28812 2100 28868 3724
rect 28924 3444 28980 7422
rect 29036 6916 29092 10670
rect 29036 6850 29092 6860
rect 29148 10052 29204 10062
rect 29148 6130 29204 9996
rect 29260 8036 29316 8046
rect 29260 7942 29316 7980
rect 29372 6692 29428 11116
rect 29708 9940 29764 11452
rect 29820 11442 29876 11452
rect 29932 10724 29988 20972
rect 30044 16996 30100 21196
rect 30604 20914 30660 20926
rect 30604 20862 30606 20914
rect 30658 20862 30660 20914
rect 30268 20692 30324 20702
rect 30156 19348 30212 19358
rect 30156 19254 30212 19292
rect 30156 17780 30212 17790
rect 30156 17686 30212 17724
rect 30044 16940 30212 16996
rect 30044 16772 30100 16782
rect 30044 16678 30100 16716
rect 30156 16660 30212 16940
rect 30156 16594 30212 16604
rect 30268 16436 30324 20636
rect 30492 19906 30548 19918
rect 30492 19854 30494 19906
rect 30546 19854 30548 19906
rect 30492 17892 30548 19854
rect 30604 18450 30660 20862
rect 30940 19124 30996 29260
rect 31164 28530 31220 28542
rect 31164 28478 31166 28530
rect 31218 28478 31220 28530
rect 31164 26964 31220 28478
rect 31276 27076 31332 30046
rect 31724 29202 31780 29214
rect 31724 29150 31726 29202
rect 31778 29150 31780 29202
rect 31500 28084 31556 28094
rect 31500 27990 31556 28028
rect 31276 27010 31332 27020
rect 31724 27076 31780 29150
rect 31948 28532 32004 28542
rect 31948 28438 32004 28476
rect 31724 27010 31780 27020
rect 31164 26898 31220 26908
rect 31948 26962 32004 26974
rect 31948 26910 31950 26962
rect 32002 26910 32004 26962
rect 31276 26516 31332 26526
rect 31276 26514 31444 26516
rect 31276 26462 31278 26514
rect 31330 26462 31444 26514
rect 31276 26460 31444 26462
rect 31276 26450 31332 26460
rect 31164 22258 31220 22270
rect 31164 22206 31166 22258
rect 31218 22206 31220 22258
rect 31164 21924 31220 22206
rect 31164 21858 31220 21868
rect 31052 21698 31108 21710
rect 31052 21646 31054 21698
rect 31106 21646 31108 21698
rect 31052 20580 31108 21646
rect 31052 20514 31108 20524
rect 30940 19058 30996 19068
rect 31164 19122 31220 19134
rect 31164 19070 31166 19122
rect 31218 19070 31220 19122
rect 30604 18398 30606 18450
rect 30658 18398 30660 18450
rect 30604 18386 30660 18398
rect 31164 18228 31220 19070
rect 31276 18452 31332 18462
rect 31388 18452 31444 26460
rect 31836 26068 31892 26078
rect 31612 26066 31892 26068
rect 31612 26014 31838 26066
rect 31890 26014 31892 26066
rect 31612 26012 31892 26014
rect 31500 25394 31556 25406
rect 31500 25342 31502 25394
rect 31554 25342 31556 25394
rect 31500 24948 31556 25342
rect 31500 24882 31556 24892
rect 31500 23828 31556 23838
rect 31612 23828 31668 26012
rect 31836 26002 31892 26012
rect 31500 23826 31668 23828
rect 31500 23774 31502 23826
rect 31554 23774 31668 23826
rect 31500 23772 31668 23774
rect 31724 24946 31780 24958
rect 31724 24894 31726 24946
rect 31778 24894 31780 24946
rect 31500 23762 31556 23772
rect 31500 23042 31556 23054
rect 31500 22990 31502 23042
rect 31554 22990 31556 23042
rect 31500 22932 31556 22990
rect 31500 22866 31556 22876
rect 31500 21476 31556 21486
rect 31500 20914 31556 21420
rect 31500 20862 31502 20914
rect 31554 20862 31556 20914
rect 31500 20850 31556 20862
rect 31500 20130 31556 20142
rect 31500 20078 31502 20130
rect 31554 20078 31556 20130
rect 31500 19460 31556 20078
rect 31500 19394 31556 19404
rect 31500 18452 31556 18462
rect 31388 18450 31556 18452
rect 31388 18398 31502 18450
rect 31554 18398 31556 18450
rect 31388 18396 31556 18398
rect 31276 18358 31332 18396
rect 31500 18386 31556 18396
rect 31164 18162 31220 18172
rect 30492 17826 30548 17836
rect 31164 17556 31220 17566
rect 31164 17462 31220 17500
rect 29932 10658 29988 10668
rect 30044 16380 30324 16436
rect 31052 16994 31108 17006
rect 31052 16942 31054 16994
rect 31106 16942 31108 16994
rect 29820 10388 29876 10398
rect 29820 10386 29988 10388
rect 29820 10334 29822 10386
rect 29874 10334 29988 10386
rect 29820 10332 29988 10334
rect 29820 10322 29876 10332
rect 29820 9940 29876 9950
rect 29708 9938 29876 9940
rect 29708 9886 29822 9938
rect 29874 9886 29876 9938
rect 29708 9884 29876 9886
rect 29708 8484 29764 9884
rect 29820 9874 29876 9884
rect 29708 8372 29764 8428
rect 29708 8370 29876 8372
rect 29708 8318 29710 8370
rect 29762 8318 29876 8370
rect 29708 8316 29876 8318
rect 29708 8306 29764 8316
rect 29372 6626 29428 6636
rect 29148 6078 29150 6130
rect 29202 6078 29204 6130
rect 29148 6066 29204 6078
rect 29036 5684 29092 5694
rect 29036 3668 29092 5628
rect 29820 5234 29876 8316
rect 29932 5908 29988 10332
rect 30044 10164 30100 16380
rect 30156 16212 30212 16222
rect 30156 16118 30212 16156
rect 31052 15652 31108 16942
rect 31724 16996 31780 24894
rect 31948 21700 32004 26910
rect 32060 23826 32116 30268
rect 32172 29316 32228 29326
rect 32172 29222 32228 29260
rect 32284 28980 32340 31612
rect 32460 29820 32724 29830
rect 32516 29764 32564 29820
rect 32620 29764 32668 29820
rect 32460 29754 32724 29764
rect 32172 28924 32340 28980
rect 32172 26514 32228 28924
rect 32460 28252 32724 28262
rect 32516 28196 32564 28252
rect 32620 28196 32668 28252
rect 32460 28186 32724 28196
rect 32172 26462 32174 26514
rect 32226 26462 32228 26514
rect 32172 26450 32228 26462
rect 32284 27634 32340 27646
rect 32284 27582 32286 27634
rect 32338 27582 32340 27634
rect 32172 25620 32228 25630
rect 32172 25394 32228 25564
rect 32172 25342 32174 25394
rect 32226 25342 32228 25394
rect 32172 25330 32228 25342
rect 32284 25172 32340 27582
rect 32460 26684 32724 26694
rect 32516 26628 32564 26684
rect 32620 26628 32668 26684
rect 32460 26618 32724 26628
rect 32060 23774 32062 23826
rect 32114 23774 32116 23826
rect 32060 23762 32116 23774
rect 32172 25116 32340 25172
rect 32460 25116 32724 25126
rect 32172 23154 32228 25116
rect 32516 25060 32564 25116
rect 32620 25060 32668 25116
rect 32460 25050 32724 25060
rect 32284 24948 32340 24958
rect 32284 24854 32340 24892
rect 32460 23548 32724 23558
rect 32516 23492 32564 23548
rect 32620 23492 32668 23548
rect 32460 23482 32724 23492
rect 32172 23102 32174 23154
rect 32226 23102 32228 23154
rect 32172 23090 32228 23102
rect 32460 21980 32724 21990
rect 32516 21924 32564 21980
rect 32620 21924 32668 21980
rect 32460 21914 32724 21924
rect 31948 21644 32116 21700
rect 31836 21476 31892 21486
rect 31836 18562 31892 21420
rect 31948 21474 32004 21486
rect 31948 21422 31950 21474
rect 32002 21422 32004 21474
rect 31948 20244 32004 21422
rect 31948 20178 32004 20188
rect 32060 19236 32116 21644
rect 32172 21476 32228 21486
rect 32172 21382 32228 21420
rect 32460 20412 32724 20422
rect 32516 20356 32564 20412
rect 32620 20356 32668 20412
rect 32460 20346 32724 20356
rect 31836 18510 31838 18562
rect 31890 18510 31892 18562
rect 31836 18116 31892 18510
rect 31948 19180 32116 19236
rect 31948 18340 32004 19180
rect 32060 19010 32116 19022
rect 32060 18958 32062 19010
rect 32114 18958 32116 19010
rect 32060 18452 32116 18958
rect 32460 18844 32724 18854
rect 32516 18788 32564 18844
rect 32620 18788 32668 18844
rect 32460 18778 32724 18788
rect 32060 18386 32116 18396
rect 31948 18274 32004 18284
rect 31836 18060 32116 18116
rect 32060 17778 32116 18060
rect 32060 17726 32062 17778
rect 32114 17726 32116 17778
rect 32060 17668 32116 17726
rect 31836 16996 31892 17006
rect 31724 16994 31892 16996
rect 31724 16942 31838 16994
rect 31890 16942 31892 16994
rect 31724 16940 31892 16942
rect 31836 16930 31892 16940
rect 32060 16882 32116 17612
rect 32460 17276 32724 17286
rect 32516 17220 32564 17276
rect 32620 17220 32668 17276
rect 32460 17210 32724 17220
rect 32060 16830 32062 16882
rect 32114 16830 32116 16882
rect 32060 16210 32116 16830
rect 32060 16158 32062 16210
rect 32114 16158 32116 16210
rect 32060 16146 32116 16158
rect 31164 15988 31220 15998
rect 31164 15894 31220 15932
rect 32460 15708 32724 15718
rect 32516 15652 32564 15708
rect 32620 15652 32668 15708
rect 32460 15642 32724 15652
rect 31052 15586 31108 15596
rect 30716 15314 30772 15326
rect 30716 15262 30718 15314
rect 30770 15262 30772 15314
rect 30716 15092 30772 15262
rect 31612 15314 31668 15326
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 30156 14644 30212 14654
rect 30156 14550 30212 14588
rect 30716 14308 30772 15036
rect 30716 14242 30772 14252
rect 30828 15202 30884 15214
rect 30828 15150 30830 15202
rect 30882 15150 30884 15202
rect 30380 14196 30436 14206
rect 30156 14084 30212 14094
rect 30156 12068 30212 14028
rect 30380 13074 30436 14140
rect 30380 13022 30382 13074
rect 30434 13022 30436 13074
rect 30380 13010 30436 13022
rect 30268 12068 30324 12078
rect 30156 12066 30324 12068
rect 30156 12014 30270 12066
rect 30322 12014 30324 12066
rect 30156 12012 30324 12014
rect 30268 12002 30324 12012
rect 30156 11506 30212 11518
rect 30156 11454 30158 11506
rect 30210 11454 30212 11506
rect 30156 11060 30212 11454
rect 30156 10994 30212 11004
rect 30268 11172 30324 11182
rect 30044 10098 30100 10108
rect 30156 10836 30212 10846
rect 30044 9940 30100 9950
rect 30044 6804 30100 9884
rect 30156 9938 30212 10780
rect 30268 10834 30324 11116
rect 30268 10782 30270 10834
rect 30322 10782 30324 10834
rect 30268 10770 30324 10782
rect 30604 10724 30660 10734
rect 30604 10630 30660 10668
rect 30156 9886 30158 9938
rect 30210 9886 30212 9938
rect 30156 9874 30212 9886
rect 30828 9266 30884 15150
rect 31500 15092 31556 15102
rect 31052 15090 31556 15092
rect 31052 15038 31502 15090
rect 31554 15038 31556 15090
rect 31052 15036 31556 15038
rect 30940 10612 30996 10622
rect 30940 10518 30996 10556
rect 30828 9214 30830 9266
rect 30882 9214 30884 9266
rect 30828 9202 30884 9214
rect 30156 8820 30212 8830
rect 30156 8428 30212 8764
rect 30156 8372 30324 8428
rect 30268 8370 30324 8372
rect 30268 8318 30270 8370
rect 30322 8318 30324 8370
rect 30268 8306 30324 8318
rect 30156 7812 30212 7822
rect 30156 7028 30212 7756
rect 31052 7700 31108 15036
rect 31500 15026 31556 15036
rect 31612 15092 31668 15262
rect 31612 15026 31668 15036
rect 31500 14418 31556 14430
rect 31500 14366 31502 14418
rect 31554 14366 31556 14418
rect 31276 13636 31332 13646
rect 31276 12290 31332 13580
rect 31276 12238 31278 12290
rect 31330 12238 31332 12290
rect 31276 12226 31332 12238
rect 31164 11284 31220 11294
rect 31164 11190 31220 11228
rect 31164 9716 31220 9726
rect 31164 9622 31220 9660
rect 31500 9266 31556 14366
rect 32060 14308 32116 14318
rect 32060 14214 32116 14252
rect 32460 14140 32724 14150
rect 32516 14084 32564 14140
rect 32620 14084 32668 14140
rect 32460 14074 32724 14084
rect 32460 12572 32724 12582
rect 32516 12516 32564 12572
rect 32620 12516 32668 12572
rect 32460 12506 32724 12516
rect 32060 11508 32116 11518
rect 32060 11414 32116 11452
rect 32460 11004 32724 11014
rect 32516 10948 32564 11004
rect 32620 10948 32668 11004
rect 32460 10938 32724 10948
rect 32284 10724 32340 10734
rect 32284 10630 32340 10668
rect 31724 10388 31780 10398
rect 31724 10386 31892 10388
rect 31724 10334 31726 10386
rect 31778 10334 31892 10386
rect 31724 10332 31892 10334
rect 31724 10322 31780 10332
rect 31500 9214 31502 9266
rect 31554 9214 31556 9266
rect 31500 9202 31556 9214
rect 31724 9828 31780 9838
rect 31724 9266 31780 9772
rect 31724 9214 31726 9266
rect 31778 9214 31780 9266
rect 31724 9202 31780 9214
rect 31164 8148 31220 8158
rect 31164 8054 31220 8092
rect 31164 7700 31220 7710
rect 31052 7698 31220 7700
rect 31052 7646 31166 7698
rect 31218 7646 31220 7698
rect 31052 7644 31220 7646
rect 31164 7634 31220 7644
rect 31836 7476 31892 10332
rect 32172 10052 32228 10062
rect 32172 9940 32228 9996
rect 32060 9938 32228 9940
rect 32060 9886 32174 9938
rect 32226 9886 32228 9938
rect 32060 9884 32228 9886
rect 32060 9154 32116 9884
rect 32172 9874 32228 9884
rect 32460 9436 32724 9446
rect 32516 9380 32564 9436
rect 32620 9380 32668 9436
rect 32460 9370 32724 9380
rect 32060 9102 32062 9154
rect 32114 9102 32116 9154
rect 32060 9090 32116 9102
rect 31836 7410 31892 7420
rect 32060 8034 32116 8046
rect 32060 7982 32062 8034
rect 32114 7982 32116 8034
rect 31948 7252 32004 7262
rect 31500 7250 32004 7252
rect 31500 7198 31950 7250
rect 32002 7198 32004 7250
rect 31500 7196 32004 7198
rect 30156 6972 30324 7028
rect 30156 6804 30212 6814
rect 30044 6802 30212 6804
rect 30044 6750 30158 6802
rect 30210 6750 30212 6802
rect 30044 6748 30212 6750
rect 30156 6738 30212 6748
rect 30268 6580 30324 6972
rect 29932 5842 29988 5852
rect 30156 6524 30324 6580
rect 31164 6692 31220 6702
rect 29820 5182 29822 5234
rect 29874 5182 29876 5234
rect 29820 4340 29876 5182
rect 30156 5234 30212 6524
rect 30156 5182 30158 5234
rect 30210 5182 30212 5234
rect 30156 5170 30212 5182
rect 31052 5908 31108 5918
rect 29820 3668 29876 4284
rect 30044 5124 30100 5134
rect 30044 3892 30100 5068
rect 30044 3836 30324 3892
rect 29932 3668 29988 3678
rect 30156 3668 30212 3678
rect 29820 3666 29988 3668
rect 29820 3614 29934 3666
rect 29986 3614 29988 3666
rect 29820 3612 29988 3614
rect 29036 3602 29092 3612
rect 29932 3602 29988 3612
rect 30044 3666 30212 3668
rect 30044 3614 30158 3666
rect 30210 3614 30212 3666
rect 30044 3612 30212 3614
rect 30044 3444 30100 3612
rect 30156 3602 30212 3612
rect 30268 3444 30324 3836
rect 28924 3388 30100 3444
rect 30156 3388 30324 3444
rect 31052 3444 31108 5852
rect 31164 5010 31220 6636
rect 31500 6578 31556 7196
rect 31948 7186 32004 7196
rect 32060 6804 32116 7982
rect 32460 7868 32724 7878
rect 32516 7812 32564 7868
rect 32620 7812 32668 7868
rect 32460 7802 32724 7812
rect 32060 6748 32340 6804
rect 31500 6526 31502 6578
rect 31554 6526 31556 6578
rect 31500 6514 31556 6526
rect 32060 6468 32116 6478
rect 32060 6466 32228 6468
rect 32060 6414 32062 6466
rect 32114 6414 32228 6466
rect 32060 6412 32228 6414
rect 32060 6402 32116 6412
rect 31388 5906 31444 5918
rect 31388 5854 31390 5906
rect 31442 5854 31444 5906
rect 31388 5236 31444 5854
rect 31388 5170 31444 5180
rect 32060 5906 32116 5918
rect 32060 5854 32062 5906
rect 32114 5854 32116 5906
rect 32060 5234 32116 5854
rect 32060 5182 32062 5234
rect 32114 5182 32116 5234
rect 32060 5124 32116 5182
rect 31164 4958 31166 5010
rect 31218 4958 31220 5010
rect 31164 4946 31220 4958
rect 31836 5068 32116 5124
rect 31164 4788 31220 4798
rect 31164 4338 31220 4732
rect 31164 4286 31166 4338
rect 31218 4286 31220 4338
rect 31164 4274 31220 4286
rect 31612 4340 31668 4350
rect 31836 4340 31892 5068
rect 32172 5012 32228 6412
rect 31668 4284 31892 4340
rect 32060 4956 32228 5012
rect 31612 4246 31668 4284
rect 31164 3444 31220 3454
rect 31052 3442 31220 3444
rect 31052 3390 31166 3442
rect 31218 3390 31220 3442
rect 31052 3388 31220 3390
rect 28812 2034 28868 2044
rect 30156 1428 30212 3388
rect 31164 3378 31220 3388
rect 30156 1362 30212 1372
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32060 756 32116 4956
rect 32172 4450 32228 4462
rect 32172 4398 32174 4450
rect 32226 4398 32228 4450
rect 32172 2772 32228 4398
rect 32284 4116 32340 6748
rect 32460 6300 32724 6310
rect 32516 6244 32564 6300
rect 32620 6244 32668 6300
rect 32460 6234 32724 6244
rect 32460 4732 32724 4742
rect 32516 4676 32564 4732
rect 32620 4676 32668 4732
rect 32460 4666 32724 4676
rect 32284 4050 32340 4060
rect 32460 3164 32724 3174
rect 32516 3108 32564 3164
rect 32620 3108 32668 3164
rect 32460 3098 32724 3108
rect 32172 2706 32228 2716
rect 32060 690 32116 700
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
<< via2 >>
rect 140 28700 196 28756
rect 1820 32844 1876 32900
rect 2156 30940 2212 30996
rect 2044 30268 2100 30324
rect 1932 29372 1988 29428
rect 1372 28812 1428 28868
rect 2268 29484 2324 29540
rect 2156 27970 2212 27972
rect 2156 27918 2158 27970
rect 2158 27918 2210 27970
rect 2210 27918 2212 27970
rect 2156 27916 2212 27918
rect 2044 27132 2100 27188
rect 2268 27020 2324 27076
rect 2604 29260 2660 29316
rect 2156 26012 2212 26068
rect 2380 25676 2436 25732
rect 1932 25618 1988 25620
rect 1932 25566 1934 25618
rect 1934 25566 1986 25618
rect 1986 25566 1988 25618
rect 1932 25564 1988 25566
rect 812 25116 868 25172
rect 2044 25004 2100 25060
rect 1932 24610 1988 24612
rect 1932 24558 1934 24610
rect 1934 24558 1986 24610
rect 1986 24558 1988 24610
rect 1932 24556 1988 24558
rect 140 18172 196 18228
rect 1820 22876 1876 22932
rect 1708 21196 1764 21252
rect 1596 19794 1652 19796
rect 1596 19742 1598 19794
rect 1598 19742 1650 19794
rect 1650 19742 1652 19794
rect 1596 19740 1652 19742
rect 1260 15820 1316 15876
rect 1596 14364 1652 14420
rect 2044 23996 2100 24052
rect 2156 22428 2212 22484
rect 2268 22540 2324 22596
rect 2156 22092 2212 22148
rect 2156 21644 2212 21700
rect 2268 21980 2324 22036
rect 2156 20860 2212 20916
rect 2044 20802 2100 20804
rect 2044 20750 2046 20802
rect 2046 20750 2098 20802
rect 2098 20750 2100 20802
rect 2044 20748 2100 20750
rect 2044 19292 2100 19348
rect 1932 17500 1988 17556
rect 2492 22428 2548 22484
rect 2604 25228 2660 25284
rect 3724 32284 3780 32340
rect 3388 30156 3444 30212
rect 3276 29708 3332 29764
rect 2940 29426 2996 29428
rect 2940 29374 2942 29426
rect 2942 29374 2994 29426
rect 2994 29374 2996 29426
rect 2940 29372 2996 29374
rect 3052 29148 3108 29204
rect 3164 27804 3220 27860
rect 3052 27580 3108 27636
rect 2940 25564 2996 25620
rect 3164 26402 3220 26404
rect 3164 26350 3166 26402
rect 3166 26350 3218 26402
rect 3218 26350 3220 26402
rect 3164 26348 3220 26350
rect 2940 25228 2996 25284
rect 2940 24556 2996 24612
rect 3052 24444 3108 24500
rect 2380 20130 2436 20132
rect 2380 20078 2382 20130
rect 2382 20078 2434 20130
rect 2434 20078 2436 20130
rect 2380 20076 2436 20078
rect 2268 15874 2324 15876
rect 2268 15822 2270 15874
rect 2270 15822 2322 15874
rect 2322 15822 2324 15874
rect 2268 15820 2324 15822
rect 2604 21420 2660 21476
rect 2492 14476 2548 14532
rect 1708 12962 1764 12964
rect 1708 12910 1710 12962
rect 1710 12910 1762 12962
rect 1762 12910 1764 12962
rect 1708 12908 1764 12910
rect 1484 9996 1540 10052
rect 2044 13132 2100 13188
rect 2380 13970 2436 13972
rect 2380 13918 2382 13970
rect 2382 13918 2434 13970
rect 2434 13918 2436 13970
rect 2380 13916 2436 13918
rect 2492 12348 2548 12404
rect 2380 11564 2436 11620
rect 2268 11452 2324 11508
rect 1932 11394 1988 11396
rect 1932 11342 1934 11394
rect 1934 11342 1986 11394
rect 1986 11342 1988 11394
rect 1932 11340 1988 11342
rect 1820 9548 1876 9604
rect 1932 10444 1988 10500
rect 1596 8316 1652 8372
rect 1820 8764 1876 8820
rect 2044 9324 2100 9380
rect 1260 6412 1316 6468
rect 2044 7644 2100 7700
rect 1820 6188 1876 6244
rect 1932 5404 1988 5460
rect 1596 3388 1652 3444
rect 2828 19852 2884 19908
rect 2716 19740 2772 19796
rect 3164 21532 3220 21588
rect 3052 20690 3108 20692
rect 3052 20638 3054 20690
rect 3054 20638 3106 20690
rect 3106 20638 3108 20690
rect 3052 20636 3108 20638
rect 2940 18450 2996 18452
rect 2940 18398 2942 18450
rect 2942 18398 2994 18450
rect 2994 18398 2996 18450
rect 2940 18396 2996 18398
rect 3052 17836 3108 17892
rect 3052 17554 3108 17556
rect 3052 17502 3054 17554
rect 3054 17502 3106 17554
rect 3106 17502 3108 17554
rect 3052 17500 3108 17502
rect 2828 16828 2884 16884
rect 2716 14418 2772 14420
rect 2716 14366 2718 14418
rect 2718 14366 2770 14418
rect 2770 14366 2772 14418
rect 2716 14364 2772 14366
rect 2604 10892 2660 10948
rect 2716 9996 2772 10052
rect 3164 15260 3220 15316
rect 3052 14700 3108 14756
rect 3052 13468 3108 13524
rect 2940 12962 2996 12964
rect 2940 12910 2942 12962
rect 2942 12910 2994 12962
rect 2994 12910 2996 12962
rect 2940 12908 2996 12910
rect 3612 31612 3668 31668
rect 3836 29708 3892 29764
rect 3948 29596 4004 29652
rect 3724 25676 3780 25732
rect 4620 32956 4676 33012
rect 4172 29986 4228 29988
rect 4172 29934 4174 29986
rect 4174 29934 4226 29986
rect 4226 29934 4228 29986
rect 4172 29932 4228 29934
rect 4172 29314 4228 29316
rect 4172 29262 4174 29314
rect 4174 29262 4226 29314
rect 4226 29262 4228 29314
rect 4172 29260 4228 29262
rect 4060 29036 4116 29092
rect 4060 28754 4116 28756
rect 4060 28702 4062 28754
rect 4062 28702 4114 28754
rect 4114 28702 4116 28754
rect 4060 28700 4116 28702
rect 4172 28252 4228 28308
rect 4396 29202 4452 29204
rect 4396 29150 4398 29202
rect 4398 29150 4450 29202
rect 4450 29150 4452 29202
rect 4396 29148 4452 29150
rect 4508 28364 4564 28420
rect 5118 30602 5174 30604
rect 5118 30550 5120 30602
rect 5120 30550 5172 30602
rect 5172 30550 5174 30602
rect 5118 30548 5174 30550
rect 5222 30602 5278 30604
rect 5222 30550 5224 30602
rect 5224 30550 5276 30602
rect 5276 30550 5278 30602
rect 5222 30548 5278 30550
rect 5326 30602 5382 30604
rect 5326 30550 5328 30602
rect 5328 30550 5380 30602
rect 5380 30550 5382 30602
rect 5326 30548 5382 30550
rect 4956 30098 5012 30100
rect 4956 30046 4958 30098
rect 4958 30046 5010 30098
rect 5010 30046 5012 30098
rect 4956 30044 5012 30046
rect 5628 29820 5684 29876
rect 5740 29708 5796 29764
rect 5180 29148 5236 29204
rect 5118 29034 5174 29036
rect 5118 28982 5120 29034
rect 5120 28982 5172 29034
rect 5172 28982 5174 29034
rect 5118 28980 5174 28982
rect 5222 29034 5278 29036
rect 5222 28982 5224 29034
rect 5224 28982 5276 29034
rect 5276 28982 5278 29034
rect 5222 28980 5278 28982
rect 5326 29034 5382 29036
rect 5326 28982 5328 29034
rect 5328 28982 5380 29034
rect 5380 28982 5382 29034
rect 5326 28980 5382 28982
rect 4844 28588 4900 28644
rect 5628 28588 5684 28644
rect 4396 27634 4452 27636
rect 4396 27582 4398 27634
rect 4398 27582 4450 27634
rect 4450 27582 4452 27634
rect 4396 27580 4452 27582
rect 4172 26460 4228 26516
rect 4060 26236 4116 26292
rect 4172 25452 4228 25508
rect 3500 24668 3556 24724
rect 4172 24498 4228 24500
rect 4172 24446 4174 24498
rect 4174 24446 4226 24498
rect 4226 24446 4228 24498
rect 4172 24444 4228 24446
rect 3724 23884 3780 23940
rect 3948 24220 4004 24276
rect 3388 21980 3444 22036
rect 3500 23548 3556 23604
rect 4060 23100 4116 23156
rect 4172 23884 4228 23940
rect 4172 22540 4228 22596
rect 4172 22092 4228 22148
rect 4060 21532 4116 21588
rect 4172 20748 4228 20804
rect 4060 19964 4116 20020
rect 4060 19180 4116 19236
rect 3724 18450 3780 18452
rect 3724 18398 3726 18450
rect 3726 18398 3778 18450
rect 3778 18398 3780 18450
rect 3724 18396 3780 18398
rect 3948 17612 4004 17668
rect 3500 16828 3556 16884
rect 3948 16044 4004 16100
rect 3276 12348 3332 12404
rect 3724 14476 3780 14532
rect 3836 13074 3892 13076
rect 3836 13022 3838 13074
rect 3838 13022 3890 13074
rect 3890 13022 3892 13074
rect 3836 13020 3892 13022
rect 4060 12460 4116 12516
rect 3052 10332 3108 10388
rect 4508 27186 4564 27188
rect 4508 27134 4510 27186
rect 4510 27134 4562 27186
rect 4562 27134 4564 27186
rect 4508 27132 4564 27134
rect 4732 25618 4788 25620
rect 4732 25566 4734 25618
rect 4734 25566 4786 25618
rect 4786 25566 4788 25618
rect 4732 25564 4788 25566
rect 5118 27466 5174 27468
rect 5118 27414 5120 27466
rect 5120 27414 5172 27466
rect 5172 27414 5174 27466
rect 5118 27412 5174 27414
rect 5222 27466 5278 27468
rect 5222 27414 5224 27466
rect 5224 27414 5276 27466
rect 5276 27414 5278 27466
rect 5222 27412 5278 27414
rect 5326 27466 5382 27468
rect 5326 27414 5328 27466
rect 5328 27414 5380 27466
rect 5380 27414 5382 27466
rect 5326 27412 5382 27414
rect 5068 26178 5124 26180
rect 5068 26126 5070 26178
rect 5070 26126 5122 26178
rect 5122 26126 5124 26178
rect 5068 26124 5124 26126
rect 5118 25898 5174 25900
rect 5118 25846 5120 25898
rect 5120 25846 5172 25898
rect 5172 25846 5174 25898
rect 5118 25844 5174 25846
rect 5222 25898 5278 25900
rect 5222 25846 5224 25898
rect 5224 25846 5276 25898
rect 5276 25846 5278 25898
rect 5222 25844 5278 25846
rect 5326 25898 5382 25900
rect 5326 25846 5328 25898
rect 5328 25846 5380 25898
rect 5380 25846 5382 25898
rect 5326 25844 5382 25846
rect 5740 28252 5796 28308
rect 5516 25676 5572 25732
rect 5964 28028 6020 28084
rect 6636 30380 6692 30436
rect 6412 29820 6468 29876
rect 6188 29148 6244 29204
rect 6188 28642 6244 28644
rect 6188 28590 6190 28642
rect 6190 28590 6242 28642
rect 6242 28590 6244 28642
rect 6188 28588 6244 28590
rect 6076 27692 6132 27748
rect 5964 26290 6020 26292
rect 5964 26238 5966 26290
rect 5966 26238 6018 26290
rect 6018 26238 6020 26290
rect 5964 26236 6020 26238
rect 4620 25228 4676 25284
rect 5740 25282 5796 25284
rect 5740 25230 5742 25282
rect 5742 25230 5794 25282
rect 5794 25230 5796 25282
rect 5740 25228 5796 25230
rect 6300 25004 6356 25060
rect 6524 26962 6580 26964
rect 6524 26910 6526 26962
rect 6526 26910 6578 26962
rect 6578 26910 6580 26962
rect 6524 26908 6580 26910
rect 6412 25228 6468 25284
rect 4956 24834 5012 24836
rect 4956 24782 4958 24834
rect 4958 24782 5010 24834
rect 5010 24782 5012 24834
rect 4956 24780 5012 24782
rect 5964 24780 6020 24836
rect 5118 24330 5174 24332
rect 5118 24278 5120 24330
rect 5120 24278 5172 24330
rect 5172 24278 5174 24330
rect 5118 24276 5174 24278
rect 5222 24330 5278 24332
rect 5222 24278 5224 24330
rect 5224 24278 5276 24330
rect 5276 24278 5278 24330
rect 5222 24276 5278 24278
rect 5326 24330 5382 24332
rect 5326 24278 5328 24330
rect 5328 24278 5380 24330
rect 5380 24278 5382 24330
rect 5326 24276 5382 24278
rect 4508 24050 4564 24052
rect 4508 23998 4510 24050
rect 4510 23998 4562 24050
rect 4562 23998 4564 24050
rect 4508 23996 4564 23998
rect 5068 23938 5124 23940
rect 5068 23886 5070 23938
rect 5070 23886 5122 23938
rect 5122 23886 5124 23938
rect 5068 23884 5124 23886
rect 6300 23884 6356 23940
rect 4956 23154 5012 23156
rect 4956 23102 4958 23154
rect 4958 23102 5010 23154
rect 5010 23102 5012 23154
rect 4956 23100 5012 23102
rect 5118 22762 5174 22764
rect 5118 22710 5120 22762
rect 5120 22710 5172 22762
rect 5172 22710 5174 22762
rect 5118 22708 5174 22710
rect 5222 22762 5278 22764
rect 5222 22710 5224 22762
rect 5224 22710 5276 22762
rect 5276 22710 5278 22762
rect 5222 22708 5278 22710
rect 5326 22762 5382 22764
rect 5326 22710 5328 22762
rect 5328 22710 5380 22762
rect 5380 22710 5382 22762
rect 5326 22708 5382 22710
rect 4620 22428 4676 22484
rect 5068 22482 5124 22484
rect 5068 22430 5070 22482
rect 5070 22430 5122 22482
rect 5122 22430 5124 22482
rect 5068 22428 5124 22430
rect 5628 22428 5684 22484
rect 4620 22146 4676 22148
rect 4620 22094 4622 22146
rect 4622 22094 4674 22146
rect 4674 22094 4676 22146
rect 4620 22092 4676 22094
rect 4956 22092 5012 22148
rect 4620 21698 4676 21700
rect 4620 21646 4622 21698
rect 4622 21646 4674 21698
rect 4674 21646 4676 21698
rect 4620 21644 4676 21646
rect 4620 20972 4676 21028
rect 4508 19346 4564 19348
rect 4508 19294 4510 19346
rect 4510 19294 4562 19346
rect 4562 19294 4564 19346
rect 4508 19292 4564 19294
rect 4508 17836 4564 17892
rect 4732 20860 4788 20916
rect 5118 21194 5174 21196
rect 5118 21142 5120 21194
rect 5120 21142 5172 21194
rect 5172 21142 5174 21194
rect 5118 21140 5174 21142
rect 5222 21194 5278 21196
rect 5222 21142 5224 21194
rect 5224 21142 5276 21194
rect 5276 21142 5278 21194
rect 5222 21140 5278 21142
rect 5326 21194 5382 21196
rect 5326 21142 5328 21194
rect 5328 21142 5380 21194
rect 5380 21142 5382 21194
rect 5326 21140 5382 21142
rect 4956 20188 5012 20244
rect 5964 21586 6020 21588
rect 5964 21534 5966 21586
rect 5966 21534 6018 21586
rect 6018 21534 6020 21586
rect 5964 21532 6020 21534
rect 6524 22146 6580 22148
rect 6524 22094 6526 22146
rect 6526 22094 6578 22146
rect 6578 22094 6580 22146
rect 6524 22092 6580 22094
rect 5852 20076 5908 20132
rect 5118 19626 5174 19628
rect 5118 19574 5120 19626
rect 5120 19574 5172 19626
rect 5172 19574 5174 19626
rect 5118 19572 5174 19574
rect 5222 19626 5278 19628
rect 5222 19574 5224 19626
rect 5224 19574 5276 19626
rect 5276 19574 5278 19626
rect 5222 19572 5278 19574
rect 5326 19626 5382 19628
rect 5326 19574 5328 19626
rect 5328 19574 5380 19626
rect 5380 19574 5382 19626
rect 5326 19572 5382 19574
rect 5964 20018 6020 20020
rect 5964 19966 5966 20018
rect 5966 19966 6018 20018
rect 6018 19966 6020 20018
rect 5964 19964 6020 19966
rect 6412 19292 6468 19348
rect 6076 19234 6132 19236
rect 6076 19182 6078 19234
rect 6078 19182 6130 19234
rect 6130 19182 6132 19234
rect 6076 19180 6132 19182
rect 5628 18396 5684 18452
rect 4956 18284 5012 18340
rect 4956 18060 5012 18116
rect 5118 18058 5174 18060
rect 5118 18006 5120 18058
rect 5120 18006 5172 18058
rect 5172 18006 5174 18058
rect 5118 18004 5174 18006
rect 5222 18058 5278 18060
rect 5222 18006 5224 18058
rect 5224 18006 5276 18058
rect 5276 18006 5278 18058
rect 5222 18004 5278 18006
rect 5326 18058 5382 18060
rect 5326 18006 5328 18058
rect 5328 18006 5380 18058
rect 5380 18006 5382 18058
rect 5326 18004 5382 18006
rect 4732 16210 4788 16212
rect 4732 16158 4734 16210
rect 4734 16158 4786 16210
rect 4786 16158 4788 16210
rect 4732 16156 4788 16158
rect 4620 15314 4676 15316
rect 4620 15262 4622 15314
rect 4622 15262 4674 15314
rect 4674 15262 4676 15314
rect 4620 15260 4676 15262
rect 4396 14588 4452 14644
rect 4396 14028 4452 14084
rect 4732 14588 4788 14644
rect 4620 14306 4676 14308
rect 4620 14254 4622 14306
rect 4622 14254 4674 14306
rect 4674 14254 4676 14306
rect 4620 14252 4676 14254
rect 4508 13020 4564 13076
rect 4732 13580 4788 13636
rect 4396 12348 4452 12404
rect 4172 11340 4228 11396
rect 4508 11228 4564 11284
rect 5404 17500 5460 17556
rect 6188 16994 6244 16996
rect 6188 16942 6190 16994
rect 6190 16942 6242 16994
rect 6242 16942 6244 16994
rect 6188 16940 6244 16942
rect 6076 16716 6132 16772
rect 5118 16490 5174 16492
rect 5118 16438 5120 16490
rect 5120 16438 5172 16490
rect 5172 16438 5174 16490
rect 5118 16436 5174 16438
rect 5222 16490 5278 16492
rect 5222 16438 5224 16490
rect 5224 16438 5276 16490
rect 5276 16438 5278 16490
rect 5222 16436 5278 16438
rect 5326 16490 5382 16492
rect 5326 16438 5328 16490
rect 5328 16438 5380 16490
rect 5380 16438 5382 16490
rect 5326 16436 5382 16438
rect 5068 16210 5124 16212
rect 5068 16158 5070 16210
rect 5070 16158 5122 16210
rect 5122 16158 5124 16210
rect 5068 16156 5124 16158
rect 5964 16156 6020 16212
rect 5628 15260 5684 15316
rect 5118 14922 5174 14924
rect 5118 14870 5120 14922
rect 5120 14870 5172 14922
rect 5172 14870 5174 14922
rect 5118 14868 5174 14870
rect 5222 14922 5278 14924
rect 5222 14870 5224 14922
rect 5224 14870 5276 14922
rect 5276 14870 5278 14922
rect 5222 14868 5278 14870
rect 5326 14922 5382 14924
rect 5326 14870 5328 14922
rect 5328 14870 5380 14922
rect 5380 14870 5382 14922
rect 5326 14868 5382 14870
rect 5628 14700 5684 14756
rect 4956 14252 5012 14308
rect 5964 15314 6020 15316
rect 5964 15262 5966 15314
rect 5966 15262 6018 15314
rect 6018 15262 6020 15314
rect 5964 15260 6020 15262
rect 5740 13916 5796 13972
rect 5404 13858 5460 13860
rect 5404 13806 5406 13858
rect 5406 13806 5458 13858
rect 5458 13806 5460 13858
rect 5404 13804 5460 13806
rect 5292 13468 5348 13524
rect 5118 13354 5174 13356
rect 5118 13302 5120 13354
rect 5120 13302 5172 13354
rect 5172 13302 5174 13354
rect 5118 13300 5174 13302
rect 5222 13354 5278 13356
rect 5222 13302 5224 13354
rect 5224 13302 5276 13354
rect 5276 13302 5278 13354
rect 5222 13300 5278 13302
rect 5326 13354 5382 13356
rect 5326 13302 5328 13354
rect 5328 13302 5380 13354
rect 5380 13302 5382 13354
rect 5326 13300 5382 13302
rect 4844 13020 4900 13076
rect 4956 12850 5012 12852
rect 4956 12798 4958 12850
rect 4958 12798 5010 12850
rect 5010 12798 5012 12850
rect 4956 12796 5012 12798
rect 5516 12402 5572 12404
rect 5516 12350 5518 12402
rect 5518 12350 5570 12402
rect 5570 12350 5572 12402
rect 5516 12348 5572 12350
rect 5118 11786 5174 11788
rect 5118 11734 5120 11786
rect 5120 11734 5172 11786
rect 5172 11734 5174 11786
rect 5118 11732 5174 11734
rect 5222 11786 5278 11788
rect 5222 11734 5224 11786
rect 5224 11734 5276 11786
rect 5276 11734 5278 11786
rect 5222 11732 5278 11734
rect 5326 11786 5382 11788
rect 5326 11734 5328 11786
rect 5328 11734 5380 11786
rect 5380 11734 5382 11786
rect 5326 11732 5382 11734
rect 5740 11618 5796 11620
rect 5740 11566 5742 11618
rect 5742 11566 5794 11618
rect 5794 11566 5796 11618
rect 5740 11564 5796 11566
rect 3836 9660 3892 9716
rect 2828 8764 2884 8820
rect 3276 8316 3332 8372
rect 3052 6300 3108 6356
rect 2268 5852 2324 5908
rect 2940 5292 2996 5348
rect 3500 7308 3556 7364
rect 3388 6636 3444 6692
rect 3388 5740 3444 5796
rect 2380 3724 2436 3780
rect 2604 3442 2660 3444
rect 2604 3390 2606 3442
rect 2606 3390 2658 3442
rect 2658 3390 2660 3442
rect 2604 3388 2660 3390
rect 3948 9212 4004 9268
rect 4508 10444 4564 10500
rect 5292 10386 5348 10388
rect 5292 10334 5294 10386
rect 5294 10334 5346 10386
rect 5346 10334 5348 10386
rect 5292 10332 5348 10334
rect 5118 10218 5174 10220
rect 5118 10166 5120 10218
rect 5120 10166 5172 10218
rect 5172 10166 5174 10218
rect 5118 10164 5174 10166
rect 5222 10218 5278 10220
rect 5222 10166 5224 10218
rect 5224 10166 5276 10218
rect 5276 10166 5278 10218
rect 5222 10164 5278 10166
rect 5326 10218 5382 10220
rect 5326 10166 5328 10218
rect 5328 10166 5380 10218
rect 5380 10166 5382 10218
rect 5326 10164 5382 10166
rect 4620 9548 4676 9604
rect 5068 9602 5124 9604
rect 5068 9550 5070 9602
rect 5070 9550 5122 9602
rect 5122 9550 5124 9602
rect 5068 9548 5124 9550
rect 5964 10668 6020 10724
rect 5964 9548 6020 9604
rect 5852 9324 5908 9380
rect 6748 29932 6804 29988
rect 6972 30044 7028 30100
rect 6860 29260 6916 29316
rect 7644 29596 7700 29652
rect 7308 28924 7364 28980
rect 7420 28700 7476 28756
rect 7532 27186 7588 27188
rect 7532 27134 7534 27186
rect 7534 27134 7586 27186
rect 7586 27134 7588 27186
rect 7532 27132 7588 27134
rect 6860 25564 6916 25620
rect 7308 24780 7364 24836
rect 7084 22092 7140 22148
rect 6860 20914 6916 20916
rect 6860 20862 6862 20914
rect 6862 20862 6914 20914
rect 6914 20862 6916 20914
rect 6860 20860 6916 20862
rect 6972 17724 7028 17780
rect 6412 15820 6468 15876
rect 6636 15426 6692 15428
rect 6636 15374 6638 15426
rect 6638 15374 6690 15426
rect 6690 15374 6692 15426
rect 6636 15372 6692 15374
rect 7084 16828 7140 16884
rect 7420 17948 7476 18004
rect 7420 17778 7476 17780
rect 7420 17726 7422 17778
rect 7422 17726 7474 17778
rect 7474 17726 7476 17778
rect 7420 17724 7476 17726
rect 7420 16156 7476 16212
rect 6748 12908 6804 12964
rect 7308 15874 7364 15876
rect 7308 15822 7310 15874
rect 7310 15822 7362 15874
rect 7362 15822 7364 15874
rect 7308 15820 7364 15822
rect 7420 13356 7476 13412
rect 7420 12348 7476 12404
rect 8652 30380 8708 30436
rect 7980 28252 8036 28308
rect 8092 28588 8148 28644
rect 8652 29932 8708 29988
rect 9324 30156 9380 30212
rect 9436 30268 9492 30324
rect 9772 30098 9828 30100
rect 9772 30046 9774 30098
rect 9774 30046 9826 30098
rect 9826 30046 9828 30098
rect 9772 30044 9828 30046
rect 8764 29708 8820 29764
rect 9024 29818 9080 29820
rect 9024 29766 9026 29818
rect 9026 29766 9078 29818
rect 9078 29766 9080 29818
rect 9024 29764 9080 29766
rect 9128 29818 9184 29820
rect 9128 29766 9130 29818
rect 9130 29766 9182 29818
rect 9182 29766 9184 29818
rect 9128 29764 9184 29766
rect 9232 29818 9288 29820
rect 9232 29766 9234 29818
rect 9234 29766 9286 29818
rect 9286 29766 9288 29818
rect 9232 29764 9288 29766
rect 9996 29820 10052 29876
rect 9548 29650 9604 29652
rect 9548 29598 9550 29650
rect 9550 29598 9602 29650
rect 9602 29598 9604 29650
rect 9548 29596 9604 29598
rect 8764 29484 8820 29540
rect 9996 29484 10052 29540
rect 9548 29260 9604 29316
rect 8988 28476 9044 28532
rect 9024 28250 9080 28252
rect 9024 28198 9026 28250
rect 9026 28198 9078 28250
rect 9078 28198 9080 28250
rect 9024 28196 9080 28198
rect 9128 28250 9184 28252
rect 9128 28198 9130 28250
rect 9130 28198 9182 28250
rect 9182 28198 9184 28250
rect 9128 28196 9184 28198
rect 9232 28250 9288 28252
rect 9232 28198 9234 28250
rect 9234 28198 9286 28250
rect 9286 28198 9288 28250
rect 9232 28196 9288 28198
rect 8764 27916 8820 27972
rect 7756 25228 7812 25284
rect 8092 25116 8148 25172
rect 7756 24892 7812 24948
rect 8204 24892 8260 24948
rect 9024 26682 9080 26684
rect 9024 26630 9026 26682
rect 9026 26630 9078 26682
rect 9078 26630 9080 26682
rect 9024 26628 9080 26630
rect 9128 26682 9184 26684
rect 9128 26630 9130 26682
rect 9130 26630 9182 26682
rect 9182 26630 9184 26682
rect 9128 26628 9184 26630
rect 9232 26682 9288 26684
rect 9232 26630 9234 26682
rect 9234 26630 9286 26682
rect 9286 26630 9288 26682
rect 9232 26628 9288 26630
rect 9100 26402 9156 26404
rect 9100 26350 9102 26402
rect 9102 26350 9154 26402
rect 9154 26350 9156 26402
rect 9100 26348 9156 26350
rect 8540 25116 8596 25172
rect 8540 24668 8596 24724
rect 8652 24892 8708 24948
rect 9024 25114 9080 25116
rect 9024 25062 9026 25114
rect 9026 25062 9078 25114
rect 9078 25062 9080 25114
rect 9024 25060 9080 25062
rect 9128 25114 9184 25116
rect 9128 25062 9130 25114
rect 9130 25062 9182 25114
rect 9182 25062 9184 25114
rect 9128 25060 9184 25062
rect 9232 25114 9288 25116
rect 9232 25062 9234 25114
rect 9234 25062 9286 25114
rect 9286 25062 9288 25114
rect 9232 25060 9288 25062
rect 8988 24722 9044 24724
rect 8988 24670 8990 24722
rect 8990 24670 9042 24722
rect 9042 24670 9044 24722
rect 8988 24668 9044 24670
rect 8316 23660 8372 23716
rect 8092 23100 8148 23156
rect 8092 20636 8148 20692
rect 9100 23772 9156 23828
rect 9024 23546 9080 23548
rect 9024 23494 9026 23546
rect 9026 23494 9078 23546
rect 9078 23494 9080 23546
rect 9024 23492 9080 23494
rect 9128 23546 9184 23548
rect 9128 23494 9130 23546
rect 9130 23494 9182 23546
rect 9182 23494 9184 23546
rect 9128 23492 9184 23494
rect 9232 23546 9288 23548
rect 9232 23494 9234 23546
rect 9234 23494 9286 23546
rect 9286 23494 9288 23546
rect 9232 23492 9288 23494
rect 10108 29426 10164 29428
rect 10108 29374 10110 29426
rect 10110 29374 10162 29426
rect 10162 29374 10164 29426
rect 10108 29372 10164 29374
rect 9548 28754 9604 28756
rect 9548 28702 9550 28754
rect 9550 28702 9602 28754
rect 9602 28702 9604 28754
rect 9548 28700 9604 28702
rect 9548 28028 9604 28084
rect 9772 27020 9828 27076
rect 9884 24668 9940 24724
rect 9772 24610 9828 24612
rect 9772 24558 9774 24610
rect 9774 24558 9826 24610
rect 9826 24558 9828 24610
rect 9772 24556 9828 24558
rect 9660 24108 9716 24164
rect 9436 23436 9492 23492
rect 9548 23660 9604 23716
rect 9660 23548 9716 23604
rect 8540 22482 8596 22484
rect 8540 22430 8542 22482
rect 8542 22430 8594 22482
rect 8594 22430 8596 22482
rect 8540 22428 8596 22430
rect 9024 21978 9080 21980
rect 9024 21926 9026 21978
rect 9026 21926 9078 21978
rect 9078 21926 9080 21978
rect 9024 21924 9080 21926
rect 9128 21978 9184 21980
rect 9128 21926 9130 21978
rect 9130 21926 9182 21978
rect 9182 21926 9184 21978
rect 9128 21924 9184 21926
rect 9232 21978 9288 21980
rect 9232 21926 9234 21978
rect 9234 21926 9286 21978
rect 9286 21926 9288 21978
rect 9232 21924 9288 21926
rect 8540 21532 8596 21588
rect 8764 21644 8820 21700
rect 9548 21586 9604 21588
rect 9548 21534 9550 21586
rect 9550 21534 9602 21586
rect 9602 21534 9604 21586
rect 9548 21532 9604 21534
rect 9100 21420 9156 21476
rect 9100 20802 9156 20804
rect 9100 20750 9102 20802
rect 9102 20750 9154 20802
rect 9154 20750 9156 20802
rect 9100 20748 9156 20750
rect 9024 20410 9080 20412
rect 9024 20358 9026 20410
rect 9026 20358 9078 20410
rect 9078 20358 9080 20410
rect 9024 20356 9080 20358
rect 9128 20410 9184 20412
rect 9128 20358 9130 20410
rect 9130 20358 9182 20410
rect 9182 20358 9184 20410
rect 9128 20356 9184 20358
rect 9232 20410 9288 20412
rect 9232 20358 9234 20410
rect 9234 20358 9286 20410
rect 9286 20358 9288 20410
rect 9232 20356 9288 20358
rect 9100 19906 9156 19908
rect 9100 19854 9102 19906
rect 9102 19854 9154 19906
rect 9154 19854 9156 19906
rect 9100 19852 9156 19854
rect 8204 19740 8260 19796
rect 7644 18396 7700 18452
rect 7868 18338 7924 18340
rect 7868 18286 7870 18338
rect 7870 18286 7922 18338
rect 7922 18286 7924 18338
rect 7868 18284 7924 18286
rect 7644 17724 7700 17780
rect 7756 17948 7812 18004
rect 8204 17666 8260 17668
rect 8204 17614 8206 17666
rect 8206 17614 8258 17666
rect 8258 17614 8260 17666
rect 8204 17612 8260 17614
rect 8652 17052 8708 17108
rect 7756 16716 7812 16772
rect 8204 15372 8260 15428
rect 8540 15314 8596 15316
rect 8540 15262 8542 15314
rect 8542 15262 8594 15314
rect 8594 15262 8596 15314
rect 8540 15260 8596 15262
rect 7980 14812 8036 14868
rect 8092 13074 8148 13076
rect 8092 13022 8094 13074
rect 8094 13022 8146 13074
rect 8146 13022 8148 13074
rect 8092 13020 8148 13022
rect 7532 12236 7588 12292
rect 8652 14924 8708 14980
rect 8540 14530 8596 14532
rect 8540 14478 8542 14530
rect 8542 14478 8594 14530
rect 8594 14478 8596 14530
rect 8540 14476 8596 14478
rect 8652 13580 8708 13636
rect 9024 18842 9080 18844
rect 9024 18790 9026 18842
rect 9026 18790 9078 18842
rect 9078 18790 9080 18842
rect 9024 18788 9080 18790
rect 9128 18842 9184 18844
rect 9128 18790 9130 18842
rect 9130 18790 9182 18842
rect 9182 18790 9184 18842
rect 9128 18788 9184 18790
rect 9232 18842 9288 18844
rect 9232 18790 9234 18842
rect 9234 18790 9286 18842
rect 9286 18790 9288 18842
rect 9232 18788 9288 18790
rect 10220 29148 10276 29204
rect 10332 28924 10388 28980
rect 10108 27858 10164 27860
rect 10108 27806 10110 27858
rect 10110 27806 10162 27858
rect 10162 27806 10164 27858
rect 10108 27804 10164 27806
rect 10220 26908 10276 26964
rect 10556 28812 10612 28868
rect 10220 24108 10276 24164
rect 10108 23772 10164 23828
rect 10332 23548 10388 23604
rect 10780 29650 10836 29652
rect 10780 29598 10782 29650
rect 10782 29598 10834 29650
rect 10834 29598 10836 29650
rect 10780 29596 10836 29598
rect 10780 25004 10836 25060
rect 10780 24668 10836 24724
rect 11116 25506 11172 25508
rect 11116 25454 11118 25506
rect 11118 25454 11170 25506
rect 11170 25454 11172 25506
rect 11116 25452 11172 25454
rect 11004 24556 11060 24612
rect 10668 23996 10724 24052
rect 10780 23154 10836 23156
rect 10780 23102 10782 23154
rect 10782 23102 10834 23154
rect 10834 23102 10836 23154
rect 10780 23100 10836 23102
rect 10556 21586 10612 21588
rect 10556 21534 10558 21586
rect 10558 21534 10610 21586
rect 10610 21534 10612 21586
rect 10556 21532 10612 21534
rect 10892 20972 10948 21028
rect 8988 18450 9044 18452
rect 8988 18398 8990 18450
rect 8990 18398 9042 18450
rect 9042 18398 9044 18450
rect 8988 18396 9044 18398
rect 9024 17274 9080 17276
rect 9024 17222 9026 17274
rect 9026 17222 9078 17274
rect 9078 17222 9080 17274
rect 9024 17220 9080 17222
rect 9128 17274 9184 17276
rect 9128 17222 9130 17274
rect 9130 17222 9182 17274
rect 9182 17222 9184 17274
rect 9128 17220 9184 17222
rect 9232 17274 9288 17276
rect 9232 17222 9234 17274
rect 9234 17222 9286 17274
rect 9286 17222 9288 17274
rect 9232 17220 9288 17222
rect 9772 19346 9828 19348
rect 9772 19294 9774 19346
rect 9774 19294 9826 19346
rect 9826 19294 9828 19346
rect 9772 19292 9828 19294
rect 11340 29314 11396 29316
rect 11340 29262 11342 29314
rect 11342 29262 11394 29314
rect 11394 29262 11396 29314
rect 11340 29260 11396 29262
rect 11340 28700 11396 28756
rect 11900 30268 11956 30324
rect 11564 28588 11620 28644
rect 11788 27580 11844 27636
rect 11788 27020 11844 27076
rect 12012 30098 12068 30100
rect 12012 30046 12014 30098
rect 12014 30046 12066 30098
rect 12066 30046 12068 30098
rect 12012 30044 12068 30046
rect 12012 29538 12068 29540
rect 12012 29486 12014 29538
rect 12014 29486 12066 29538
rect 12066 29486 12068 29538
rect 12012 29484 12068 29486
rect 12930 30602 12986 30604
rect 12930 30550 12932 30602
rect 12932 30550 12984 30602
rect 12984 30550 12986 30602
rect 12930 30548 12986 30550
rect 13034 30602 13090 30604
rect 13034 30550 13036 30602
rect 13036 30550 13088 30602
rect 13088 30550 13090 30602
rect 13034 30548 13090 30550
rect 13138 30602 13194 30604
rect 13138 30550 13140 30602
rect 13140 30550 13192 30602
rect 13192 30550 13194 30602
rect 13138 30548 13194 30550
rect 13244 30380 13300 30436
rect 13580 30210 13636 30212
rect 13580 30158 13582 30210
rect 13582 30158 13634 30210
rect 13634 30158 13636 30210
rect 13580 30156 13636 30158
rect 14028 30210 14084 30212
rect 14028 30158 14030 30210
rect 14030 30158 14082 30210
rect 14082 30158 14084 30210
rect 14028 30156 14084 30158
rect 13468 29820 13524 29876
rect 13020 29314 13076 29316
rect 13020 29262 13022 29314
rect 13022 29262 13074 29314
rect 13074 29262 13076 29314
rect 13020 29260 13076 29262
rect 12930 29034 12986 29036
rect 12930 28982 12932 29034
rect 12932 28982 12984 29034
rect 12984 28982 12986 29034
rect 12930 28980 12986 28982
rect 13034 29034 13090 29036
rect 13034 28982 13036 29034
rect 13036 28982 13088 29034
rect 13088 28982 13090 29034
rect 13034 28980 13090 28982
rect 13138 29034 13194 29036
rect 13138 28982 13140 29034
rect 13140 28982 13192 29034
rect 13192 28982 13194 29034
rect 13138 28980 13194 28982
rect 12684 28364 12740 28420
rect 12124 28140 12180 28196
rect 12572 28082 12628 28084
rect 12572 28030 12574 28082
rect 12574 28030 12626 28082
rect 12626 28030 12628 28082
rect 12572 28028 12628 28030
rect 12236 27692 12292 27748
rect 12460 27074 12516 27076
rect 12460 27022 12462 27074
rect 12462 27022 12514 27074
rect 12514 27022 12516 27074
rect 12460 27020 12516 27022
rect 11788 26460 11844 26516
rect 11788 25506 11844 25508
rect 11788 25454 11790 25506
rect 11790 25454 11842 25506
rect 11842 25454 11844 25506
rect 11788 25452 11844 25454
rect 11340 25228 11396 25284
rect 11676 24892 11732 24948
rect 11564 24722 11620 24724
rect 11564 24670 11566 24722
rect 11566 24670 11618 24722
rect 11618 24670 11620 24722
rect 11564 24668 11620 24670
rect 11564 24108 11620 24164
rect 11340 23772 11396 23828
rect 11452 22204 11508 22260
rect 11564 21756 11620 21812
rect 12460 25452 12516 25508
rect 13916 28642 13972 28644
rect 13916 28590 13918 28642
rect 13918 28590 13970 28642
rect 13970 28590 13972 28642
rect 13916 28588 13972 28590
rect 13132 27634 13188 27636
rect 13132 27582 13134 27634
rect 13134 27582 13186 27634
rect 13186 27582 13188 27634
rect 13132 27580 13188 27582
rect 12930 27466 12986 27468
rect 12930 27414 12932 27466
rect 12932 27414 12984 27466
rect 12984 27414 12986 27466
rect 12930 27412 12986 27414
rect 13034 27466 13090 27468
rect 13034 27414 13036 27466
rect 13036 27414 13088 27466
rect 13088 27414 13090 27466
rect 13034 27412 13090 27414
rect 13138 27466 13194 27468
rect 13138 27414 13140 27466
rect 13140 27414 13192 27466
rect 13192 27414 13194 27466
rect 13138 27412 13194 27414
rect 13692 28028 13748 28084
rect 13804 27132 13860 27188
rect 13916 27692 13972 27748
rect 13356 27020 13412 27076
rect 13020 26290 13076 26292
rect 13020 26238 13022 26290
rect 13022 26238 13074 26290
rect 13074 26238 13076 26290
rect 13020 26236 13076 26238
rect 12930 25898 12986 25900
rect 12930 25846 12932 25898
rect 12932 25846 12984 25898
rect 12984 25846 12986 25898
rect 12930 25844 12986 25846
rect 13034 25898 13090 25900
rect 13034 25846 13036 25898
rect 13036 25846 13088 25898
rect 13088 25846 13090 25898
rect 13034 25844 13090 25846
rect 13138 25898 13194 25900
rect 13138 25846 13140 25898
rect 13140 25846 13192 25898
rect 13192 25846 13194 25898
rect 13138 25844 13194 25846
rect 12236 23884 12292 23940
rect 12908 25676 12964 25732
rect 12796 25004 12852 25060
rect 14924 30322 14980 30324
rect 14924 30270 14926 30322
rect 14926 30270 14978 30322
rect 14978 30270 14980 30322
rect 14924 30268 14980 30270
rect 16156 30156 16212 30212
rect 15484 30044 15540 30100
rect 14812 29596 14868 29652
rect 14028 27020 14084 27076
rect 14364 26962 14420 26964
rect 14364 26910 14366 26962
rect 14366 26910 14418 26962
rect 14418 26910 14420 26962
rect 14364 26908 14420 26910
rect 16836 29818 16892 29820
rect 16836 29766 16838 29818
rect 16838 29766 16890 29818
rect 16890 29766 16892 29818
rect 16836 29764 16892 29766
rect 16940 29818 16996 29820
rect 16940 29766 16942 29818
rect 16942 29766 16994 29818
rect 16994 29766 16996 29818
rect 16940 29764 16996 29766
rect 17044 29818 17100 29820
rect 17044 29766 17046 29818
rect 17046 29766 17098 29818
rect 17098 29766 17100 29818
rect 17044 29764 17100 29766
rect 17500 29820 17556 29876
rect 16268 29148 16324 29204
rect 16604 28588 16660 28644
rect 16492 28418 16548 28420
rect 16492 28366 16494 28418
rect 16494 28366 16546 28418
rect 16546 28366 16548 28418
rect 16492 28364 16548 28366
rect 15932 28140 15988 28196
rect 15596 27074 15652 27076
rect 15596 27022 15598 27074
rect 15598 27022 15650 27074
rect 15650 27022 15652 27074
rect 15596 27020 15652 27022
rect 14028 26236 14084 26292
rect 13692 26124 13748 26180
rect 13244 24668 13300 24724
rect 12930 24330 12986 24332
rect 12930 24278 12932 24330
rect 12932 24278 12984 24330
rect 12984 24278 12986 24330
rect 12930 24276 12986 24278
rect 13034 24330 13090 24332
rect 13034 24278 13036 24330
rect 13036 24278 13088 24330
rect 13088 24278 13090 24330
rect 13034 24276 13090 24278
rect 13138 24330 13194 24332
rect 13138 24278 13140 24330
rect 13140 24278 13192 24330
rect 13192 24278 13194 24330
rect 13138 24276 13194 24278
rect 12796 23772 12852 23828
rect 12930 22762 12986 22764
rect 12930 22710 12932 22762
rect 12932 22710 12984 22762
rect 12984 22710 12986 22762
rect 12930 22708 12986 22710
rect 13034 22762 13090 22764
rect 13034 22710 13036 22762
rect 13036 22710 13088 22762
rect 13088 22710 13090 22762
rect 13034 22708 13090 22710
rect 13138 22762 13194 22764
rect 13138 22710 13140 22762
rect 13140 22710 13192 22762
rect 13192 22710 13194 22762
rect 13138 22708 13194 22710
rect 12796 22370 12852 22372
rect 12796 22318 12798 22370
rect 12798 22318 12850 22370
rect 12850 22318 12852 22370
rect 12796 22316 12852 22318
rect 12572 22258 12628 22260
rect 12572 22206 12574 22258
rect 12574 22206 12626 22258
rect 12626 22206 12628 22258
rect 12572 22204 12628 22206
rect 12236 22092 12292 22148
rect 11676 21644 11732 21700
rect 12012 20748 12068 20804
rect 12460 21756 12516 21812
rect 11228 19292 11284 19348
rect 11452 19180 11508 19236
rect 11004 18172 11060 18228
rect 11452 18396 11508 18452
rect 10220 17724 10276 17780
rect 10668 17052 10724 17108
rect 8988 15874 9044 15876
rect 8988 15822 8990 15874
rect 8990 15822 9042 15874
rect 9042 15822 9044 15874
rect 8988 15820 9044 15822
rect 9024 15706 9080 15708
rect 9024 15654 9026 15706
rect 9026 15654 9078 15706
rect 9078 15654 9080 15706
rect 9024 15652 9080 15654
rect 9128 15706 9184 15708
rect 9128 15654 9130 15706
rect 9130 15654 9182 15706
rect 9182 15654 9184 15706
rect 9128 15652 9184 15654
rect 9232 15706 9288 15708
rect 9232 15654 9234 15706
rect 9234 15654 9286 15706
rect 9286 15654 9288 15706
rect 9232 15652 9288 15654
rect 8988 15538 9044 15540
rect 8988 15486 8990 15538
rect 8990 15486 9042 15538
rect 9042 15486 9044 15538
rect 8988 15484 9044 15486
rect 9436 14700 9492 14756
rect 9772 16156 9828 16212
rect 10332 16828 10388 16884
rect 9772 15484 9828 15540
rect 9884 15820 9940 15876
rect 9660 14924 9716 14980
rect 9884 14812 9940 14868
rect 9212 14530 9268 14532
rect 9212 14478 9214 14530
rect 9214 14478 9266 14530
rect 9266 14478 9268 14530
rect 9212 14476 9268 14478
rect 9024 14138 9080 14140
rect 9024 14086 9026 14138
rect 9026 14086 9078 14138
rect 9078 14086 9080 14138
rect 9024 14084 9080 14086
rect 9128 14138 9184 14140
rect 9128 14086 9130 14138
rect 9130 14086 9182 14138
rect 9182 14086 9184 14138
rect 9128 14084 9184 14086
rect 9232 14138 9288 14140
rect 9232 14086 9234 14138
rect 9234 14086 9286 14138
rect 9286 14086 9288 14138
rect 9232 14084 9288 14086
rect 8428 12460 8484 12516
rect 9024 12570 9080 12572
rect 9024 12518 9026 12570
rect 9026 12518 9078 12570
rect 9078 12518 9080 12570
rect 9024 12516 9080 12518
rect 9128 12570 9184 12572
rect 9128 12518 9130 12570
rect 9130 12518 9182 12570
rect 9182 12518 9184 12570
rect 9128 12516 9184 12518
rect 9232 12570 9288 12572
rect 9232 12518 9234 12570
rect 9234 12518 9286 12570
rect 9286 12518 9288 12570
rect 9232 12516 9288 12518
rect 8988 12402 9044 12404
rect 8988 12350 8990 12402
rect 8990 12350 9042 12402
rect 9042 12350 9044 12402
rect 8988 12348 9044 12350
rect 6188 11900 6244 11956
rect 6636 10668 6692 10724
rect 6636 9602 6692 9604
rect 6636 9550 6638 9602
rect 6638 9550 6690 9602
rect 6690 9550 6692 9602
rect 6636 9548 6692 9550
rect 5516 9212 5572 9268
rect 5118 8650 5174 8652
rect 5118 8598 5120 8650
rect 5120 8598 5172 8650
rect 5172 8598 5174 8650
rect 5118 8596 5174 8598
rect 5222 8650 5278 8652
rect 5222 8598 5224 8650
rect 5224 8598 5276 8650
rect 5276 8598 5278 8650
rect 5222 8596 5278 8598
rect 5326 8650 5382 8652
rect 5326 8598 5328 8650
rect 5328 8598 5380 8650
rect 5380 8598 5382 8650
rect 5326 8596 5382 8598
rect 4620 6860 4676 6916
rect 3836 6748 3892 6804
rect 4060 6636 4116 6692
rect 3612 6524 3668 6580
rect 4060 6300 4116 6356
rect 4508 6188 4564 6244
rect 3948 5740 4004 5796
rect 3836 5628 3892 5684
rect 4172 4060 4228 4116
rect 5404 7196 5460 7252
rect 5118 7082 5174 7084
rect 5118 7030 5120 7082
rect 5120 7030 5172 7082
rect 5172 7030 5174 7082
rect 5118 7028 5174 7030
rect 5222 7082 5278 7084
rect 5222 7030 5224 7082
rect 5224 7030 5276 7082
rect 5276 7030 5278 7082
rect 5222 7028 5278 7030
rect 5326 7082 5382 7084
rect 5326 7030 5328 7082
rect 5328 7030 5380 7082
rect 5380 7030 5382 7082
rect 5326 7028 5382 7030
rect 5068 6802 5124 6804
rect 5068 6750 5070 6802
rect 5070 6750 5122 6802
rect 5122 6750 5124 6802
rect 5068 6748 5124 6750
rect 5404 6748 5460 6804
rect 4844 5740 4900 5796
rect 5118 5514 5174 5516
rect 5118 5462 5120 5514
rect 5120 5462 5172 5514
rect 5172 5462 5174 5514
rect 5118 5460 5174 5462
rect 5222 5514 5278 5516
rect 5222 5462 5224 5514
rect 5224 5462 5276 5514
rect 5276 5462 5278 5514
rect 5222 5460 5278 5462
rect 5326 5514 5382 5516
rect 5326 5462 5328 5514
rect 5328 5462 5380 5514
rect 5380 5462 5382 5514
rect 5326 5460 5382 5462
rect 5628 6578 5684 6580
rect 5628 6526 5630 6578
rect 5630 6526 5682 6578
rect 5682 6526 5684 6578
rect 5628 6524 5684 6526
rect 5628 5852 5684 5908
rect 5068 4898 5124 4900
rect 5068 4846 5070 4898
rect 5070 4846 5122 4898
rect 5122 4846 5124 4898
rect 5068 4844 5124 4846
rect 4732 4508 4788 4564
rect 6300 6748 6356 6804
rect 6076 5628 6132 5684
rect 6412 5404 6468 5460
rect 6300 5010 6356 5012
rect 6300 4958 6302 5010
rect 6302 4958 6354 5010
rect 6354 4958 6356 5010
rect 6300 4956 6356 4958
rect 5740 4732 5796 4788
rect 5740 4396 5796 4452
rect 5118 3946 5174 3948
rect 5118 3894 5120 3946
rect 5120 3894 5172 3946
rect 5172 3894 5174 3946
rect 5118 3892 5174 3894
rect 5222 3946 5278 3948
rect 5222 3894 5224 3946
rect 5224 3894 5276 3946
rect 5276 3894 5278 3946
rect 5222 3892 5278 3894
rect 5326 3946 5382 3948
rect 5326 3894 5328 3946
rect 5328 3894 5380 3946
rect 5380 3894 5382 3946
rect 5326 3892 5382 3894
rect 5068 3724 5124 3780
rect 4620 3666 4676 3668
rect 4620 3614 4622 3666
rect 4622 3614 4674 3666
rect 4674 3614 4676 3666
rect 4620 3612 4676 3614
rect 8428 10780 8484 10836
rect 7308 10668 7364 10724
rect 8316 10668 8372 10724
rect 6748 7308 6804 7364
rect 6636 7196 6692 7252
rect 6860 6690 6916 6692
rect 6860 6638 6862 6690
rect 6862 6638 6914 6690
rect 6914 6638 6916 6690
rect 6860 6636 6916 6638
rect 7420 6076 7476 6132
rect 7532 6636 7588 6692
rect 7196 5906 7252 5908
rect 7196 5854 7198 5906
rect 7198 5854 7250 5906
rect 7250 5854 7252 5906
rect 7196 5852 7252 5854
rect 7532 5906 7588 5908
rect 7532 5854 7534 5906
rect 7534 5854 7586 5906
rect 7586 5854 7588 5906
rect 7532 5852 7588 5854
rect 7196 5516 7252 5572
rect 6748 4844 6804 4900
rect 4508 3500 4564 3556
rect 6076 3500 6132 3556
rect 4172 3276 4228 3332
rect 3500 2044 3556 2100
rect 7532 4732 7588 4788
rect 8092 6130 8148 6132
rect 8092 6078 8094 6130
rect 8094 6078 8146 6130
rect 8146 6078 8148 6130
rect 8092 6076 8148 6078
rect 8316 9826 8372 9828
rect 8316 9774 8318 9826
rect 8318 9774 8370 9826
rect 8370 9774 8372 9826
rect 8316 9772 8372 9774
rect 8316 9548 8372 9604
rect 9436 11394 9492 11396
rect 9436 11342 9438 11394
rect 9438 11342 9490 11394
rect 9490 11342 9492 11394
rect 9436 11340 9492 11342
rect 9024 11002 9080 11004
rect 9024 10950 9026 11002
rect 9026 10950 9078 11002
rect 9078 10950 9080 11002
rect 9024 10948 9080 10950
rect 9128 11002 9184 11004
rect 9128 10950 9130 11002
rect 9130 10950 9182 11002
rect 9182 10950 9184 11002
rect 9128 10948 9184 10950
rect 9232 11002 9288 11004
rect 9232 10950 9234 11002
rect 9234 10950 9286 11002
rect 9286 10950 9288 11002
rect 9232 10948 9288 10950
rect 9996 14476 10052 14532
rect 10108 13580 10164 13636
rect 9996 12348 10052 12404
rect 10108 10834 10164 10836
rect 10108 10782 10110 10834
rect 10110 10782 10162 10834
rect 10162 10782 10164 10834
rect 10108 10780 10164 10782
rect 9024 9434 9080 9436
rect 9024 9382 9026 9434
rect 9026 9382 9078 9434
rect 9078 9382 9080 9434
rect 9024 9380 9080 9382
rect 9128 9434 9184 9436
rect 9128 9382 9130 9434
rect 9130 9382 9182 9434
rect 9182 9382 9184 9434
rect 9128 9380 9184 9382
rect 9232 9434 9288 9436
rect 9232 9382 9234 9434
rect 9234 9382 9286 9434
rect 9286 9382 9288 9434
rect 9232 9380 9288 9382
rect 8540 8988 8596 9044
rect 8764 8204 8820 8260
rect 8652 8034 8708 8036
rect 8652 7982 8654 8034
rect 8654 7982 8706 8034
rect 8706 7982 8708 8034
rect 8652 7980 8708 7982
rect 9548 9154 9604 9156
rect 9548 9102 9550 9154
rect 9550 9102 9602 9154
rect 9602 9102 9604 9154
rect 9548 9100 9604 9102
rect 9100 8092 9156 8148
rect 9024 7866 9080 7868
rect 9024 7814 9026 7866
rect 9026 7814 9078 7866
rect 9078 7814 9080 7866
rect 9024 7812 9080 7814
rect 9128 7866 9184 7868
rect 9128 7814 9130 7866
rect 9130 7814 9182 7866
rect 9182 7814 9184 7866
rect 9128 7812 9184 7814
rect 9232 7866 9288 7868
rect 9232 7814 9234 7866
rect 9234 7814 9286 7866
rect 9286 7814 9288 7866
rect 9232 7812 9288 7814
rect 9024 6298 9080 6300
rect 9024 6246 9026 6298
rect 9026 6246 9078 6298
rect 9078 6246 9080 6298
rect 9024 6244 9080 6246
rect 9128 6298 9184 6300
rect 9128 6246 9130 6298
rect 9130 6246 9182 6298
rect 9182 6246 9184 6298
rect 9128 6244 9184 6246
rect 9232 6298 9288 6300
rect 9232 6246 9234 6298
rect 9234 6246 9286 6298
rect 9286 6246 9288 6298
rect 9232 6244 9288 6246
rect 8316 5852 8372 5908
rect 8092 5516 8148 5572
rect 8204 4898 8260 4900
rect 8204 4846 8206 4898
rect 8206 4846 8258 4898
rect 8258 4846 8260 4898
rect 8204 4844 8260 4846
rect 9772 7868 9828 7924
rect 9996 7868 10052 7924
rect 11004 17164 11060 17220
rect 10892 16940 10948 16996
rect 12572 21308 12628 21364
rect 12930 21194 12986 21196
rect 12930 21142 12932 21194
rect 12932 21142 12984 21194
rect 12984 21142 12986 21194
rect 12930 21140 12986 21142
rect 13034 21194 13090 21196
rect 13034 21142 13036 21194
rect 13036 21142 13088 21194
rect 13088 21142 13090 21194
rect 13034 21140 13090 21142
rect 13138 21194 13194 21196
rect 13138 21142 13140 21194
rect 13140 21142 13192 21194
rect 13192 21142 13194 21194
rect 13138 21140 13194 21142
rect 12796 20690 12852 20692
rect 12796 20638 12798 20690
rect 12798 20638 12850 20690
rect 12850 20638 12852 20690
rect 12796 20636 12852 20638
rect 13580 22370 13636 22372
rect 13580 22318 13582 22370
rect 13582 22318 13634 22370
rect 13634 22318 13636 22370
rect 13580 22316 13636 22318
rect 14028 25676 14084 25732
rect 14588 25730 14644 25732
rect 14588 25678 14590 25730
rect 14590 25678 14642 25730
rect 14642 25678 14644 25730
rect 14588 25676 14644 25678
rect 13804 25506 13860 25508
rect 13804 25454 13806 25506
rect 13806 25454 13858 25506
rect 13858 25454 13860 25506
rect 13804 25452 13860 25454
rect 13916 25228 13972 25284
rect 13916 23938 13972 23940
rect 13916 23886 13918 23938
rect 13918 23886 13970 23938
rect 13970 23886 13972 23938
rect 13916 23884 13972 23886
rect 15260 25506 15316 25508
rect 15260 25454 15262 25506
rect 15262 25454 15314 25506
rect 15314 25454 15316 25506
rect 15260 25452 15316 25454
rect 14812 24780 14868 24836
rect 14700 24556 14756 24612
rect 14140 23436 14196 23492
rect 15484 24946 15540 24948
rect 15484 24894 15486 24946
rect 15486 24894 15538 24946
rect 15538 24894 15540 24946
rect 15484 24892 15540 24894
rect 15260 24834 15316 24836
rect 15260 24782 15262 24834
rect 15262 24782 15314 24834
rect 15314 24782 15316 24834
rect 15260 24780 15316 24782
rect 16268 26908 16324 26964
rect 17052 29484 17108 29540
rect 17164 28812 17220 28868
rect 16836 28250 16892 28252
rect 16836 28198 16838 28250
rect 16838 28198 16890 28250
rect 16890 28198 16892 28250
rect 16836 28196 16892 28198
rect 16940 28250 16996 28252
rect 16940 28198 16942 28250
rect 16942 28198 16994 28250
rect 16994 28198 16996 28250
rect 16940 28196 16996 28198
rect 17044 28250 17100 28252
rect 17044 28198 17046 28250
rect 17046 28198 17098 28250
rect 17098 28198 17100 28250
rect 17044 28196 17100 28198
rect 16380 26796 16436 26852
rect 17164 27804 17220 27860
rect 16380 26348 16436 26404
rect 13804 20972 13860 21028
rect 13916 22316 13972 22372
rect 15036 22370 15092 22372
rect 15036 22318 15038 22370
rect 15038 22318 15090 22370
rect 15090 22318 15092 22370
rect 15036 22316 15092 22318
rect 13804 20802 13860 20804
rect 13804 20750 13806 20802
rect 13806 20750 13858 20802
rect 13858 20750 13860 20802
rect 13804 20748 13860 20750
rect 12930 19626 12986 19628
rect 12930 19574 12932 19626
rect 12932 19574 12984 19626
rect 12984 19574 12986 19626
rect 12930 19572 12986 19574
rect 13034 19626 13090 19628
rect 13034 19574 13036 19626
rect 13036 19574 13088 19626
rect 13088 19574 13090 19626
rect 13034 19572 13090 19574
rect 13138 19626 13194 19628
rect 13138 19574 13140 19626
rect 13140 19574 13192 19626
rect 13192 19574 13194 19626
rect 13138 19572 13194 19574
rect 12908 19346 12964 19348
rect 12908 19294 12910 19346
rect 12910 19294 12962 19346
rect 12962 19294 12964 19346
rect 12908 19292 12964 19294
rect 11676 18284 11732 18340
rect 11788 18172 11844 18228
rect 11564 17164 11620 17220
rect 14476 19740 14532 19796
rect 13692 19292 13748 19348
rect 13020 18450 13076 18452
rect 13020 18398 13022 18450
rect 13022 18398 13074 18450
rect 13074 18398 13076 18450
rect 13020 18396 13076 18398
rect 13916 18450 13972 18452
rect 13916 18398 13918 18450
rect 13918 18398 13970 18450
rect 13970 18398 13972 18450
rect 13916 18396 13972 18398
rect 14364 18172 14420 18228
rect 12012 18060 12068 18116
rect 11228 16098 11284 16100
rect 11228 16046 11230 16098
rect 11230 16046 11282 16098
rect 11282 16046 11284 16098
rect 11228 16044 11284 16046
rect 12930 18058 12986 18060
rect 12930 18006 12932 18058
rect 12932 18006 12984 18058
rect 12984 18006 12986 18058
rect 12930 18004 12986 18006
rect 13034 18058 13090 18060
rect 13034 18006 13036 18058
rect 13036 18006 13088 18058
rect 13088 18006 13090 18058
rect 13034 18004 13090 18006
rect 13138 18058 13194 18060
rect 13138 18006 13140 18058
rect 13140 18006 13192 18058
rect 13192 18006 13194 18058
rect 13138 18004 13194 18006
rect 12124 17778 12180 17780
rect 12124 17726 12126 17778
rect 12126 17726 12178 17778
rect 12178 17726 12180 17778
rect 12124 17724 12180 17726
rect 12348 17164 12404 17220
rect 12908 17164 12964 17220
rect 13580 17164 13636 17220
rect 12572 16828 12628 16884
rect 11116 15314 11172 15316
rect 11116 15262 11118 15314
rect 11118 15262 11170 15314
rect 11170 15262 11172 15314
rect 11116 15260 11172 15262
rect 10892 14252 10948 14308
rect 11676 13580 11732 13636
rect 11900 13692 11956 13748
rect 12930 16490 12986 16492
rect 12930 16438 12932 16490
rect 12932 16438 12984 16490
rect 12984 16438 12986 16490
rect 12930 16436 12986 16438
rect 13034 16490 13090 16492
rect 13034 16438 13036 16490
rect 13036 16438 13088 16490
rect 13088 16438 13090 16490
rect 13034 16436 13090 16438
rect 13138 16490 13194 16492
rect 13138 16438 13140 16490
rect 13140 16438 13192 16490
rect 13192 16438 13194 16490
rect 13138 16436 13194 16438
rect 14364 17106 14420 17108
rect 14364 17054 14366 17106
rect 14366 17054 14418 17106
rect 14418 17054 14420 17106
rect 14364 17052 14420 17054
rect 13020 16210 13076 16212
rect 13020 16158 13022 16210
rect 13022 16158 13074 16210
rect 13074 16158 13076 16210
rect 13020 16156 13076 16158
rect 14924 20748 14980 20804
rect 15148 20802 15204 20804
rect 15148 20750 15150 20802
rect 15150 20750 15202 20802
rect 15202 20750 15204 20802
rect 15148 20748 15204 20750
rect 15260 23996 15316 24052
rect 16380 23212 16436 23268
rect 14924 16658 14980 16660
rect 14924 16606 14926 16658
rect 14926 16606 14978 16658
rect 14978 16606 14980 16658
rect 14924 16604 14980 16606
rect 14812 16156 14868 16212
rect 16836 26682 16892 26684
rect 16836 26630 16838 26682
rect 16838 26630 16890 26682
rect 16890 26630 16892 26682
rect 16836 26628 16892 26630
rect 16940 26682 16996 26684
rect 16940 26630 16942 26682
rect 16942 26630 16994 26682
rect 16994 26630 16996 26682
rect 16940 26628 16996 26630
rect 17044 26682 17100 26684
rect 17044 26630 17046 26682
rect 17046 26630 17098 26682
rect 17098 26630 17100 26682
rect 17044 26628 17100 26630
rect 17276 26908 17332 26964
rect 17724 29260 17780 29316
rect 18172 30156 18228 30212
rect 20742 30602 20798 30604
rect 20742 30550 20744 30602
rect 20744 30550 20796 30602
rect 20796 30550 20798 30602
rect 20742 30548 20798 30550
rect 20846 30602 20902 30604
rect 20846 30550 20848 30602
rect 20848 30550 20900 30602
rect 20900 30550 20902 30602
rect 20846 30548 20902 30550
rect 20950 30602 21006 30604
rect 20950 30550 20952 30602
rect 20952 30550 21004 30602
rect 21004 30550 21006 30602
rect 20950 30548 21006 30550
rect 19964 30210 20020 30212
rect 19964 30158 19966 30210
rect 19966 30158 20018 30210
rect 20018 30158 20020 30210
rect 19964 30156 20020 30158
rect 21420 30210 21476 30212
rect 21420 30158 21422 30210
rect 21422 30158 21474 30210
rect 21474 30158 21476 30210
rect 21420 30156 21476 30158
rect 17948 28588 18004 28644
rect 18844 28252 18900 28308
rect 18732 27746 18788 27748
rect 18732 27694 18734 27746
rect 18734 27694 18786 27746
rect 18786 27694 18788 27746
rect 18732 27692 18788 27694
rect 17388 26402 17444 26404
rect 17388 26350 17390 26402
rect 17390 26350 17442 26402
rect 17442 26350 17444 26402
rect 17388 26348 17444 26350
rect 16828 25676 16884 25732
rect 17612 25676 17668 25732
rect 16604 24892 16660 24948
rect 16836 25114 16892 25116
rect 16836 25062 16838 25114
rect 16838 25062 16890 25114
rect 16890 25062 16892 25114
rect 16836 25060 16892 25062
rect 16940 25114 16996 25116
rect 16940 25062 16942 25114
rect 16942 25062 16994 25114
rect 16994 25062 16996 25114
rect 16940 25060 16996 25062
rect 17044 25114 17100 25116
rect 17044 25062 17046 25114
rect 17046 25062 17098 25114
rect 17098 25062 17100 25114
rect 17044 25060 17100 25062
rect 17724 24668 17780 24724
rect 17836 25564 17892 25620
rect 17612 24610 17668 24612
rect 17612 24558 17614 24610
rect 17614 24558 17666 24610
rect 17666 24558 17668 24610
rect 17612 24556 17668 24558
rect 16836 23546 16892 23548
rect 16836 23494 16838 23546
rect 16838 23494 16890 23546
rect 16890 23494 16892 23546
rect 16836 23492 16892 23494
rect 16940 23546 16996 23548
rect 16940 23494 16942 23546
rect 16942 23494 16994 23546
rect 16994 23494 16996 23546
rect 16940 23492 16996 23494
rect 17044 23546 17100 23548
rect 17044 23494 17046 23546
rect 17046 23494 17098 23546
rect 17098 23494 17100 23546
rect 17044 23492 17100 23494
rect 16716 23100 16772 23156
rect 16156 22092 16212 22148
rect 17724 23378 17780 23380
rect 17724 23326 17726 23378
rect 17726 23326 17778 23378
rect 17778 23326 17780 23378
rect 17724 23324 17780 23326
rect 17164 22092 17220 22148
rect 16836 21978 16892 21980
rect 16836 21926 16838 21978
rect 16838 21926 16890 21978
rect 16890 21926 16892 21978
rect 16836 21924 16892 21926
rect 16940 21978 16996 21980
rect 16940 21926 16942 21978
rect 16942 21926 16994 21978
rect 16994 21926 16996 21978
rect 16940 21924 16996 21926
rect 17044 21978 17100 21980
rect 17044 21926 17046 21978
rect 17046 21926 17098 21978
rect 17098 21926 17100 21978
rect 17044 21924 17100 21926
rect 16268 21756 16324 21812
rect 17500 20860 17556 20916
rect 16836 20410 16892 20412
rect 16836 20358 16838 20410
rect 16838 20358 16890 20410
rect 16890 20358 16892 20410
rect 16836 20356 16892 20358
rect 16940 20410 16996 20412
rect 16940 20358 16942 20410
rect 16942 20358 16994 20410
rect 16994 20358 16996 20410
rect 16940 20356 16996 20358
rect 17044 20410 17100 20412
rect 17044 20358 17046 20410
rect 17046 20358 17098 20410
rect 17098 20358 17100 20410
rect 17044 20356 17100 20358
rect 15932 20130 15988 20132
rect 15932 20078 15934 20130
rect 15934 20078 15986 20130
rect 15986 20078 15988 20130
rect 15932 20076 15988 20078
rect 16716 19404 16772 19460
rect 15372 17612 15428 17668
rect 15484 17164 15540 17220
rect 15260 16994 15316 16996
rect 15260 16942 15262 16994
rect 15262 16942 15314 16994
rect 15314 16942 15316 16994
rect 15260 16940 15316 16942
rect 15932 16882 15988 16884
rect 15932 16830 15934 16882
rect 15934 16830 15986 16882
rect 15986 16830 15988 16882
rect 15932 16828 15988 16830
rect 16604 18508 16660 18564
rect 16380 17052 16436 17108
rect 16836 18842 16892 18844
rect 16836 18790 16838 18842
rect 16838 18790 16890 18842
rect 16890 18790 16892 18842
rect 16836 18788 16892 18790
rect 16940 18842 16996 18844
rect 16940 18790 16942 18842
rect 16942 18790 16994 18842
rect 16994 18790 16996 18842
rect 16940 18788 16996 18790
rect 17044 18842 17100 18844
rect 17044 18790 17046 18842
rect 17046 18790 17098 18842
rect 17098 18790 17100 18842
rect 17044 18788 17100 18790
rect 16940 18226 16996 18228
rect 16940 18174 16942 18226
rect 16942 18174 16994 18226
rect 16994 18174 16996 18226
rect 16940 18172 16996 18174
rect 17164 17666 17220 17668
rect 17164 17614 17166 17666
rect 17166 17614 17218 17666
rect 17218 17614 17220 17666
rect 17164 17612 17220 17614
rect 16836 17274 16892 17276
rect 16836 17222 16838 17274
rect 16838 17222 16890 17274
rect 16890 17222 16892 17274
rect 16836 17220 16892 17222
rect 16940 17274 16996 17276
rect 16940 17222 16942 17274
rect 16942 17222 16994 17274
rect 16994 17222 16996 17274
rect 16940 17220 16996 17222
rect 17044 17274 17100 17276
rect 17044 17222 17046 17274
rect 17046 17222 17098 17274
rect 17098 17222 17100 17274
rect 17044 17220 17100 17222
rect 16828 16828 16884 16884
rect 15820 16604 15876 16660
rect 15148 15484 15204 15540
rect 12930 14922 12986 14924
rect 12930 14870 12932 14922
rect 12932 14870 12984 14922
rect 12984 14870 12986 14922
rect 12930 14868 12986 14870
rect 13034 14922 13090 14924
rect 13034 14870 13036 14922
rect 13036 14870 13088 14922
rect 13088 14870 13090 14922
rect 13034 14868 13090 14870
rect 13138 14922 13194 14924
rect 13138 14870 13140 14922
rect 13140 14870 13192 14922
rect 13192 14870 13194 14922
rect 14700 14924 14756 14980
rect 13138 14868 13194 14870
rect 12460 14588 12516 14644
rect 12348 14476 12404 14532
rect 13020 14306 13076 14308
rect 13020 14254 13022 14306
rect 13022 14254 13074 14306
rect 13074 14254 13076 14306
rect 13020 14252 13076 14254
rect 13692 13746 13748 13748
rect 13692 13694 13694 13746
rect 13694 13694 13746 13746
rect 13746 13694 13748 13746
rect 13692 13692 13748 13694
rect 14476 13692 14532 13748
rect 16380 14588 16436 14644
rect 15260 13692 15316 13748
rect 16156 13692 16212 13748
rect 12796 13634 12852 13636
rect 12796 13582 12798 13634
rect 12798 13582 12850 13634
rect 12850 13582 12852 13634
rect 12796 13580 12852 13582
rect 12930 13354 12986 13356
rect 12930 13302 12932 13354
rect 12932 13302 12984 13354
rect 12984 13302 12986 13354
rect 12930 13300 12986 13302
rect 13034 13354 13090 13356
rect 13034 13302 13036 13354
rect 13036 13302 13088 13354
rect 13088 13302 13090 13354
rect 13034 13300 13090 13302
rect 13138 13354 13194 13356
rect 13138 13302 13140 13354
rect 13140 13302 13192 13354
rect 13192 13302 13194 13354
rect 13138 13300 13194 13302
rect 13692 13244 13748 13300
rect 12460 13020 12516 13076
rect 13580 13074 13636 13076
rect 13580 13022 13582 13074
rect 13582 13022 13634 13074
rect 13634 13022 13636 13074
rect 13580 13020 13636 13022
rect 12012 12796 12068 12852
rect 15372 13244 15428 13300
rect 11676 12124 11732 12180
rect 12908 12738 12964 12740
rect 12908 12686 12910 12738
rect 12910 12686 12962 12738
rect 12962 12686 12964 12738
rect 12908 12684 12964 12686
rect 14588 12908 14644 12964
rect 13692 12684 13748 12740
rect 10892 11340 10948 11396
rect 10556 10834 10612 10836
rect 10556 10782 10558 10834
rect 10558 10782 10610 10834
rect 10610 10782 10612 10834
rect 10556 10780 10612 10782
rect 12930 11786 12986 11788
rect 12930 11734 12932 11786
rect 12932 11734 12984 11786
rect 12984 11734 12986 11786
rect 12930 11732 12986 11734
rect 13034 11786 13090 11788
rect 13034 11734 13036 11786
rect 13036 11734 13088 11786
rect 13088 11734 13090 11786
rect 13034 11732 13090 11734
rect 13138 11786 13194 11788
rect 13138 11734 13140 11786
rect 13140 11734 13192 11786
rect 13192 11734 13194 11786
rect 13138 11732 13194 11734
rect 12908 11394 12964 11396
rect 12908 11342 12910 11394
rect 12910 11342 12962 11394
rect 12962 11342 12964 11394
rect 12908 11340 12964 11342
rect 11676 10780 11732 10836
rect 13468 11116 13524 11172
rect 10444 9266 10500 9268
rect 10444 9214 10446 9266
rect 10446 9214 10498 9266
rect 10498 9214 10500 9266
rect 10444 9212 10500 9214
rect 10892 10332 10948 10388
rect 13468 10332 13524 10388
rect 14364 12178 14420 12180
rect 14364 12126 14366 12178
rect 14366 12126 14418 12178
rect 14418 12126 14420 12178
rect 14364 12124 14420 12126
rect 12930 10218 12986 10220
rect 12930 10166 12932 10218
rect 12932 10166 12984 10218
rect 12984 10166 12986 10218
rect 12930 10164 12986 10166
rect 13034 10218 13090 10220
rect 13034 10166 13036 10218
rect 13036 10166 13088 10218
rect 13088 10166 13090 10218
rect 13034 10164 13090 10166
rect 13138 10218 13194 10220
rect 13138 10166 13140 10218
rect 13140 10166 13192 10218
rect 13192 10166 13194 10218
rect 13138 10164 13194 10166
rect 10892 9772 10948 9828
rect 10668 8876 10724 8932
rect 9772 6412 9828 6468
rect 9548 6130 9604 6132
rect 9548 6078 9550 6130
rect 9550 6078 9602 6130
rect 9602 6078 9604 6130
rect 9548 6076 9604 6078
rect 9436 5292 9492 5348
rect 8764 4956 8820 5012
rect 9024 4730 9080 4732
rect 9024 4678 9026 4730
rect 9026 4678 9078 4730
rect 9078 4678 9080 4730
rect 9024 4676 9080 4678
rect 9128 4730 9184 4732
rect 9128 4678 9130 4730
rect 9130 4678 9182 4730
rect 9182 4678 9184 4730
rect 9128 4676 9184 4678
rect 9232 4730 9288 4732
rect 9232 4678 9234 4730
rect 9234 4678 9286 4730
rect 9286 4678 9288 4730
rect 9232 4676 9288 4678
rect 9660 4508 9716 4564
rect 8652 3442 8708 3444
rect 8652 3390 8654 3442
rect 8654 3390 8706 3442
rect 8706 3390 8708 3442
rect 8652 3388 8708 3390
rect 10332 6690 10388 6692
rect 10332 6638 10334 6690
rect 10334 6638 10386 6690
rect 10386 6638 10388 6690
rect 10332 6636 10388 6638
rect 10444 6076 10500 6132
rect 10780 9324 10836 9380
rect 11340 9772 11396 9828
rect 11228 9266 11284 9268
rect 11228 9214 11230 9266
rect 11230 9214 11282 9266
rect 11282 9214 11284 9266
rect 11228 9212 11284 9214
rect 11228 7868 11284 7924
rect 12460 9548 12516 9604
rect 12236 8092 12292 8148
rect 11340 6860 11396 6916
rect 10780 6690 10836 6692
rect 10780 6638 10782 6690
rect 10782 6638 10834 6690
rect 10834 6638 10836 6690
rect 10780 6636 10836 6638
rect 11676 6636 11732 6692
rect 10668 6524 10724 6580
rect 10108 5068 10164 5124
rect 10108 4844 10164 4900
rect 13580 9602 13636 9604
rect 13580 9550 13582 9602
rect 13582 9550 13634 9602
rect 13634 9550 13636 9602
rect 13580 9548 13636 9550
rect 13468 9212 13524 9268
rect 13244 8876 13300 8932
rect 12930 8650 12986 8652
rect 12930 8598 12932 8650
rect 12932 8598 12984 8650
rect 12984 8598 12986 8650
rect 12930 8596 12986 8598
rect 13034 8650 13090 8652
rect 13034 8598 13036 8650
rect 13036 8598 13088 8650
rect 13088 8598 13090 8650
rect 13034 8596 13090 8598
rect 13138 8650 13194 8652
rect 13138 8598 13140 8650
rect 13140 8598 13192 8650
rect 13192 8598 13194 8650
rect 13138 8596 13194 8598
rect 12930 7082 12986 7084
rect 12930 7030 12932 7082
rect 12932 7030 12984 7082
rect 12984 7030 12986 7082
rect 12930 7028 12986 7030
rect 13034 7082 13090 7084
rect 13034 7030 13036 7082
rect 13036 7030 13088 7082
rect 13088 7030 13090 7082
rect 13034 7028 13090 7030
rect 13138 7082 13194 7084
rect 13138 7030 13140 7082
rect 13140 7030 13192 7082
rect 13192 7030 13194 7082
rect 13138 7028 13194 7030
rect 12124 3554 12180 3556
rect 12124 3502 12126 3554
rect 12126 3502 12178 3554
rect 12178 3502 12180 3554
rect 12124 3500 12180 3502
rect 9024 3162 9080 3164
rect 9024 3110 9026 3162
rect 9026 3110 9078 3162
rect 9078 3110 9080 3162
rect 9024 3108 9080 3110
rect 9128 3162 9184 3164
rect 9128 3110 9130 3162
rect 9130 3110 9182 3162
rect 9182 3110 9184 3162
rect 9128 3108 9184 3110
rect 9232 3162 9288 3164
rect 9232 3110 9234 3162
rect 9234 3110 9286 3162
rect 9286 3110 9288 3162
rect 9232 3108 9288 3110
rect 12572 5404 12628 5460
rect 13468 5964 13524 6020
rect 15148 12178 15204 12180
rect 15148 12126 15150 12178
rect 15150 12126 15202 12178
rect 15202 12126 15204 12178
rect 15148 12124 15204 12126
rect 14924 12066 14980 12068
rect 14924 12014 14926 12066
rect 14926 12014 14978 12066
rect 14978 12014 14980 12066
rect 14924 12012 14980 12014
rect 14700 11452 14756 11508
rect 15260 11954 15316 11956
rect 15260 11902 15262 11954
rect 15262 11902 15314 11954
rect 15314 11902 15316 11954
rect 15260 11900 15316 11902
rect 15372 11676 15428 11732
rect 15260 10498 15316 10500
rect 15260 10446 15262 10498
rect 15262 10446 15314 10498
rect 15314 10446 15316 10498
rect 15260 10444 15316 10446
rect 14028 9660 14084 9716
rect 14812 9660 14868 9716
rect 14252 9212 14308 9268
rect 13804 8876 13860 8932
rect 14252 8316 14308 8372
rect 14028 7084 14084 7140
rect 14476 6018 14532 6020
rect 14476 5966 14478 6018
rect 14478 5966 14530 6018
rect 14530 5966 14532 6018
rect 14476 5964 14532 5966
rect 13916 5852 13972 5908
rect 12930 5514 12986 5516
rect 12930 5462 12932 5514
rect 12932 5462 12984 5514
rect 12984 5462 12986 5514
rect 12930 5460 12986 5462
rect 13034 5514 13090 5516
rect 13034 5462 13036 5514
rect 13036 5462 13088 5514
rect 13088 5462 13090 5514
rect 13034 5460 13090 5462
rect 13138 5514 13194 5516
rect 13138 5462 13140 5514
rect 13140 5462 13192 5514
rect 13192 5462 13194 5514
rect 13138 5460 13194 5462
rect 12572 5122 12628 5124
rect 12572 5070 12574 5122
rect 12574 5070 12626 5122
rect 12626 5070 12628 5122
rect 12572 5068 12628 5070
rect 13916 5122 13972 5124
rect 13916 5070 13918 5122
rect 13918 5070 13970 5122
rect 13970 5070 13972 5122
rect 13916 5068 13972 5070
rect 12796 4338 12852 4340
rect 12796 4286 12798 4338
rect 12798 4286 12850 4338
rect 12850 4286 12852 4338
rect 12796 4284 12852 4286
rect 13244 4060 13300 4116
rect 12930 3946 12986 3948
rect 12930 3894 12932 3946
rect 12932 3894 12984 3946
rect 12984 3894 12986 3946
rect 12930 3892 12986 3894
rect 13034 3946 13090 3948
rect 13034 3894 13036 3946
rect 13036 3894 13088 3946
rect 13088 3894 13090 3946
rect 13034 3892 13090 3894
rect 13138 3946 13194 3948
rect 13138 3894 13140 3946
rect 13140 3894 13192 3946
rect 13192 3894 13194 3946
rect 13138 3892 13194 3894
rect 14140 4898 14196 4900
rect 14140 4846 14142 4898
rect 14142 4846 14194 4898
rect 14194 4846 14196 4898
rect 14140 4844 14196 4846
rect 13356 3554 13412 3556
rect 13356 3502 13358 3554
rect 13358 3502 13410 3554
rect 13410 3502 13412 3554
rect 13356 3500 13412 3502
rect 13132 3442 13188 3444
rect 13132 3390 13134 3442
rect 13134 3390 13186 3442
rect 13186 3390 13188 3442
rect 13132 3388 13188 3390
rect 14812 9100 14868 9156
rect 15260 8428 15316 8484
rect 15036 8316 15092 8372
rect 16604 15148 16660 15204
rect 16604 13692 16660 13748
rect 16492 13244 16548 13300
rect 16836 15706 16892 15708
rect 16836 15654 16838 15706
rect 16838 15654 16890 15706
rect 16890 15654 16892 15706
rect 16836 15652 16892 15654
rect 16940 15706 16996 15708
rect 16940 15654 16942 15706
rect 16942 15654 16994 15706
rect 16994 15654 16996 15706
rect 16940 15652 16996 15654
rect 17044 15706 17100 15708
rect 17044 15654 17046 15706
rect 17046 15654 17098 15706
rect 17098 15654 17100 15706
rect 17044 15652 17100 15654
rect 17052 15036 17108 15092
rect 17612 19852 17668 19908
rect 17612 18060 17668 18116
rect 17612 17388 17668 17444
rect 17500 16882 17556 16884
rect 17500 16830 17502 16882
rect 17502 16830 17554 16882
rect 17554 16830 17556 16882
rect 17500 16828 17556 16830
rect 18060 26796 18116 26852
rect 18284 26796 18340 26852
rect 18060 23266 18116 23268
rect 18060 23214 18062 23266
rect 18062 23214 18114 23266
rect 18114 23214 18116 23266
rect 18060 23212 18116 23214
rect 20188 30044 20244 30100
rect 19404 29932 19460 29988
rect 19180 27804 19236 27860
rect 19292 25618 19348 25620
rect 19292 25566 19294 25618
rect 19294 25566 19346 25618
rect 19346 25566 19348 25618
rect 19292 25564 19348 25566
rect 18396 24722 18452 24724
rect 18396 24670 18398 24722
rect 18398 24670 18450 24722
rect 18450 24670 18452 24722
rect 18396 24668 18452 24670
rect 18956 24722 19012 24724
rect 18956 24670 18958 24722
rect 18958 24670 19010 24722
rect 19010 24670 19012 24722
rect 18956 24668 19012 24670
rect 18732 23266 18788 23268
rect 18732 23214 18734 23266
rect 18734 23214 18786 23266
rect 18786 23214 18788 23266
rect 18732 23212 18788 23214
rect 18396 22092 18452 22148
rect 18060 21810 18116 21812
rect 18060 21758 18062 21810
rect 18062 21758 18114 21810
rect 18114 21758 18116 21810
rect 18060 21756 18116 21758
rect 17948 20636 18004 20692
rect 18956 21586 19012 21588
rect 18956 21534 18958 21586
rect 18958 21534 19010 21586
rect 19010 21534 19012 21586
rect 18956 21532 19012 21534
rect 20742 29034 20798 29036
rect 20742 28982 20744 29034
rect 20744 28982 20796 29034
rect 20796 28982 20798 29034
rect 20742 28980 20798 28982
rect 20846 29034 20902 29036
rect 20846 28982 20848 29034
rect 20848 28982 20900 29034
rect 20900 28982 20902 29034
rect 20846 28980 20902 28982
rect 20950 29034 21006 29036
rect 20950 28982 20952 29034
rect 20952 28982 21004 29034
rect 21004 28982 21006 29034
rect 20950 28980 21006 28982
rect 20860 28866 20916 28868
rect 20860 28814 20862 28866
rect 20862 28814 20914 28866
rect 20914 28814 20916 28866
rect 20860 28812 20916 28814
rect 19740 28588 19796 28644
rect 19964 28364 20020 28420
rect 20076 28140 20132 28196
rect 21308 29484 21364 29540
rect 21308 28812 21364 28868
rect 21308 28530 21364 28532
rect 21308 28478 21310 28530
rect 21310 28478 21362 28530
rect 21362 28478 21364 28530
rect 21308 28476 21364 28478
rect 21868 29820 21924 29876
rect 22540 29260 22596 29316
rect 22652 29372 22708 29428
rect 21756 28252 21812 28308
rect 20742 27466 20798 27468
rect 20742 27414 20744 27466
rect 20744 27414 20796 27466
rect 20796 27414 20798 27466
rect 20742 27412 20798 27414
rect 20846 27466 20902 27468
rect 20846 27414 20848 27466
rect 20848 27414 20900 27466
rect 20900 27414 20902 27466
rect 20846 27412 20902 27414
rect 20950 27466 21006 27468
rect 20950 27414 20952 27466
rect 20952 27414 21004 27466
rect 21004 27414 21006 27466
rect 20950 27412 21006 27414
rect 20300 26962 20356 26964
rect 20300 26910 20302 26962
rect 20302 26910 20354 26962
rect 20354 26910 20356 26962
rect 20300 26908 20356 26910
rect 20748 26796 20804 26852
rect 21644 27804 21700 27860
rect 22204 27298 22260 27300
rect 22204 27246 22206 27298
rect 22206 27246 22258 27298
rect 22258 27246 22260 27298
rect 22204 27244 22260 27246
rect 21532 26908 21588 26964
rect 21756 26908 21812 26964
rect 21084 26124 21140 26180
rect 20742 25898 20798 25900
rect 20742 25846 20744 25898
rect 20744 25846 20796 25898
rect 20796 25846 20798 25898
rect 20742 25844 20798 25846
rect 20846 25898 20902 25900
rect 20846 25846 20848 25898
rect 20848 25846 20900 25898
rect 20900 25846 20902 25898
rect 20846 25844 20902 25846
rect 20950 25898 21006 25900
rect 20950 25846 20952 25898
rect 20952 25846 21004 25898
rect 21004 25846 21006 25898
rect 20950 25844 21006 25846
rect 20076 25676 20132 25732
rect 22204 26796 22260 26852
rect 21980 26402 22036 26404
rect 21980 26350 21982 26402
rect 21982 26350 22034 26402
rect 22034 26350 22036 26402
rect 21980 26348 22036 26350
rect 19740 24946 19796 24948
rect 19740 24894 19742 24946
rect 19742 24894 19794 24946
rect 19794 24894 19796 24946
rect 19740 24892 19796 24894
rect 21084 25228 21140 25284
rect 20524 24834 20580 24836
rect 20524 24782 20526 24834
rect 20526 24782 20578 24834
rect 20578 24782 20580 24834
rect 20524 24780 20580 24782
rect 20742 24330 20798 24332
rect 20742 24278 20744 24330
rect 20744 24278 20796 24330
rect 20796 24278 20798 24330
rect 20742 24276 20798 24278
rect 20846 24330 20902 24332
rect 20846 24278 20848 24330
rect 20848 24278 20900 24330
rect 20900 24278 20902 24330
rect 20846 24276 20902 24278
rect 20950 24330 21006 24332
rect 20950 24278 20952 24330
rect 20952 24278 21004 24330
rect 21004 24278 21006 24330
rect 20950 24276 21006 24278
rect 20524 24108 20580 24164
rect 20300 23772 20356 23828
rect 21532 24668 21588 24724
rect 21196 24220 21252 24276
rect 20524 23212 20580 23268
rect 20860 23154 20916 23156
rect 20860 23102 20862 23154
rect 20862 23102 20914 23154
rect 20914 23102 20916 23154
rect 20860 23100 20916 23102
rect 20742 22762 20798 22764
rect 20742 22710 20744 22762
rect 20744 22710 20796 22762
rect 20796 22710 20798 22762
rect 20742 22708 20798 22710
rect 20846 22762 20902 22764
rect 20846 22710 20848 22762
rect 20848 22710 20900 22762
rect 20900 22710 20902 22762
rect 20846 22708 20902 22710
rect 20950 22762 21006 22764
rect 20950 22710 20952 22762
rect 20952 22710 21004 22762
rect 21004 22710 21006 22762
rect 20950 22708 21006 22710
rect 21644 24108 21700 24164
rect 21308 23826 21364 23828
rect 21308 23774 21310 23826
rect 21310 23774 21362 23826
rect 21362 23774 21364 23826
rect 21308 23772 21364 23774
rect 19964 22146 20020 22148
rect 19964 22094 19966 22146
rect 19966 22094 20018 22146
rect 20018 22094 20020 22146
rect 19964 22092 20020 22094
rect 20636 22092 20692 22148
rect 19516 21308 19572 21364
rect 20742 21194 20798 21196
rect 20742 21142 20744 21194
rect 20744 21142 20796 21194
rect 20796 21142 20798 21194
rect 20742 21140 20798 21142
rect 20846 21194 20902 21196
rect 20846 21142 20848 21194
rect 20848 21142 20900 21194
rect 20900 21142 20902 21194
rect 20846 21140 20902 21142
rect 20950 21194 21006 21196
rect 20950 21142 20952 21194
rect 20952 21142 21004 21194
rect 21004 21142 21006 21194
rect 20950 21140 21006 21142
rect 23548 30098 23604 30100
rect 23548 30046 23550 30098
rect 23550 30046 23602 30098
rect 23602 30046 23604 30098
rect 23548 30044 23604 30046
rect 24780 30098 24836 30100
rect 24780 30046 24782 30098
rect 24782 30046 24834 30098
rect 24834 30046 24836 30098
rect 24780 30044 24836 30046
rect 25228 30210 25284 30212
rect 25228 30158 25230 30210
rect 25230 30158 25282 30210
rect 25282 30158 25284 30210
rect 25228 30156 25284 30158
rect 24892 29932 24948 29988
rect 24648 29818 24704 29820
rect 24648 29766 24650 29818
rect 24650 29766 24702 29818
rect 24702 29766 24704 29818
rect 24648 29764 24704 29766
rect 24752 29818 24808 29820
rect 24752 29766 24754 29818
rect 24754 29766 24806 29818
rect 24806 29766 24808 29818
rect 24752 29764 24808 29766
rect 24856 29818 24912 29820
rect 24856 29766 24858 29818
rect 24858 29766 24910 29818
rect 24910 29766 24912 29818
rect 24856 29764 24912 29766
rect 23996 29650 24052 29652
rect 23996 29598 23998 29650
rect 23998 29598 24050 29650
rect 24050 29598 24052 29650
rect 23996 29596 24052 29598
rect 24556 29596 24612 29652
rect 22764 28588 22820 28644
rect 22876 29148 22932 29204
rect 23324 28924 23380 28980
rect 24332 29426 24388 29428
rect 24332 29374 24334 29426
rect 24334 29374 24386 29426
rect 24386 29374 24388 29426
rect 24332 29372 24388 29374
rect 23436 28588 23492 28644
rect 22988 26962 23044 26964
rect 22988 26910 22990 26962
rect 22990 26910 23042 26962
rect 23042 26910 23044 26962
rect 22988 26908 23044 26910
rect 23660 29148 23716 29204
rect 24332 28140 24388 28196
rect 24108 27970 24164 27972
rect 24108 27918 24110 27970
rect 24110 27918 24162 27970
rect 24162 27918 24164 27970
rect 24108 27916 24164 27918
rect 25340 29426 25396 29428
rect 25340 29374 25342 29426
rect 25342 29374 25394 29426
rect 25394 29374 25396 29426
rect 25340 29372 25396 29374
rect 24648 28250 24704 28252
rect 24648 28198 24650 28250
rect 24650 28198 24702 28250
rect 24702 28198 24704 28250
rect 24648 28196 24704 28198
rect 24752 28250 24808 28252
rect 24752 28198 24754 28250
rect 24754 28198 24806 28250
rect 24806 28198 24808 28250
rect 24752 28196 24808 28198
rect 24856 28250 24912 28252
rect 24856 28198 24858 28250
rect 24858 28198 24910 28250
rect 24910 28198 24912 28250
rect 24856 28196 24912 28198
rect 24444 27804 24500 27860
rect 25228 27692 25284 27748
rect 25004 27020 25060 27076
rect 22316 25228 22372 25284
rect 22204 24668 22260 24724
rect 22988 24162 23044 24164
rect 22988 24110 22990 24162
rect 22990 24110 23042 24162
rect 23042 24110 23044 24162
rect 22988 24108 23044 24110
rect 21980 21868 22036 21924
rect 21868 20914 21924 20916
rect 21868 20862 21870 20914
rect 21870 20862 21922 20914
rect 21922 20862 21924 20914
rect 21868 20860 21924 20862
rect 22204 21420 22260 21476
rect 19068 20802 19124 20804
rect 19068 20750 19070 20802
rect 19070 20750 19122 20802
rect 19122 20750 19124 20802
rect 19068 20748 19124 20750
rect 22316 22316 22372 22372
rect 22988 22652 23044 22708
rect 22204 20748 22260 20804
rect 18396 19906 18452 19908
rect 18396 19854 18398 19906
rect 18398 19854 18450 19906
rect 18450 19854 18452 19906
rect 18396 19852 18452 19854
rect 19404 20130 19460 20132
rect 19404 20078 19406 20130
rect 19406 20078 19458 20130
rect 19458 20078 19460 20130
rect 19404 20076 19460 20078
rect 20300 20076 20356 20132
rect 19068 19852 19124 19908
rect 18060 18508 18116 18564
rect 18396 18508 18452 18564
rect 18172 18060 18228 18116
rect 18508 17724 18564 17780
rect 17836 16716 17892 16772
rect 18732 17388 18788 17444
rect 18620 16044 18676 16100
rect 17724 15596 17780 15652
rect 18284 15484 18340 15540
rect 18172 15426 18228 15428
rect 18172 15374 18174 15426
rect 18174 15374 18226 15426
rect 18226 15374 18228 15426
rect 18172 15372 18228 15374
rect 17500 15202 17556 15204
rect 17500 15150 17502 15202
rect 17502 15150 17554 15202
rect 17554 15150 17556 15202
rect 17500 15148 17556 15150
rect 17388 14700 17444 14756
rect 16836 14138 16892 14140
rect 16836 14086 16838 14138
rect 16838 14086 16890 14138
rect 16890 14086 16892 14138
rect 16836 14084 16892 14086
rect 16940 14138 16996 14140
rect 16940 14086 16942 14138
rect 16942 14086 16994 14138
rect 16994 14086 16996 14138
rect 16940 14084 16996 14086
rect 17044 14138 17100 14140
rect 17044 14086 17046 14138
rect 17046 14086 17098 14138
rect 17098 14086 17100 14138
rect 17044 14084 17100 14086
rect 18060 13970 18116 13972
rect 18060 13918 18062 13970
rect 18062 13918 18114 13970
rect 18114 13918 18116 13970
rect 18060 13916 18116 13918
rect 18284 13580 18340 13636
rect 19180 19404 19236 19460
rect 18956 17164 19012 17220
rect 19404 17052 19460 17108
rect 21196 19906 21252 19908
rect 21196 19854 21198 19906
rect 21198 19854 21250 19906
rect 21250 19854 21252 19906
rect 21196 19852 21252 19854
rect 22204 20130 22260 20132
rect 22204 20078 22206 20130
rect 22206 20078 22258 20130
rect 22258 20078 22260 20130
rect 22204 20076 22260 20078
rect 21420 19852 21476 19908
rect 20742 19626 20798 19628
rect 20742 19574 20744 19626
rect 20744 19574 20796 19626
rect 20796 19574 20798 19626
rect 20742 19572 20798 19574
rect 20846 19626 20902 19628
rect 20846 19574 20848 19626
rect 20848 19574 20900 19626
rect 20900 19574 20902 19626
rect 20846 19572 20902 19574
rect 20950 19626 21006 19628
rect 20950 19574 20952 19626
rect 20952 19574 21004 19626
rect 21004 19574 21006 19626
rect 20950 19572 21006 19574
rect 19628 15932 19684 15988
rect 17724 13132 17780 13188
rect 17612 13020 17668 13076
rect 16836 12570 16892 12572
rect 16836 12518 16838 12570
rect 16838 12518 16890 12570
rect 16890 12518 16892 12570
rect 16836 12516 16892 12518
rect 16940 12570 16996 12572
rect 16940 12518 16942 12570
rect 16942 12518 16994 12570
rect 16994 12518 16996 12570
rect 16940 12516 16996 12518
rect 17044 12570 17100 12572
rect 17044 12518 17046 12570
rect 17046 12518 17098 12570
rect 17098 12518 17100 12570
rect 17044 12516 17100 12518
rect 17388 12290 17444 12292
rect 17388 12238 17390 12290
rect 17390 12238 17442 12290
rect 17442 12238 17444 12290
rect 17388 12236 17444 12238
rect 16492 12012 16548 12068
rect 15484 8988 15540 9044
rect 15036 7420 15092 7476
rect 14588 4620 14644 4676
rect 14700 6578 14756 6580
rect 14700 6526 14702 6578
rect 14702 6526 14754 6578
rect 14754 6526 14756 6578
rect 14700 6524 14756 6526
rect 15036 6524 15092 6580
rect 15372 7084 15428 7140
rect 15148 6466 15204 6468
rect 15148 6414 15150 6466
rect 15150 6414 15202 6466
rect 15202 6414 15204 6466
rect 15148 6412 15204 6414
rect 15148 5852 15204 5908
rect 16836 11002 16892 11004
rect 16836 10950 16838 11002
rect 16838 10950 16890 11002
rect 16890 10950 16892 11002
rect 16836 10948 16892 10950
rect 16940 11002 16996 11004
rect 16940 10950 16942 11002
rect 16942 10950 16994 11002
rect 16994 10950 16996 11002
rect 16940 10948 16996 10950
rect 17044 11002 17100 11004
rect 17044 10950 17046 11002
rect 17046 10950 17098 11002
rect 17098 10950 17100 11002
rect 17044 10948 17100 10950
rect 15820 8428 15876 8484
rect 15820 7644 15876 7700
rect 16268 9324 16324 9380
rect 16156 9154 16212 9156
rect 16156 9102 16158 9154
rect 16158 9102 16210 9154
rect 16210 9102 16212 9154
rect 16156 9100 16212 9102
rect 16836 9434 16892 9436
rect 16836 9382 16838 9434
rect 16838 9382 16890 9434
rect 16890 9382 16892 9434
rect 16836 9380 16892 9382
rect 16940 9434 16996 9436
rect 16940 9382 16942 9434
rect 16942 9382 16994 9434
rect 16994 9382 16996 9434
rect 16940 9380 16996 9382
rect 17044 9434 17100 9436
rect 17044 9382 17046 9434
rect 17046 9382 17098 9434
rect 17098 9382 17100 9434
rect 17044 9380 17100 9382
rect 16492 8876 16548 8932
rect 15932 7532 15988 7588
rect 16044 6636 16100 6692
rect 16044 6412 16100 6468
rect 16940 8092 16996 8148
rect 16836 7866 16892 7868
rect 16836 7814 16838 7866
rect 16838 7814 16890 7866
rect 16890 7814 16892 7866
rect 16836 7812 16892 7814
rect 16940 7866 16996 7868
rect 16940 7814 16942 7866
rect 16942 7814 16994 7866
rect 16994 7814 16996 7866
rect 16940 7812 16996 7814
rect 17044 7866 17100 7868
rect 17044 7814 17046 7866
rect 17046 7814 17098 7866
rect 17098 7814 17100 7866
rect 17044 7812 17100 7814
rect 16828 7698 16884 7700
rect 16828 7646 16830 7698
rect 16830 7646 16882 7698
rect 16882 7646 16884 7698
rect 16828 7644 16884 7646
rect 16268 7308 16324 7364
rect 16716 7196 16772 7252
rect 16156 5964 16212 6020
rect 16380 6524 16436 6580
rect 16836 6298 16892 6300
rect 16836 6246 16838 6298
rect 16838 6246 16890 6298
rect 16890 6246 16892 6298
rect 16836 6244 16892 6246
rect 16940 6298 16996 6300
rect 16940 6246 16942 6298
rect 16942 6246 16994 6298
rect 16994 6246 16996 6298
rect 16940 6244 16996 6246
rect 17044 6298 17100 6300
rect 17044 6246 17046 6298
rect 17046 6246 17098 6298
rect 17098 6246 17100 6298
rect 17044 6244 17100 6246
rect 19628 15372 19684 15428
rect 19180 14252 19236 14308
rect 20300 15932 20356 15988
rect 20748 19122 20804 19124
rect 20748 19070 20750 19122
rect 20750 19070 20802 19122
rect 20802 19070 20804 19122
rect 20748 19068 20804 19070
rect 21868 19234 21924 19236
rect 21868 19182 21870 19234
rect 21870 19182 21922 19234
rect 21922 19182 21924 19234
rect 21868 19180 21924 19182
rect 21196 18396 21252 18452
rect 20742 18058 20798 18060
rect 20742 18006 20744 18058
rect 20744 18006 20796 18058
rect 20796 18006 20798 18058
rect 20742 18004 20798 18006
rect 20846 18058 20902 18060
rect 20846 18006 20848 18058
rect 20848 18006 20900 18058
rect 20900 18006 20902 18058
rect 20846 18004 20902 18006
rect 20950 18058 21006 18060
rect 20950 18006 20952 18058
rect 20952 18006 21004 18058
rect 21004 18006 21006 18058
rect 20950 18004 21006 18006
rect 20748 17778 20804 17780
rect 20748 17726 20750 17778
rect 20750 17726 20802 17778
rect 20802 17726 20804 17778
rect 20748 17724 20804 17726
rect 22764 21474 22820 21476
rect 22764 21422 22766 21474
rect 22766 21422 22818 21474
rect 22818 21422 22820 21474
rect 22764 21420 22820 21422
rect 22652 21308 22708 21364
rect 22428 18450 22484 18452
rect 22428 18398 22430 18450
rect 22430 18398 22482 18450
rect 22482 18398 22484 18450
rect 22428 18396 22484 18398
rect 22092 18226 22148 18228
rect 22092 18174 22094 18226
rect 22094 18174 22146 18226
rect 22146 18174 22148 18226
rect 22092 18172 22148 18174
rect 23212 24722 23268 24724
rect 23212 24670 23214 24722
rect 23214 24670 23266 24722
rect 23266 24670 23268 24722
rect 23212 24668 23268 24670
rect 23100 21868 23156 21924
rect 24108 26796 24164 26852
rect 24648 26682 24704 26684
rect 24648 26630 24650 26682
rect 24650 26630 24702 26682
rect 24702 26630 24704 26682
rect 24648 26628 24704 26630
rect 24752 26682 24808 26684
rect 24752 26630 24754 26682
rect 24754 26630 24806 26682
rect 24806 26630 24808 26682
rect 24752 26628 24808 26630
rect 24856 26682 24912 26684
rect 24856 26630 24858 26682
rect 24858 26630 24910 26682
rect 24910 26630 24912 26682
rect 24856 26628 24912 26630
rect 24892 25730 24948 25732
rect 24892 25678 24894 25730
rect 24894 25678 24946 25730
rect 24946 25678 24948 25730
rect 24892 25676 24948 25678
rect 23660 24834 23716 24836
rect 23660 24782 23662 24834
rect 23662 24782 23714 24834
rect 23714 24782 23716 24834
rect 23660 24780 23716 24782
rect 23996 24834 24052 24836
rect 23996 24782 23998 24834
rect 23998 24782 24050 24834
rect 24050 24782 24052 24834
rect 23996 24780 24052 24782
rect 23996 24108 24052 24164
rect 23100 20242 23156 20244
rect 23100 20190 23102 20242
rect 23102 20190 23154 20242
rect 23154 20190 23156 20242
rect 23100 20188 23156 20190
rect 23548 21308 23604 21364
rect 23436 20188 23492 20244
rect 23548 19964 23604 20020
rect 23212 18284 23268 18340
rect 24648 25114 24704 25116
rect 24648 25062 24650 25114
rect 24650 25062 24702 25114
rect 24702 25062 24704 25114
rect 24648 25060 24704 25062
rect 24752 25114 24808 25116
rect 24752 25062 24754 25114
rect 24754 25062 24806 25114
rect 24806 25062 24808 25114
rect 24752 25060 24808 25062
rect 24856 25114 24912 25116
rect 24856 25062 24858 25114
rect 24858 25062 24910 25114
rect 24910 25062 24912 25114
rect 24856 25060 24912 25062
rect 24332 24834 24388 24836
rect 24332 24782 24334 24834
rect 24334 24782 24386 24834
rect 24386 24782 24388 24834
rect 24332 24780 24388 24782
rect 24648 23546 24704 23548
rect 24648 23494 24650 23546
rect 24650 23494 24702 23546
rect 24702 23494 24704 23546
rect 24648 23492 24704 23494
rect 24752 23546 24808 23548
rect 24752 23494 24754 23546
rect 24754 23494 24806 23546
rect 24806 23494 24808 23546
rect 24752 23492 24808 23494
rect 24856 23546 24912 23548
rect 24856 23494 24858 23546
rect 24858 23494 24910 23546
rect 24910 23494 24912 23546
rect 24856 23492 24912 23494
rect 24444 22988 24500 23044
rect 25900 29986 25956 29988
rect 25900 29934 25902 29986
rect 25902 29934 25954 29986
rect 25954 29934 25956 29986
rect 25900 29932 25956 29934
rect 26348 30156 26404 30212
rect 26236 29314 26292 29316
rect 26236 29262 26238 29314
rect 26238 29262 26290 29314
rect 26290 29262 26292 29314
rect 26236 29260 26292 29262
rect 25900 28812 25956 28868
rect 26236 28642 26292 28644
rect 26236 28590 26238 28642
rect 26238 28590 26290 28642
rect 26290 28590 26292 28642
rect 26236 28588 26292 28590
rect 26236 27746 26292 27748
rect 26236 27694 26238 27746
rect 26238 27694 26290 27746
rect 26290 27694 26292 27746
rect 26236 27692 26292 27694
rect 25788 26908 25844 26964
rect 24668 22370 24724 22372
rect 24668 22318 24670 22370
rect 24670 22318 24722 22370
rect 24722 22318 24724 22370
rect 24668 22316 24724 22318
rect 25788 23100 25844 23156
rect 25116 22316 25172 22372
rect 25676 22988 25732 23044
rect 24648 21978 24704 21980
rect 24648 21926 24650 21978
rect 24650 21926 24702 21978
rect 24702 21926 24704 21978
rect 24648 21924 24704 21926
rect 24752 21978 24808 21980
rect 24752 21926 24754 21978
rect 24754 21926 24806 21978
rect 24806 21926 24808 21978
rect 24752 21924 24808 21926
rect 24856 21978 24912 21980
rect 24856 21926 24858 21978
rect 24858 21926 24910 21978
rect 24910 21926 24912 21978
rect 24856 21924 24912 21926
rect 25116 21868 25172 21924
rect 24332 19740 24388 19796
rect 24648 20410 24704 20412
rect 24648 20358 24650 20410
rect 24650 20358 24702 20410
rect 24702 20358 24704 20410
rect 24648 20356 24704 20358
rect 24752 20410 24808 20412
rect 24752 20358 24754 20410
rect 24754 20358 24806 20410
rect 24806 20358 24808 20410
rect 24752 20356 24808 20358
rect 24856 20410 24912 20412
rect 24856 20358 24858 20410
rect 24858 20358 24910 20410
rect 24910 20358 24912 20410
rect 24856 20356 24912 20358
rect 25564 22146 25620 22148
rect 25564 22094 25566 22146
rect 25566 22094 25618 22146
rect 25618 22094 25620 22146
rect 25564 22092 25620 22094
rect 25788 20636 25844 20692
rect 25004 19964 25060 20020
rect 24892 19458 24948 19460
rect 24892 19406 24894 19458
rect 24894 19406 24946 19458
rect 24946 19406 24948 19458
rect 24892 19404 24948 19406
rect 25564 20018 25620 20020
rect 25564 19966 25566 20018
rect 25566 19966 25618 20018
rect 25618 19966 25620 20018
rect 25564 19964 25620 19966
rect 25564 19740 25620 19796
rect 24648 18842 24704 18844
rect 24648 18790 24650 18842
rect 24650 18790 24702 18842
rect 24702 18790 24704 18842
rect 24648 18788 24704 18790
rect 24752 18842 24808 18844
rect 24752 18790 24754 18842
rect 24754 18790 24806 18842
rect 24806 18790 24808 18842
rect 24752 18788 24808 18790
rect 24856 18842 24912 18844
rect 24856 18790 24858 18842
rect 24858 18790 24910 18842
rect 24910 18790 24912 18842
rect 24856 18788 24912 18790
rect 23324 18060 23380 18116
rect 20742 16490 20798 16492
rect 20742 16438 20744 16490
rect 20744 16438 20796 16490
rect 20796 16438 20798 16490
rect 20742 16436 20798 16438
rect 20846 16490 20902 16492
rect 20846 16438 20848 16490
rect 20848 16438 20900 16490
rect 20900 16438 20902 16490
rect 20846 16436 20902 16438
rect 20950 16490 21006 16492
rect 20950 16438 20952 16490
rect 20952 16438 21004 16490
rect 21004 16438 21006 16490
rect 20950 16436 21006 16438
rect 22540 17164 22596 17220
rect 21420 16098 21476 16100
rect 21420 16046 21422 16098
rect 21422 16046 21474 16098
rect 21474 16046 21476 16098
rect 21420 16044 21476 16046
rect 21308 15932 21364 15988
rect 20412 14924 20468 14980
rect 20742 14922 20798 14924
rect 20742 14870 20744 14922
rect 20744 14870 20796 14922
rect 20796 14870 20798 14922
rect 20742 14868 20798 14870
rect 20846 14922 20902 14924
rect 20846 14870 20848 14922
rect 20848 14870 20900 14922
rect 20900 14870 20902 14922
rect 20846 14868 20902 14870
rect 20950 14922 21006 14924
rect 20950 14870 20952 14922
rect 20952 14870 21004 14922
rect 21004 14870 21006 14922
rect 20950 14868 21006 14870
rect 20748 14418 20804 14420
rect 20748 14366 20750 14418
rect 20750 14366 20802 14418
rect 20802 14366 20804 14418
rect 20748 14364 20804 14366
rect 19068 13692 19124 13748
rect 18956 13580 19012 13636
rect 19292 13074 19348 13076
rect 19292 13022 19294 13074
rect 19294 13022 19346 13074
rect 19346 13022 19348 13074
rect 19292 13020 19348 13022
rect 20524 14252 20580 14308
rect 20748 13804 20804 13860
rect 20742 13354 20798 13356
rect 20742 13302 20744 13354
rect 20744 13302 20796 13354
rect 20796 13302 20798 13354
rect 20742 13300 20798 13302
rect 20846 13354 20902 13356
rect 20846 13302 20848 13354
rect 20848 13302 20900 13354
rect 20900 13302 20902 13354
rect 20846 13300 20902 13302
rect 20950 13354 21006 13356
rect 20950 13302 20952 13354
rect 20952 13302 21004 13354
rect 21004 13302 21006 13354
rect 20950 13300 21006 13302
rect 20188 12236 20244 12292
rect 18508 11676 18564 11732
rect 20742 11786 20798 11788
rect 20742 11734 20744 11786
rect 20744 11734 20796 11786
rect 20796 11734 20798 11786
rect 20742 11732 20798 11734
rect 20846 11786 20902 11788
rect 20846 11734 20848 11786
rect 20848 11734 20900 11786
rect 20900 11734 20902 11786
rect 20846 11732 20902 11734
rect 20950 11786 21006 11788
rect 20950 11734 20952 11786
rect 20952 11734 21004 11786
rect 21004 11734 21006 11786
rect 20950 11732 21006 11734
rect 19180 11452 19236 11508
rect 18172 11340 18228 11396
rect 18172 10610 18228 10612
rect 18172 10558 18174 10610
rect 18174 10558 18226 10610
rect 18226 10558 18228 10610
rect 18172 10556 18228 10558
rect 17724 9548 17780 9604
rect 19180 11170 19236 11172
rect 19180 11118 19182 11170
rect 19182 11118 19234 11170
rect 19234 11118 19236 11170
rect 19180 11116 19236 11118
rect 19068 10668 19124 10724
rect 19404 10610 19460 10612
rect 19404 10558 19406 10610
rect 19406 10558 19458 10610
rect 19458 10558 19460 10610
rect 19404 10556 19460 10558
rect 21420 13804 21476 13860
rect 21196 11394 21252 11396
rect 21196 11342 21198 11394
rect 21198 11342 21250 11394
rect 21250 11342 21252 11394
rect 21196 11340 21252 11342
rect 21084 11228 21140 11284
rect 20972 10722 21028 10724
rect 20972 10670 20974 10722
rect 20974 10670 21026 10722
rect 21026 10670 21028 10722
rect 20972 10668 21028 10670
rect 20524 10444 20580 10500
rect 20742 10218 20798 10220
rect 20742 10166 20744 10218
rect 20744 10166 20796 10218
rect 20796 10166 20798 10218
rect 20742 10164 20798 10166
rect 20846 10218 20902 10220
rect 20846 10166 20848 10218
rect 20848 10166 20900 10218
rect 20900 10166 20902 10218
rect 20846 10164 20902 10166
rect 20950 10218 21006 10220
rect 20950 10166 20952 10218
rect 20952 10166 21004 10218
rect 21004 10166 21006 10218
rect 20950 10164 21006 10166
rect 21868 14924 21924 14980
rect 21980 16044 22036 16100
rect 22988 16716 23044 16772
rect 23100 16604 23156 16660
rect 22652 16156 22708 16212
rect 22092 15090 22148 15092
rect 22092 15038 22094 15090
rect 22094 15038 22146 15090
rect 22146 15038 22148 15090
rect 22092 15036 22148 15038
rect 21756 14418 21812 14420
rect 21756 14366 21758 14418
rect 21758 14366 21810 14418
rect 21810 14366 21812 14418
rect 21756 14364 21812 14366
rect 23324 17666 23380 17668
rect 23324 17614 23326 17666
rect 23326 17614 23378 17666
rect 23378 17614 23380 17666
rect 23324 17612 23380 17614
rect 23660 17052 23716 17108
rect 23324 16994 23380 16996
rect 23324 16942 23326 16994
rect 23326 16942 23378 16994
rect 23378 16942 23380 16994
rect 23324 16940 23380 16942
rect 24332 17052 24388 17108
rect 23996 16940 24052 16996
rect 23212 15932 23268 15988
rect 23548 15820 23604 15876
rect 23996 16770 24052 16772
rect 23996 16718 23998 16770
rect 23998 16718 24050 16770
rect 24050 16718 24052 16770
rect 23996 16716 24052 16718
rect 24108 15874 24164 15876
rect 24108 15822 24110 15874
rect 24110 15822 24162 15874
rect 24162 15822 24164 15874
rect 24108 15820 24164 15822
rect 24332 15596 24388 15652
rect 24556 18060 24612 18116
rect 24648 17274 24704 17276
rect 24648 17222 24650 17274
rect 24650 17222 24702 17274
rect 24702 17222 24704 17274
rect 24648 17220 24704 17222
rect 24752 17274 24808 17276
rect 24752 17222 24754 17274
rect 24754 17222 24806 17274
rect 24806 17222 24808 17274
rect 24752 17220 24808 17222
rect 24856 17274 24912 17276
rect 24856 17222 24858 17274
rect 24858 17222 24910 17274
rect 24910 17222 24912 17274
rect 24856 17220 24912 17222
rect 25564 18284 25620 18340
rect 25452 18060 25508 18116
rect 25340 16882 25396 16884
rect 25340 16830 25342 16882
rect 25342 16830 25394 16882
rect 25394 16830 25396 16882
rect 25340 16828 25396 16830
rect 24668 16044 24724 16100
rect 24892 15986 24948 15988
rect 24892 15934 24894 15986
rect 24894 15934 24946 15986
rect 24946 15934 24948 15986
rect 24892 15932 24948 15934
rect 24648 15706 24704 15708
rect 24648 15654 24650 15706
rect 24650 15654 24702 15706
rect 24702 15654 24704 15706
rect 24648 15652 24704 15654
rect 24752 15706 24808 15708
rect 24752 15654 24754 15706
rect 24754 15654 24806 15706
rect 24806 15654 24808 15706
rect 24752 15652 24808 15654
rect 24856 15706 24912 15708
rect 24856 15654 24858 15706
rect 24858 15654 24910 15706
rect 24910 15654 24912 15706
rect 24856 15652 24912 15654
rect 24668 15426 24724 15428
rect 24668 15374 24670 15426
rect 24670 15374 24722 15426
rect 24722 15374 24724 15426
rect 24668 15372 24724 15374
rect 25788 17724 25844 17780
rect 25900 16940 25956 16996
rect 25564 16716 25620 16772
rect 25788 16716 25844 16772
rect 25676 15596 25732 15652
rect 24556 14588 24612 14644
rect 26796 30156 26852 30212
rect 26684 28924 26740 28980
rect 26908 29596 26964 29652
rect 27580 30156 27636 30212
rect 28554 30602 28610 30604
rect 28554 30550 28556 30602
rect 28556 30550 28608 30602
rect 28608 30550 28610 30602
rect 28554 30548 28610 30550
rect 28658 30602 28714 30604
rect 28658 30550 28660 30602
rect 28660 30550 28712 30602
rect 28712 30550 28714 30602
rect 28658 30548 28714 30550
rect 28762 30602 28818 30604
rect 28762 30550 28764 30602
rect 28764 30550 28816 30602
rect 28816 30550 28818 30602
rect 28762 30548 28818 30550
rect 28252 30044 28308 30100
rect 27356 29596 27412 29652
rect 27244 29538 27300 29540
rect 27244 29486 27246 29538
rect 27246 29486 27298 29538
rect 27298 29486 27300 29538
rect 27244 29484 27300 29486
rect 27468 29148 27524 29204
rect 28028 29596 28084 29652
rect 26236 26178 26292 26180
rect 26236 26126 26238 26178
rect 26238 26126 26290 26178
rect 26290 26126 26292 26178
rect 26236 26124 26292 26126
rect 26236 22652 26292 22708
rect 26572 25228 26628 25284
rect 26684 25564 26740 25620
rect 26572 24556 26628 24612
rect 26348 21756 26404 21812
rect 26348 20690 26404 20692
rect 26348 20638 26350 20690
rect 26350 20638 26402 20690
rect 26402 20638 26404 20690
rect 26348 20636 26404 20638
rect 26124 20578 26180 20580
rect 26124 20526 26126 20578
rect 26126 20526 26178 20578
rect 26178 20526 26180 20578
rect 26124 20524 26180 20526
rect 27244 27970 27300 27972
rect 27244 27918 27246 27970
rect 27246 27918 27298 27970
rect 27298 27918 27300 27970
rect 27244 27916 27300 27918
rect 27244 26402 27300 26404
rect 27244 26350 27246 26402
rect 27246 26350 27298 26402
rect 27298 26350 27300 26402
rect 27244 26348 27300 26350
rect 27132 25228 27188 25284
rect 27244 24220 27300 24276
rect 28554 29034 28610 29036
rect 28554 28982 28556 29034
rect 28556 28982 28608 29034
rect 28608 28982 28610 29034
rect 28554 28980 28610 28982
rect 28658 29034 28714 29036
rect 28658 28982 28660 29034
rect 28660 28982 28712 29034
rect 28712 28982 28714 29034
rect 28658 28980 28714 28982
rect 28762 29034 28818 29036
rect 28762 28982 28764 29034
rect 28764 28982 28816 29034
rect 28816 28982 28818 29034
rect 28762 28980 28818 28982
rect 28588 28476 28644 28532
rect 29036 28812 29092 28868
rect 28924 28028 28980 28084
rect 29036 28588 29092 28644
rect 27916 25228 27972 25284
rect 28554 27466 28610 27468
rect 28554 27414 28556 27466
rect 28556 27414 28608 27466
rect 28608 27414 28610 27466
rect 28554 27412 28610 27414
rect 28658 27466 28714 27468
rect 28658 27414 28660 27466
rect 28660 27414 28712 27466
rect 28712 27414 28714 27466
rect 28658 27412 28714 27414
rect 28762 27466 28818 27468
rect 28762 27414 28764 27466
rect 28764 27414 28816 27466
rect 28816 27414 28818 27466
rect 28762 27412 28818 27414
rect 28364 26908 28420 26964
rect 28812 26572 28868 26628
rect 28554 25898 28610 25900
rect 28554 25846 28556 25898
rect 28556 25846 28608 25898
rect 28608 25846 28610 25898
rect 28554 25844 28610 25846
rect 28658 25898 28714 25900
rect 28658 25846 28660 25898
rect 28660 25846 28712 25898
rect 28712 25846 28714 25898
rect 28658 25844 28714 25846
rect 28762 25898 28818 25900
rect 28762 25846 28764 25898
rect 28764 25846 28816 25898
rect 28816 25846 28818 25898
rect 28762 25844 28818 25846
rect 28252 24780 28308 24836
rect 27020 23324 27076 23380
rect 26684 23154 26740 23156
rect 26684 23102 26686 23154
rect 26686 23102 26738 23154
rect 26738 23102 26740 23154
rect 26684 23100 26740 23102
rect 26684 20914 26740 20916
rect 26684 20862 26686 20914
rect 26686 20862 26738 20914
rect 26738 20862 26740 20914
rect 26684 20860 26740 20862
rect 26684 18562 26740 18564
rect 26684 18510 26686 18562
rect 26686 18510 26738 18562
rect 26738 18510 26740 18562
rect 26684 18508 26740 18510
rect 26124 18284 26180 18340
rect 26460 18284 26516 18340
rect 26572 18060 26628 18116
rect 26348 17554 26404 17556
rect 26348 17502 26350 17554
rect 26350 17502 26402 17554
rect 26402 17502 26404 17554
rect 26348 17500 26404 17502
rect 26124 17052 26180 17108
rect 26012 15372 26068 15428
rect 27132 18284 27188 18340
rect 27132 17612 27188 17668
rect 26908 17052 26964 17108
rect 26908 16044 26964 16100
rect 24648 14138 24704 14140
rect 24648 14086 24650 14138
rect 24650 14086 24702 14138
rect 24702 14086 24704 14138
rect 24648 14084 24704 14086
rect 24752 14138 24808 14140
rect 24752 14086 24754 14138
rect 24754 14086 24806 14138
rect 24806 14086 24808 14138
rect 24752 14084 24808 14086
rect 24856 14138 24912 14140
rect 24856 14086 24858 14138
rect 24858 14086 24910 14138
rect 24910 14086 24912 14138
rect 24856 14084 24912 14086
rect 22876 13692 22932 13748
rect 22540 13634 22596 13636
rect 22540 13582 22542 13634
rect 22542 13582 22594 13634
rect 22594 13582 22596 13634
rect 22540 13580 22596 13582
rect 21868 13132 21924 13188
rect 21756 11676 21812 11732
rect 21644 10668 21700 10724
rect 21532 9996 21588 10052
rect 21868 10498 21924 10500
rect 21868 10446 21870 10498
rect 21870 10446 21922 10498
rect 21922 10446 21924 10498
rect 21868 10444 21924 10446
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 25676 13580 25732 13636
rect 26348 13580 26404 13636
rect 26796 14924 26852 14980
rect 32284 31612 32340 31668
rect 29932 30940 29988 30996
rect 29148 28476 29204 28532
rect 29036 25228 29092 25284
rect 29148 28252 29204 28308
rect 28364 24610 28420 24612
rect 28364 24558 28366 24610
rect 28366 24558 28418 24610
rect 28418 24558 28420 24610
rect 28364 24556 28420 24558
rect 28554 24330 28610 24332
rect 28554 24278 28556 24330
rect 28556 24278 28608 24330
rect 28608 24278 28610 24330
rect 28554 24276 28610 24278
rect 28658 24330 28714 24332
rect 28658 24278 28660 24330
rect 28660 24278 28712 24330
rect 28712 24278 28714 24330
rect 28658 24276 28714 24278
rect 28762 24330 28818 24332
rect 28762 24278 28764 24330
rect 28764 24278 28816 24330
rect 28816 24278 28818 24330
rect 28762 24276 28818 24278
rect 28554 22762 28610 22764
rect 28554 22710 28556 22762
rect 28556 22710 28608 22762
rect 28608 22710 28610 22762
rect 28554 22708 28610 22710
rect 28658 22762 28714 22764
rect 28658 22710 28660 22762
rect 28660 22710 28712 22762
rect 28712 22710 28714 22762
rect 28658 22708 28714 22710
rect 28762 22762 28818 22764
rect 28762 22710 28764 22762
rect 28764 22710 28816 22762
rect 28816 22710 28818 22762
rect 28762 22708 28818 22710
rect 28140 22428 28196 22484
rect 28252 21420 28308 21476
rect 28554 21194 28610 21196
rect 28554 21142 28556 21194
rect 28556 21142 28608 21194
rect 28608 21142 28610 21194
rect 28554 21140 28610 21142
rect 28658 21194 28714 21196
rect 28658 21142 28660 21194
rect 28660 21142 28712 21194
rect 28712 21142 28714 21194
rect 28658 21140 28714 21142
rect 28762 21194 28818 21196
rect 28762 21142 28764 21194
rect 28764 21142 28816 21194
rect 28816 21142 28818 21194
rect 28762 21140 28818 21142
rect 29372 27580 29428 27636
rect 29708 26908 29764 26964
rect 29260 25788 29316 25844
rect 32060 30268 32116 30324
rect 30268 27244 30324 27300
rect 30940 29260 30996 29316
rect 29708 26124 29764 26180
rect 29148 20636 29204 20692
rect 28476 20188 28532 20244
rect 30044 26572 30100 26628
rect 30716 25788 30772 25844
rect 30156 25618 30212 25620
rect 30156 25566 30158 25618
rect 30158 25566 30210 25618
rect 30210 25566 30212 25618
rect 30156 25564 30212 25566
rect 30156 22482 30212 22484
rect 30156 22430 30158 22482
rect 30158 22430 30210 22482
rect 30210 22430 30212 22482
rect 30156 22428 30212 22430
rect 30044 21756 30100 21812
rect 30044 21474 30100 21476
rect 30044 21422 30046 21474
rect 30046 21422 30098 21474
rect 30098 21422 30100 21474
rect 30044 21420 30100 21422
rect 27356 19516 27412 19572
rect 28554 19626 28610 19628
rect 28554 19574 28556 19626
rect 28556 19574 28608 19626
rect 28608 19574 28610 19626
rect 28554 19572 28610 19574
rect 28658 19626 28714 19628
rect 28658 19574 28660 19626
rect 28660 19574 28712 19626
rect 28712 19574 28714 19626
rect 28658 19572 28714 19574
rect 28762 19626 28818 19628
rect 28762 19574 28764 19626
rect 28764 19574 28816 19626
rect 28816 19574 28818 19626
rect 28762 19572 28818 19574
rect 28700 19234 28756 19236
rect 28700 19182 28702 19234
rect 28702 19182 28754 19234
rect 28754 19182 28756 19234
rect 28700 19180 28756 19182
rect 29484 19180 29540 19236
rect 28140 18674 28196 18676
rect 28140 18622 28142 18674
rect 28142 18622 28194 18674
rect 28194 18622 28196 18674
rect 28140 18620 28196 18622
rect 29148 18396 29204 18452
rect 27580 18338 27636 18340
rect 27580 18286 27582 18338
rect 27582 18286 27634 18338
rect 27634 18286 27636 18338
rect 27580 18284 27636 18286
rect 28554 18058 28610 18060
rect 28554 18006 28556 18058
rect 28556 18006 28608 18058
rect 28608 18006 28610 18058
rect 28554 18004 28610 18006
rect 28658 18058 28714 18060
rect 28658 18006 28660 18058
rect 28660 18006 28712 18058
rect 28712 18006 28714 18058
rect 28658 18004 28714 18006
rect 28762 18058 28818 18060
rect 28762 18006 28764 18058
rect 28764 18006 28816 18058
rect 28816 18006 28818 18058
rect 28762 18004 28818 18006
rect 27356 17666 27412 17668
rect 27356 17614 27358 17666
rect 27358 17614 27410 17666
rect 27410 17614 27412 17666
rect 27356 17612 27412 17614
rect 28028 17106 28084 17108
rect 28028 17054 28030 17106
rect 28030 17054 28082 17106
rect 28082 17054 28084 17106
rect 28028 17052 28084 17054
rect 27244 14364 27300 14420
rect 27916 15036 27972 15092
rect 28140 14028 28196 14084
rect 23100 11116 23156 11172
rect 18956 9772 19012 9828
rect 19404 9826 19460 9828
rect 19404 9774 19406 9826
rect 19406 9774 19458 9826
rect 19458 9774 19460 9826
rect 19404 9772 19460 9774
rect 20748 9826 20804 9828
rect 20748 9774 20750 9826
rect 20750 9774 20802 9826
rect 20802 9774 20804 9826
rect 20748 9772 20804 9774
rect 21532 9826 21588 9828
rect 21532 9774 21534 9826
rect 21534 9774 21586 9826
rect 21586 9774 21588 9826
rect 21532 9772 21588 9774
rect 19180 9602 19236 9604
rect 19180 9550 19182 9602
rect 19182 9550 19234 9602
rect 19234 9550 19236 9602
rect 19180 9548 19236 9550
rect 18956 9042 19012 9044
rect 18956 8990 18958 9042
rect 18958 8990 19010 9042
rect 19010 8990 19012 9042
rect 18956 8988 19012 8990
rect 19180 8988 19236 9044
rect 21532 9212 21588 9268
rect 21644 9548 21700 9604
rect 21420 8988 21476 9044
rect 17500 8204 17556 8260
rect 17500 7420 17556 7476
rect 17164 5180 17220 5236
rect 14700 4284 14756 4340
rect 17500 6412 17556 6468
rect 17276 5068 17332 5124
rect 17388 5964 17444 6020
rect 16604 4956 16660 5012
rect 15484 4844 15540 4900
rect 16268 4450 16324 4452
rect 16268 4398 16270 4450
rect 16270 4398 16322 4450
rect 16322 4398 16324 4450
rect 16268 4396 16324 4398
rect 17164 4956 17220 5012
rect 16836 4730 16892 4732
rect 16836 4678 16838 4730
rect 16838 4678 16890 4730
rect 16890 4678 16892 4730
rect 16836 4676 16892 4678
rect 16940 4730 16996 4732
rect 16940 4678 16942 4730
rect 16942 4678 16994 4730
rect 16994 4678 16996 4730
rect 16940 4676 16996 4678
rect 17044 4730 17100 4732
rect 17044 4678 17046 4730
rect 17046 4678 17098 4730
rect 17098 4678 17100 4730
rect 17044 4676 17100 4678
rect 15148 4172 15204 4228
rect 14812 4060 14868 4116
rect 18396 8204 18452 8260
rect 19292 8764 19348 8820
rect 20742 8650 20798 8652
rect 20742 8598 20744 8650
rect 20744 8598 20796 8650
rect 20796 8598 20798 8650
rect 20742 8596 20798 8598
rect 20846 8650 20902 8652
rect 20846 8598 20848 8650
rect 20848 8598 20900 8650
rect 20900 8598 20902 8650
rect 20846 8596 20902 8598
rect 20950 8650 21006 8652
rect 20950 8598 20952 8650
rect 20952 8598 21004 8650
rect 21004 8598 21006 8650
rect 20950 8596 21006 8598
rect 19404 8092 19460 8148
rect 17948 7698 18004 7700
rect 17948 7646 17950 7698
rect 17950 7646 18002 7698
rect 18002 7646 18004 7698
rect 17948 7644 18004 7646
rect 17836 6748 17892 6804
rect 17836 6300 17892 6356
rect 17724 5068 17780 5124
rect 18732 7420 18788 7476
rect 18396 7362 18452 7364
rect 18396 7310 18398 7362
rect 18398 7310 18450 7362
rect 18450 7310 18452 7362
rect 18396 7308 18452 7310
rect 18172 6524 18228 6580
rect 18060 5740 18116 5796
rect 18284 6466 18340 6468
rect 18284 6414 18286 6466
rect 18286 6414 18338 6466
rect 18338 6414 18340 6466
rect 18284 6412 18340 6414
rect 18620 6300 18676 6356
rect 17724 3666 17780 3668
rect 17724 3614 17726 3666
rect 17726 3614 17778 3666
rect 17778 3614 17780 3666
rect 17724 3612 17780 3614
rect 18508 4284 18564 4340
rect 18396 4226 18452 4228
rect 18396 4174 18398 4226
rect 18398 4174 18450 4226
rect 18450 4174 18452 4226
rect 18396 4172 18452 4174
rect 19180 6802 19236 6804
rect 19180 6750 19182 6802
rect 19182 6750 19234 6802
rect 19234 6750 19236 6802
rect 19180 6748 19236 6750
rect 18844 6690 18900 6692
rect 18844 6638 18846 6690
rect 18846 6638 18898 6690
rect 18898 6638 18900 6690
rect 18844 6636 18900 6638
rect 21196 8258 21252 8260
rect 21196 8206 21198 8258
rect 21198 8206 21250 8258
rect 21250 8206 21252 8258
rect 21196 8204 21252 8206
rect 19516 6636 19572 6692
rect 18620 3724 18676 3780
rect 18956 4508 19012 4564
rect 18396 3612 18452 3668
rect 16828 3500 16884 3556
rect 14252 3388 14308 3444
rect 15820 3442 15876 3444
rect 15820 3390 15822 3442
rect 15822 3390 15874 3442
rect 15874 3390 15876 3442
rect 15820 3388 15876 3390
rect 19404 4450 19460 4452
rect 19404 4398 19406 4450
rect 19406 4398 19458 4450
rect 19458 4398 19460 4450
rect 19404 4396 19460 4398
rect 20524 7980 20580 8036
rect 20076 7250 20132 7252
rect 20076 7198 20078 7250
rect 20078 7198 20130 7250
rect 20130 7198 20132 7250
rect 20076 7196 20132 7198
rect 20300 6636 20356 6692
rect 20188 6578 20244 6580
rect 20188 6526 20190 6578
rect 20190 6526 20242 6578
rect 20242 6526 20244 6578
rect 20188 6524 20244 6526
rect 19852 5122 19908 5124
rect 19852 5070 19854 5122
rect 19854 5070 19906 5122
rect 19906 5070 19908 5122
rect 19852 5068 19908 5070
rect 20300 5292 20356 5348
rect 20412 5180 20468 5236
rect 20188 4172 20244 4228
rect 20300 4284 20356 4340
rect 19628 3948 19684 4004
rect 19852 3554 19908 3556
rect 19852 3502 19854 3554
rect 19854 3502 19906 3554
rect 19906 3502 19908 3554
rect 19852 3500 19908 3502
rect 20748 7644 20804 7700
rect 20742 7082 20798 7084
rect 20742 7030 20744 7082
rect 20744 7030 20796 7082
rect 20796 7030 20798 7082
rect 20742 7028 20798 7030
rect 20846 7082 20902 7084
rect 20846 7030 20848 7082
rect 20848 7030 20900 7082
rect 20900 7030 20902 7082
rect 20846 7028 20902 7030
rect 20950 7082 21006 7084
rect 20950 7030 20952 7082
rect 20952 7030 21004 7082
rect 21004 7030 21006 7082
rect 20950 7028 21006 7030
rect 20972 6018 21028 6020
rect 20972 5966 20974 6018
rect 20974 5966 21026 6018
rect 21026 5966 21028 6018
rect 20972 5964 21028 5966
rect 20742 5514 20798 5516
rect 20742 5462 20744 5514
rect 20744 5462 20796 5514
rect 20796 5462 20798 5514
rect 20742 5460 20798 5462
rect 20846 5514 20902 5516
rect 20846 5462 20848 5514
rect 20848 5462 20900 5514
rect 20900 5462 20902 5514
rect 20846 5460 20902 5462
rect 20950 5514 21006 5516
rect 20950 5462 20952 5514
rect 20952 5462 21004 5514
rect 21004 5462 21006 5514
rect 20950 5460 21006 5462
rect 21532 6524 21588 6580
rect 22316 9266 22372 9268
rect 22316 9214 22318 9266
rect 22318 9214 22370 9266
rect 22370 9214 22372 9266
rect 22316 9212 22372 9214
rect 21980 7308 22036 7364
rect 21980 6748 22036 6804
rect 22316 6524 22372 6580
rect 21308 5628 21364 5684
rect 21196 5292 21252 5348
rect 20748 4898 20804 4900
rect 20748 4846 20750 4898
rect 20750 4846 20802 4898
rect 20802 4846 20804 4898
rect 20748 4844 20804 4846
rect 21756 5404 21812 5460
rect 21980 5346 22036 5348
rect 21980 5294 21982 5346
rect 21982 5294 22034 5346
rect 22034 5294 22036 5346
rect 21980 5292 22036 5294
rect 22092 5122 22148 5124
rect 22092 5070 22094 5122
rect 22094 5070 22146 5122
rect 22146 5070 22148 5122
rect 22092 5068 22148 5070
rect 21308 4172 21364 4228
rect 22316 6018 22372 6020
rect 22316 5966 22318 6018
rect 22318 5966 22370 6018
rect 22370 5966 22372 6018
rect 22316 5964 22372 5966
rect 22428 5628 22484 5684
rect 22876 9266 22932 9268
rect 22876 9214 22878 9266
rect 22878 9214 22930 9266
rect 22930 9214 22932 9266
rect 22876 9212 22932 9214
rect 24648 12570 24704 12572
rect 24648 12518 24650 12570
rect 24650 12518 24702 12570
rect 24702 12518 24704 12570
rect 24648 12516 24704 12518
rect 24752 12570 24808 12572
rect 24752 12518 24754 12570
rect 24754 12518 24806 12570
rect 24806 12518 24808 12570
rect 24752 12516 24808 12518
rect 24856 12570 24912 12572
rect 24856 12518 24858 12570
rect 24858 12518 24910 12570
rect 24910 12518 24912 12570
rect 24856 12516 24912 12518
rect 26460 13132 26516 13188
rect 27804 13356 27860 13412
rect 23884 12290 23940 12292
rect 23884 12238 23886 12290
rect 23886 12238 23938 12290
rect 23938 12238 23940 12290
rect 23884 12236 23940 12238
rect 27804 12124 27860 12180
rect 25228 11452 25284 11508
rect 26348 11452 26404 11508
rect 25116 11228 25172 11284
rect 24108 11170 24164 11172
rect 24108 11118 24110 11170
rect 24110 11118 24162 11170
rect 24162 11118 24164 11170
rect 24108 11116 24164 11118
rect 24648 11002 24704 11004
rect 24648 10950 24650 11002
rect 24650 10950 24702 11002
rect 24702 10950 24704 11002
rect 24648 10948 24704 10950
rect 24752 11002 24808 11004
rect 24752 10950 24754 11002
rect 24754 10950 24806 11002
rect 24806 10950 24808 11002
rect 24752 10948 24808 10950
rect 24856 11002 24912 11004
rect 24856 10950 24858 11002
rect 24858 10950 24910 11002
rect 24910 10950 24912 11002
rect 24856 10948 24912 10950
rect 23884 10722 23940 10724
rect 23884 10670 23886 10722
rect 23886 10670 23938 10722
rect 23938 10670 23940 10722
rect 23884 10668 23940 10670
rect 24444 10556 24500 10612
rect 23212 8930 23268 8932
rect 23212 8878 23214 8930
rect 23214 8878 23266 8930
rect 23266 8878 23268 8930
rect 23212 8876 23268 8878
rect 22988 8652 23044 8708
rect 23548 8204 23604 8260
rect 23100 6802 23156 6804
rect 23100 6750 23102 6802
rect 23102 6750 23154 6802
rect 23154 6750 23156 6802
rect 23100 6748 23156 6750
rect 24220 9154 24276 9156
rect 24220 9102 24222 9154
rect 24222 9102 24274 9154
rect 24274 9102 24276 9154
rect 24220 9100 24276 9102
rect 24332 8764 24388 8820
rect 25004 9660 25060 9716
rect 25676 9884 25732 9940
rect 25564 9548 25620 9604
rect 25788 9548 25844 9604
rect 24648 9434 24704 9436
rect 24648 9382 24650 9434
rect 24650 9382 24702 9434
rect 24702 9382 24704 9434
rect 24648 9380 24704 9382
rect 24752 9434 24808 9436
rect 24752 9382 24754 9434
rect 24754 9382 24806 9434
rect 24806 9382 24808 9434
rect 24752 9380 24808 9382
rect 24856 9434 24912 9436
rect 24856 9382 24858 9434
rect 24858 9382 24910 9434
rect 24910 9382 24912 9434
rect 24856 9380 24912 9382
rect 25228 9212 25284 9268
rect 25340 8818 25396 8820
rect 25340 8766 25342 8818
rect 25342 8766 25394 8818
rect 25394 8766 25396 8818
rect 25340 8764 25396 8766
rect 24648 7866 24704 7868
rect 24648 7814 24650 7866
rect 24650 7814 24702 7866
rect 24702 7814 24704 7866
rect 24648 7812 24704 7814
rect 24752 7866 24808 7868
rect 24752 7814 24754 7866
rect 24754 7814 24806 7866
rect 24806 7814 24808 7866
rect 24752 7812 24808 7814
rect 24856 7866 24912 7868
rect 24856 7814 24858 7866
rect 24858 7814 24910 7866
rect 24910 7814 24912 7866
rect 24856 7812 24912 7814
rect 24332 7474 24388 7476
rect 24332 7422 24334 7474
rect 24334 7422 24386 7474
rect 24386 7422 24388 7474
rect 24332 7420 24388 7422
rect 23996 6748 24052 6804
rect 24108 7308 24164 7364
rect 24648 6298 24704 6300
rect 24648 6246 24650 6298
rect 24650 6246 24702 6298
rect 24702 6246 24704 6298
rect 24648 6244 24704 6246
rect 24752 6298 24808 6300
rect 24752 6246 24754 6298
rect 24754 6246 24806 6298
rect 24806 6246 24808 6298
rect 24752 6244 24808 6246
rect 24856 6298 24912 6300
rect 24856 6246 24858 6298
rect 24858 6246 24910 6298
rect 24910 6246 24912 6298
rect 24856 6244 24912 6246
rect 26796 11004 26852 11060
rect 28252 10780 28308 10836
rect 28588 17388 28644 17444
rect 29260 17666 29316 17668
rect 29260 17614 29262 17666
rect 29262 17614 29314 17666
rect 29314 17614 29316 17666
rect 29260 17612 29316 17614
rect 29596 17388 29652 17444
rect 29260 16828 29316 16884
rect 28554 16490 28610 16492
rect 28554 16438 28556 16490
rect 28556 16438 28608 16490
rect 28608 16438 28610 16490
rect 28554 16436 28610 16438
rect 28658 16490 28714 16492
rect 28658 16438 28660 16490
rect 28660 16438 28712 16490
rect 28712 16438 28714 16490
rect 28658 16436 28714 16438
rect 28762 16490 28818 16492
rect 28762 16438 28764 16490
rect 28764 16438 28816 16490
rect 28816 16438 28818 16490
rect 28762 16436 28818 16438
rect 28924 16380 28980 16436
rect 29372 16380 29428 16436
rect 28554 14922 28610 14924
rect 28554 14870 28556 14922
rect 28556 14870 28608 14922
rect 28608 14870 28610 14922
rect 28554 14868 28610 14870
rect 28658 14922 28714 14924
rect 28658 14870 28660 14922
rect 28660 14870 28712 14922
rect 28712 14870 28714 14922
rect 28658 14868 28714 14870
rect 28762 14922 28818 14924
rect 28762 14870 28764 14922
rect 28764 14870 28816 14922
rect 28816 14870 28818 14922
rect 28762 14868 28818 14870
rect 29372 14140 29428 14196
rect 28554 13354 28610 13356
rect 28554 13302 28556 13354
rect 28556 13302 28608 13354
rect 28608 13302 28610 13354
rect 28554 13300 28610 13302
rect 28658 13354 28714 13356
rect 28658 13302 28660 13354
rect 28660 13302 28712 13354
rect 28712 13302 28714 13354
rect 28658 13300 28714 13302
rect 28762 13354 28818 13356
rect 28762 13302 28764 13354
rect 28764 13302 28816 13354
rect 28816 13302 28818 13354
rect 28762 13300 28818 13302
rect 29596 14252 29652 14308
rect 29820 14306 29876 14308
rect 29820 14254 29822 14306
rect 29822 14254 29874 14306
rect 29874 14254 29876 14306
rect 29820 14252 29876 14254
rect 29148 12178 29204 12180
rect 29148 12126 29150 12178
rect 29150 12126 29202 12178
rect 29202 12126 29204 12178
rect 29148 12124 29204 12126
rect 28554 11786 28610 11788
rect 28554 11734 28556 11786
rect 28556 11734 28608 11786
rect 28608 11734 28610 11786
rect 28554 11732 28610 11734
rect 28658 11786 28714 11788
rect 28658 11734 28660 11786
rect 28660 11734 28712 11786
rect 28712 11734 28714 11786
rect 28658 11732 28714 11734
rect 28762 11786 28818 11788
rect 28762 11734 28764 11786
rect 28764 11734 28816 11786
rect 28816 11734 28818 11786
rect 28762 11732 28818 11734
rect 29820 12124 29876 12180
rect 29260 11506 29316 11508
rect 29260 11454 29262 11506
rect 29262 11454 29314 11506
rect 29314 11454 29316 11506
rect 29260 11452 29316 11454
rect 29820 11452 29876 11508
rect 28554 10218 28610 10220
rect 28554 10166 28556 10218
rect 28556 10166 28608 10218
rect 28608 10166 28610 10218
rect 28554 10164 28610 10166
rect 28658 10218 28714 10220
rect 28658 10166 28660 10218
rect 28660 10166 28712 10218
rect 28712 10166 28714 10218
rect 28658 10164 28714 10166
rect 28762 10218 28818 10220
rect 28762 10166 28764 10218
rect 28764 10166 28816 10218
rect 28816 10166 28818 10218
rect 28762 10164 28818 10166
rect 28364 9996 28420 10052
rect 26348 8652 26404 8708
rect 27468 9602 27524 9604
rect 27468 9550 27470 9602
rect 27470 9550 27522 9602
rect 27522 9550 27524 9602
rect 27468 9548 27524 9550
rect 27356 9436 27412 9492
rect 28588 9436 28644 9492
rect 27356 8652 27412 8708
rect 28028 8428 28084 8484
rect 28140 8764 28196 8820
rect 27132 8092 27188 8148
rect 25900 7980 25956 8036
rect 26236 7362 26292 7364
rect 26236 7310 26238 7362
rect 26238 7310 26290 7362
rect 26290 7310 26292 7362
rect 26236 7308 26292 7310
rect 25116 6524 25172 6580
rect 25004 5964 25060 6020
rect 23772 5346 23828 5348
rect 23772 5294 23774 5346
rect 23774 5294 23826 5346
rect 23826 5294 23828 5346
rect 23772 5292 23828 5294
rect 24332 5234 24388 5236
rect 24332 5182 24334 5234
rect 24334 5182 24386 5234
rect 24386 5182 24388 5234
rect 24332 5180 24388 5182
rect 22540 5068 22596 5124
rect 22764 4844 22820 4900
rect 24668 5122 24724 5124
rect 24668 5070 24670 5122
rect 24670 5070 24722 5122
rect 24722 5070 24724 5122
rect 24668 5068 24724 5070
rect 25340 4844 25396 4900
rect 24648 4730 24704 4732
rect 24648 4678 24650 4730
rect 24650 4678 24702 4730
rect 24702 4678 24704 4730
rect 24648 4676 24704 4678
rect 24752 4730 24808 4732
rect 24752 4678 24754 4730
rect 24754 4678 24806 4730
rect 24806 4678 24808 4730
rect 24752 4676 24808 4678
rect 24856 4730 24912 4732
rect 24856 4678 24858 4730
rect 24858 4678 24910 4730
rect 24910 4678 24912 4730
rect 24856 4676 24912 4678
rect 23548 4338 23604 4340
rect 23548 4286 23550 4338
rect 23550 4286 23602 4338
rect 23602 4286 23604 4338
rect 23548 4284 23604 4286
rect 20742 3946 20798 3948
rect 20742 3894 20744 3946
rect 20744 3894 20796 3946
rect 20796 3894 20798 3946
rect 20742 3892 20798 3894
rect 20846 3946 20902 3948
rect 20846 3894 20848 3946
rect 20848 3894 20900 3946
rect 20900 3894 20902 3946
rect 20846 3892 20902 3894
rect 20950 3946 21006 3948
rect 20950 3894 20952 3946
rect 20952 3894 21004 3946
rect 21004 3894 21006 3946
rect 20950 3892 21006 3894
rect 22204 3554 22260 3556
rect 22204 3502 22206 3554
rect 22206 3502 22258 3554
rect 22258 3502 22260 3554
rect 22204 3500 22260 3502
rect 24108 4172 24164 4228
rect 23436 3836 23492 3892
rect 24668 4226 24724 4228
rect 24668 4174 24670 4226
rect 24670 4174 24722 4226
rect 24722 4174 24724 4226
rect 24668 4172 24724 4174
rect 24220 4114 24276 4116
rect 24220 4062 24222 4114
rect 24222 4062 24274 4114
rect 24274 4062 24276 4114
rect 24220 4060 24276 4062
rect 25004 3612 25060 3668
rect 24220 3500 24276 3556
rect 22428 3442 22484 3444
rect 22428 3390 22430 3442
rect 22430 3390 22482 3442
rect 22482 3390 22484 3442
rect 22428 3388 22484 3390
rect 12348 3330 12404 3332
rect 12348 3278 12350 3330
rect 12350 3278 12402 3330
rect 12402 3278 12404 3330
rect 12348 3276 12404 3278
rect 22876 3276 22932 3332
rect 16836 3162 16892 3164
rect 16836 3110 16838 3162
rect 16838 3110 16890 3162
rect 16890 3110 16892 3162
rect 16836 3108 16892 3110
rect 16940 3162 16996 3164
rect 16940 3110 16942 3162
rect 16942 3110 16994 3162
rect 16994 3110 16996 3162
rect 16940 3108 16996 3110
rect 17044 3162 17100 3164
rect 17044 3110 17046 3162
rect 17046 3110 17098 3162
rect 17098 3110 17100 3162
rect 17044 3108 17100 3110
rect 12236 2716 12292 2772
rect 24556 3330 24612 3332
rect 24556 3278 24558 3330
rect 24558 3278 24610 3330
rect 24610 3278 24612 3330
rect 24556 3276 24612 3278
rect 24648 3162 24704 3164
rect 24648 3110 24650 3162
rect 24650 3110 24702 3162
rect 24702 3110 24704 3162
rect 24648 3108 24704 3110
rect 24752 3162 24808 3164
rect 24752 3110 24754 3162
rect 24754 3110 24806 3162
rect 24806 3110 24808 3162
rect 24752 3108 24808 3110
rect 24856 3162 24912 3164
rect 24856 3110 24858 3162
rect 24858 3110 24910 3162
rect 24910 3110 24912 3162
rect 24856 3108 24912 3110
rect 25116 3554 25172 3556
rect 25116 3502 25118 3554
rect 25118 3502 25170 3554
rect 25170 3502 25172 3554
rect 25116 3500 25172 3502
rect 25228 3388 25284 3444
rect 25452 3388 25508 3444
rect 25900 6802 25956 6804
rect 25900 6750 25902 6802
rect 25902 6750 25954 6802
rect 25954 6750 25956 6802
rect 25900 6748 25956 6750
rect 28554 8650 28610 8652
rect 28554 8598 28556 8650
rect 28556 8598 28608 8650
rect 28608 8598 28610 8650
rect 28554 8596 28610 8598
rect 28658 8650 28714 8652
rect 28658 8598 28660 8650
rect 28660 8598 28712 8650
rect 28712 8598 28714 8650
rect 28658 8596 28714 8598
rect 28762 8650 28818 8652
rect 28762 8598 28764 8650
rect 28764 8598 28816 8650
rect 28816 8598 28818 8650
rect 28762 8596 28818 8598
rect 28700 8428 28756 8484
rect 28364 7756 28420 7812
rect 26908 6578 26964 6580
rect 26908 6526 26910 6578
rect 26910 6526 26962 6578
rect 26962 6526 26964 6578
rect 26908 6524 26964 6526
rect 27356 6076 27412 6132
rect 25788 6018 25844 6020
rect 25788 5966 25790 6018
rect 25790 5966 25842 6018
rect 25842 5966 25844 6018
rect 25788 5964 25844 5966
rect 26236 5404 26292 5460
rect 26124 4956 26180 5012
rect 26012 3666 26068 3668
rect 26012 3614 26014 3666
rect 26014 3614 26066 3666
rect 26066 3614 26068 3666
rect 26012 3612 26068 3614
rect 26572 5010 26628 5012
rect 26572 4958 26574 5010
rect 26574 4958 26626 5010
rect 26626 4958 26628 5010
rect 26572 4956 26628 4958
rect 27132 4732 27188 4788
rect 26796 4562 26852 4564
rect 26796 4510 26798 4562
rect 26798 4510 26850 4562
rect 26850 4510 26852 4562
rect 26796 4508 26852 4510
rect 28554 7082 28610 7084
rect 28554 7030 28556 7082
rect 28556 7030 28608 7082
rect 28608 7030 28610 7082
rect 28554 7028 28610 7030
rect 28658 7082 28714 7084
rect 28658 7030 28660 7082
rect 28660 7030 28712 7082
rect 28712 7030 28714 7082
rect 28658 7028 28714 7030
rect 28762 7082 28818 7084
rect 28762 7030 28764 7082
rect 28764 7030 28816 7082
rect 28816 7030 28818 7082
rect 28762 7028 28818 7030
rect 28476 6860 28532 6916
rect 28554 5514 28610 5516
rect 28554 5462 28556 5514
rect 28556 5462 28608 5514
rect 28608 5462 28610 5514
rect 28554 5460 28610 5462
rect 28658 5514 28714 5516
rect 28658 5462 28660 5514
rect 28660 5462 28712 5514
rect 28712 5462 28714 5514
rect 28658 5460 28714 5462
rect 28762 5514 28818 5516
rect 28762 5462 28764 5514
rect 28764 5462 28816 5514
rect 28816 5462 28818 5514
rect 28762 5460 28818 5462
rect 27580 5234 27636 5236
rect 27580 5182 27582 5234
rect 27582 5182 27634 5234
rect 27634 5182 27636 5234
rect 27580 5180 27636 5182
rect 28140 4956 28196 5012
rect 27468 4508 27524 4564
rect 27692 4508 27748 4564
rect 27580 4060 27636 4116
rect 26908 3388 26964 3444
rect 28700 4562 28756 4564
rect 28700 4510 28702 4562
rect 28702 4510 28754 4562
rect 28754 4510 28756 4562
rect 28700 4508 28756 4510
rect 28252 3836 28308 3892
rect 28554 3946 28610 3948
rect 28554 3894 28556 3946
rect 28556 3894 28608 3946
rect 28608 3894 28610 3946
rect 28554 3892 28610 3894
rect 28658 3946 28714 3948
rect 28658 3894 28660 3946
rect 28660 3894 28712 3946
rect 28712 3894 28714 3946
rect 28658 3892 28714 3894
rect 28762 3946 28818 3948
rect 28762 3894 28764 3946
rect 28764 3894 28816 3946
rect 28816 3894 28818 3946
rect 28762 3892 28818 3894
rect 28588 3724 28644 3780
rect 28812 3724 28868 3780
rect 29036 6860 29092 6916
rect 29148 9996 29204 10052
rect 29260 8034 29316 8036
rect 29260 7982 29262 8034
rect 29262 7982 29314 8034
rect 29314 7982 29316 8034
rect 29260 7980 29316 7982
rect 30268 20636 30324 20692
rect 30156 19346 30212 19348
rect 30156 19294 30158 19346
rect 30158 19294 30210 19346
rect 30210 19294 30212 19346
rect 30156 19292 30212 19294
rect 30156 17778 30212 17780
rect 30156 17726 30158 17778
rect 30158 17726 30210 17778
rect 30210 17726 30212 17778
rect 30156 17724 30212 17726
rect 30044 16770 30100 16772
rect 30044 16718 30046 16770
rect 30046 16718 30098 16770
rect 30098 16718 30100 16770
rect 30044 16716 30100 16718
rect 30156 16604 30212 16660
rect 31500 28082 31556 28084
rect 31500 28030 31502 28082
rect 31502 28030 31554 28082
rect 31554 28030 31556 28082
rect 31500 28028 31556 28030
rect 31276 27020 31332 27076
rect 31948 28530 32004 28532
rect 31948 28478 31950 28530
rect 31950 28478 32002 28530
rect 32002 28478 32004 28530
rect 31948 28476 32004 28478
rect 31724 27020 31780 27076
rect 31164 26908 31220 26964
rect 31164 21868 31220 21924
rect 31052 20524 31108 20580
rect 30940 19068 30996 19124
rect 31276 18450 31332 18452
rect 31276 18398 31278 18450
rect 31278 18398 31330 18450
rect 31330 18398 31332 18450
rect 31276 18396 31332 18398
rect 31500 24892 31556 24948
rect 31500 22876 31556 22932
rect 31500 21420 31556 21476
rect 31500 19404 31556 19460
rect 31164 18172 31220 18228
rect 30492 17836 30548 17892
rect 31164 17554 31220 17556
rect 31164 17502 31166 17554
rect 31166 17502 31218 17554
rect 31218 17502 31220 17554
rect 31164 17500 31220 17502
rect 29932 10668 29988 10724
rect 29708 8428 29764 8484
rect 29372 6636 29428 6692
rect 29036 5628 29092 5684
rect 29036 3612 29092 3668
rect 30156 16210 30212 16212
rect 30156 16158 30158 16210
rect 30158 16158 30210 16210
rect 30210 16158 30212 16210
rect 30156 16156 30212 16158
rect 32172 29314 32228 29316
rect 32172 29262 32174 29314
rect 32174 29262 32226 29314
rect 32226 29262 32228 29314
rect 32172 29260 32228 29262
rect 32460 29818 32516 29820
rect 32460 29766 32462 29818
rect 32462 29766 32514 29818
rect 32514 29766 32516 29818
rect 32460 29764 32516 29766
rect 32564 29818 32620 29820
rect 32564 29766 32566 29818
rect 32566 29766 32618 29818
rect 32618 29766 32620 29818
rect 32564 29764 32620 29766
rect 32668 29818 32724 29820
rect 32668 29766 32670 29818
rect 32670 29766 32722 29818
rect 32722 29766 32724 29818
rect 32668 29764 32724 29766
rect 32460 28250 32516 28252
rect 32460 28198 32462 28250
rect 32462 28198 32514 28250
rect 32514 28198 32516 28250
rect 32460 28196 32516 28198
rect 32564 28250 32620 28252
rect 32564 28198 32566 28250
rect 32566 28198 32618 28250
rect 32618 28198 32620 28250
rect 32564 28196 32620 28198
rect 32668 28250 32724 28252
rect 32668 28198 32670 28250
rect 32670 28198 32722 28250
rect 32722 28198 32724 28250
rect 32668 28196 32724 28198
rect 32172 25564 32228 25620
rect 32460 26682 32516 26684
rect 32460 26630 32462 26682
rect 32462 26630 32514 26682
rect 32514 26630 32516 26682
rect 32460 26628 32516 26630
rect 32564 26682 32620 26684
rect 32564 26630 32566 26682
rect 32566 26630 32618 26682
rect 32618 26630 32620 26682
rect 32564 26628 32620 26630
rect 32668 26682 32724 26684
rect 32668 26630 32670 26682
rect 32670 26630 32722 26682
rect 32722 26630 32724 26682
rect 32668 26628 32724 26630
rect 32460 25114 32516 25116
rect 32460 25062 32462 25114
rect 32462 25062 32514 25114
rect 32514 25062 32516 25114
rect 32460 25060 32516 25062
rect 32564 25114 32620 25116
rect 32564 25062 32566 25114
rect 32566 25062 32618 25114
rect 32618 25062 32620 25114
rect 32564 25060 32620 25062
rect 32668 25114 32724 25116
rect 32668 25062 32670 25114
rect 32670 25062 32722 25114
rect 32722 25062 32724 25114
rect 32668 25060 32724 25062
rect 32284 24946 32340 24948
rect 32284 24894 32286 24946
rect 32286 24894 32338 24946
rect 32338 24894 32340 24946
rect 32284 24892 32340 24894
rect 32460 23546 32516 23548
rect 32460 23494 32462 23546
rect 32462 23494 32514 23546
rect 32514 23494 32516 23546
rect 32460 23492 32516 23494
rect 32564 23546 32620 23548
rect 32564 23494 32566 23546
rect 32566 23494 32618 23546
rect 32618 23494 32620 23546
rect 32564 23492 32620 23494
rect 32668 23546 32724 23548
rect 32668 23494 32670 23546
rect 32670 23494 32722 23546
rect 32722 23494 32724 23546
rect 32668 23492 32724 23494
rect 32460 21978 32516 21980
rect 32460 21926 32462 21978
rect 32462 21926 32514 21978
rect 32514 21926 32516 21978
rect 32460 21924 32516 21926
rect 32564 21978 32620 21980
rect 32564 21926 32566 21978
rect 32566 21926 32618 21978
rect 32618 21926 32620 21978
rect 32564 21924 32620 21926
rect 32668 21978 32724 21980
rect 32668 21926 32670 21978
rect 32670 21926 32722 21978
rect 32722 21926 32724 21978
rect 32668 21924 32724 21926
rect 31836 21420 31892 21476
rect 31948 20188 32004 20244
rect 32172 21474 32228 21476
rect 32172 21422 32174 21474
rect 32174 21422 32226 21474
rect 32226 21422 32228 21474
rect 32172 21420 32228 21422
rect 32460 20410 32516 20412
rect 32460 20358 32462 20410
rect 32462 20358 32514 20410
rect 32514 20358 32516 20410
rect 32460 20356 32516 20358
rect 32564 20410 32620 20412
rect 32564 20358 32566 20410
rect 32566 20358 32618 20410
rect 32618 20358 32620 20410
rect 32564 20356 32620 20358
rect 32668 20410 32724 20412
rect 32668 20358 32670 20410
rect 32670 20358 32722 20410
rect 32722 20358 32724 20410
rect 32668 20356 32724 20358
rect 32460 18842 32516 18844
rect 32460 18790 32462 18842
rect 32462 18790 32514 18842
rect 32514 18790 32516 18842
rect 32460 18788 32516 18790
rect 32564 18842 32620 18844
rect 32564 18790 32566 18842
rect 32566 18790 32618 18842
rect 32618 18790 32620 18842
rect 32564 18788 32620 18790
rect 32668 18842 32724 18844
rect 32668 18790 32670 18842
rect 32670 18790 32722 18842
rect 32722 18790 32724 18842
rect 32668 18788 32724 18790
rect 32060 18396 32116 18452
rect 31948 18284 32004 18340
rect 32060 17612 32116 17668
rect 32460 17274 32516 17276
rect 32460 17222 32462 17274
rect 32462 17222 32514 17274
rect 32514 17222 32516 17274
rect 32460 17220 32516 17222
rect 32564 17274 32620 17276
rect 32564 17222 32566 17274
rect 32566 17222 32618 17274
rect 32618 17222 32620 17274
rect 32564 17220 32620 17222
rect 32668 17274 32724 17276
rect 32668 17222 32670 17274
rect 32670 17222 32722 17274
rect 32722 17222 32724 17274
rect 32668 17220 32724 17222
rect 31164 15986 31220 15988
rect 31164 15934 31166 15986
rect 31166 15934 31218 15986
rect 31218 15934 31220 15986
rect 31164 15932 31220 15934
rect 31052 15596 31108 15652
rect 32460 15706 32516 15708
rect 32460 15654 32462 15706
rect 32462 15654 32514 15706
rect 32514 15654 32516 15706
rect 32460 15652 32516 15654
rect 32564 15706 32620 15708
rect 32564 15654 32566 15706
rect 32566 15654 32618 15706
rect 32618 15654 32620 15706
rect 32564 15652 32620 15654
rect 32668 15706 32724 15708
rect 32668 15654 32670 15706
rect 32670 15654 32722 15706
rect 32722 15654 32724 15706
rect 32668 15652 32724 15654
rect 30716 15036 30772 15092
rect 30156 14642 30212 14644
rect 30156 14590 30158 14642
rect 30158 14590 30210 14642
rect 30210 14590 30212 14642
rect 30156 14588 30212 14590
rect 30716 14252 30772 14308
rect 30380 14140 30436 14196
rect 30156 14028 30212 14084
rect 30156 11004 30212 11060
rect 30268 11116 30324 11172
rect 30044 10108 30100 10164
rect 30156 10780 30212 10836
rect 30044 9884 30100 9940
rect 30604 10722 30660 10724
rect 30604 10670 30606 10722
rect 30606 10670 30658 10722
rect 30658 10670 30660 10722
rect 30604 10668 30660 10670
rect 30940 10610 30996 10612
rect 30940 10558 30942 10610
rect 30942 10558 30994 10610
rect 30994 10558 30996 10610
rect 30940 10556 30996 10558
rect 30156 8764 30212 8820
rect 30156 7756 30212 7812
rect 31612 15036 31668 15092
rect 31276 13580 31332 13636
rect 31164 11282 31220 11284
rect 31164 11230 31166 11282
rect 31166 11230 31218 11282
rect 31218 11230 31220 11282
rect 31164 11228 31220 11230
rect 31164 9714 31220 9716
rect 31164 9662 31166 9714
rect 31166 9662 31218 9714
rect 31218 9662 31220 9714
rect 31164 9660 31220 9662
rect 32060 14306 32116 14308
rect 32060 14254 32062 14306
rect 32062 14254 32114 14306
rect 32114 14254 32116 14306
rect 32060 14252 32116 14254
rect 32460 14138 32516 14140
rect 32460 14086 32462 14138
rect 32462 14086 32514 14138
rect 32514 14086 32516 14138
rect 32460 14084 32516 14086
rect 32564 14138 32620 14140
rect 32564 14086 32566 14138
rect 32566 14086 32618 14138
rect 32618 14086 32620 14138
rect 32564 14084 32620 14086
rect 32668 14138 32724 14140
rect 32668 14086 32670 14138
rect 32670 14086 32722 14138
rect 32722 14086 32724 14138
rect 32668 14084 32724 14086
rect 32460 12570 32516 12572
rect 32460 12518 32462 12570
rect 32462 12518 32514 12570
rect 32514 12518 32516 12570
rect 32460 12516 32516 12518
rect 32564 12570 32620 12572
rect 32564 12518 32566 12570
rect 32566 12518 32618 12570
rect 32618 12518 32620 12570
rect 32564 12516 32620 12518
rect 32668 12570 32724 12572
rect 32668 12518 32670 12570
rect 32670 12518 32722 12570
rect 32722 12518 32724 12570
rect 32668 12516 32724 12518
rect 32060 11506 32116 11508
rect 32060 11454 32062 11506
rect 32062 11454 32114 11506
rect 32114 11454 32116 11506
rect 32060 11452 32116 11454
rect 32460 11002 32516 11004
rect 32460 10950 32462 11002
rect 32462 10950 32514 11002
rect 32514 10950 32516 11002
rect 32460 10948 32516 10950
rect 32564 11002 32620 11004
rect 32564 10950 32566 11002
rect 32566 10950 32618 11002
rect 32618 10950 32620 11002
rect 32564 10948 32620 10950
rect 32668 11002 32724 11004
rect 32668 10950 32670 11002
rect 32670 10950 32722 11002
rect 32722 10950 32724 11002
rect 32668 10948 32724 10950
rect 32284 10722 32340 10724
rect 32284 10670 32286 10722
rect 32286 10670 32338 10722
rect 32338 10670 32340 10722
rect 32284 10668 32340 10670
rect 31724 9772 31780 9828
rect 31164 8146 31220 8148
rect 31164 8094 31166 8146
rect 31166 8094 31218 8146
rect 31218 8094 31220 8146
rect 31164 8092 31220 8094
rect 32172 9996 32228 10052
rect 32460 9434 32516 9436
rect 32460 9382 32462 9434
rect 32462 9382 32514 9434
rect 32514 9382 32516 9434
rect 32460 9380 32516 9382
rect 32564 9434 32620 9436
rect 32564 9382 32566 9434
rect 32566 9382 32618 9434
rect 32618 9382 32620 9434
rect 32564 9380 32620 9382
rect 32668 9434 32724 9436
rect 32668 9382 32670 9434
rect 32670 9382 32722 9434
rect 32722 9382 32724 9434
rect 32668 9380 32724 9382
rect 31836 7420 31892 7476
rect 29932 5852 29988 5908
rect 31164 6636 31220 6692
rect 31052 5852 31108 5908
rect 29820 4284 29876 4340
rect 30044 5068 30100 5124
rect 32460 7866 32516 7868
rect 32460 7814 32462 7866
rect 32462 7814 32514 7866
rect 32514 7814 32516 7866
rect 32460 7812 32516 7814
rect 32564 7866 32620 7868
rect 32564 7814 32566 7866
rect 32566 7814 32618 7866
rect 32618 7814 32620 7866
rect 32564 7812 32620 7814
rect 32668 7866 32724 7868
rect 32668 7814 32670 7866
rect 32670 7814 32722 7866
rect 32722 7814 32724 7866
rect 32668 7812 32724 7814
rect 31388 5180 31444 5236
rect 31164 4732 31220 4788
rect 31612 4338 31668 4340
rect 31612 4286 31614 4338
rect 31614 4286 31666 4338
rect 31666 4286 31668 4338
rect 31612 4284 31668 4286
rect 28812 2044 28868 2100
rect 30156 1372 30212 1428
rect 32460 6298 32516 6300
rect 32460 6246 32462 6298
rect 32462 6246 32514 6298
rect 32514 6246 32516 6298
rect 32460 6244 32516 6246
rect 32564 6298 32620 6300
rect 32564 6246 32566 6298
rect 32566 6246 32618 6298
rect 32618 6246 32620 6298
rect 32564 6244 32620 6246
rect 32668 6298 32724 6300
rect 32668 6246 32670 6298
rect 32670 6246 32722 6298
rect 32722 6246 32724 6298
rect 32668 6244 32724 6246
rect 32460 4730 32516 4732
rect 32460 4678 32462 4730
rect 32462 4678 32514 4730
rect 32514 4678 32516 4730
rect 32460 4676 32516 4678
rect 32564 4730 32620 4732
rect 32564 4678 32566 4730
rect 32566 4678 32618 4730
rect 32618 4678 32620 4730
rect 32564 4676 32620 4678
rect 32668 4730 32724 4732
rect 32668 4678 32670 4730
rect 32670 4678 32722 4730
rect 32722 4678 32724 4730
rect 32668 4676 32724 4678
rect 32284 4060 32340 4116
rect 32460 3162 32516 3164
rect 32460 3110 32462 3162
rect 32462 3110 32514 3162
rect 32514 3110 32516 3162
rect 32460 3108 32516 3110
rect 32564 3162 32620 3164
rect 32564 3110 32566 3162
rect 32566 3110 32618 3162
rect 32618 3110 32620 3162
rect 32564 3108 32620 3110
rect 32668 3162 32724 3164
rect 32668 3110 32670 3162
rect 32670 3110 32722 3162
rect 32722 3110 32724 3162
rect 32668 3108 32724 3110
rect 32172 2716 32228 2772
rect 32060 700 32116 756
<< metal3 >>
rect 0 33684 800 33712
rect 0 33628 4676 33684
rect 0 33600 800 33628
rect 0 33012 800 33040
rect 4620 33012 4676 33628
rect 0 32956 980 33012
rect 4610 32956 4620 33012
rect 4676 32956 4686 33012
rect 0 32928 800 32956
rect 924 32900 980 32956
rect 924 32844 1820 32900
rect 1876 32844 1886 32900
rect 0 32340 800 32368
rect 0 32284 3724 32340
rect 3780 32284 3790 32340
rect 0 32256 800 32284
rect 0 31668 800 31696
rect 33200 31668 34000 31696
rect 0 31612 3612 31668
rect 3668 31612 3678 31668
rect 32274 31612 32284 31668
rect 32340 31612 34000 31668
rect 0 31584 800 31612
rect 33200 31584 34000 31612
rect 0 30996 800 31024
rect 33200 30996 34000 31024
rect 0 30940 2156 30996
rect 2212 30940 2222 30996
rect 29922 30940 29932 30996
rect 29988 30940 34000 30996
rect 0 30912 800 30940
rect 33200 30912 34000 30940
rect 5108 30548 5118 30604
rect 5174 30548 5222 30604
rect 5278 30548 5326 30604
rect 5382 30548 5392 30604
rect 12920 30548 12930 30604
rect 12986 30548 13034 30604
rect 13090 30548 13138 30604
rect 13194 30548 13204 30604
rect 20732 30548 20742 30604
rect 20798 30548 20846 30604
rect 20902 30548 20950 30604
rect 21006 30548 21016 30604
rect 28544 30548 28554 30604
rect 28610 30548 28658 30604
rect 28714 30548 28762 30604
rect 28818 30548 28828 30604
rect 1820 30380 6636 30436
rect 6692 30380 6702 30436
rect 8642 30380 8652 30436
rect 8708 30380 13244 30436
rect 13300 30380 13310 30436
rect 0 30324 800 30352
rect 1820 30324 1876 30380
rect 33200 30324 34000 30352
rect 0 30268 1876 30324
rect 2034 30268 2044 30324
rect 2100 30268 9436 30324
rect 9492 30268 9502 30324
rect 11890 30268 11900 30324
rect 11956 30268 14924 30324
rect 14980 30268 14990 30324
rect 32050 30268 32060 30324
rect 32116 30268 34000 30324
rect 0 30240 800 30268
rect 33200 30240 34000 30268
rect 3378 30156 3388 30212
rect 3444 30156 9324 30212
rect 9380 30156 9390 30212
rect 13570 30156 13580 30212
rect 13636 30156 14028 30212
rect 14084 30156 16156 30212
rect 16212 30156 16222 30212
rect 18162 30156 18172 30212
rect 18228 30156 19964 30212
rect 20020 30156 21420 30212
rect 21476 30156 21486 30212
rect 25218 30156 25228 30212
rect 25284 30156 26348 30212
rect 26404 30156 26414 30212
rect 26786 30156 26796 30212
rect 26852 30156 27580 30212
rect 27636 30156 27646 30212
rect 4946 30044 4956 30100
rect 5012 30044 6972 30100
rect 7028 30044 7038 30100
rect 9762 30044 9772 30100
rect 9828 30044 12012 30100
rect 12068 30044 15484 30100
rect 15540 30044 15550 30100
rect 20178 30044 20188 30100
rect 20244 30044 23548 30100
rect 23604 30044 23614 30100
rect 24770 30044 24780 30100
rect 24836 30044 28252 30100
rect 28308 30044 28318 30100
rect 4162 29932 4172 29988
rect 4228 29932 6748 29988
rect 6804 29932 6814 29988
rect 8642 29932 8652 29988
rect 8708 29932 19404 29988
rect 19460 29932 19470 29988
rect 24882 29932 24892 29988
rect 24948 29932 25900 29988
rect 25956 29932 25966 29988
rect 5618 29820 5628 29876
rect 5684 29820 6412 29876
rect 6468 29820 6478 29876
rect 9986 29820 9996 29876
rect 10052 29820 13468 29876
rect 13524 29820 13534 29876
rect 17490 29820 17500 29876
rect 17556 29820 21868 29876
rect 21924 29820 21934 29876
rect 9014 29764 9024 29820
rect 9080 29764 9128 29820
rect 9184 29764 9232 29820
rect 9288 29764 9298 29820
rect 16826 29764 16836 29820
rect 16892 29764 16940 29820
rect 16996 29764 17044 29820
rect 17100 29764 17110 29820
rect 24638 29764 24648 29820
rect 24704 29764 24752 29820
rect 24808 29764 24856 29820
rect 24912 29764 24922 29820
rect 32450 29764 32460 29820
rect 32516 29764 32564 29820
rect 32620 29764 32668 29820
rect 32724 29764 32734 29820
rect 3266 29708 3276 29764
rect 3332 29708 3836 29764
rect 3892 29708 3902 29764
rect 5730 29708 5740 29764
rect 5796 29708 8764 29764
rect 8820 29708 8830 29764
rect 0 29652 800 29680
rect 33200 29652 34000 29680
rect 0 29596 3948 29652
rect 4004 29596 4014 29652
rect 7634 29596 7644 29652
rect 7700 29596 9548 29652
rect 9604 29596 9614 29652
rect 10770 29596 10780 29652
rect 10836 29596 14812 29652
rect 14868 29596 14878 29652
rect 23986 29596 23996 29652
rect 24052 29596 24556 29652
rect 24612 29596 26908 29652
rect 26964 29596 27356 29652
rect 27412 29596 27422 29652
rect 28018 29596 28028 29652
rect 28084 29596 34000 29652
rect 0 29568 800 29596
rect 33200 29568 34000 29596
rect 2258 29484 2268 29540
rect 2324 29484 8428 29540
rect 8754 29484 8764 29540
rect 8820 29484 9996 29540
rect 10052 29484 10062 29540
rect 12002 29484 12012 29540
rect 12068 29484 17052 29540
rect 17108 29484 17118 29540
rect 21298 29484 21308 29540
rect 21364 29484 27244 29540
rect 27300 29484 27310 29540
rect 8372 29428 8428 29484
rect 1922 29372 1932 29428
rect 1988 29372 2940 29428
rect 2996 29372 3006 29428
rect 8372 29372 10108 29428
rect 10164 29372 10174 29428
rect 22642 29372 22652 29428
rect 22708 29372 24332 29428
rect 24388 29372 25340 29428
rect 25396 29372 25406 29428
rect 2594 29260 2604 29316
rect 2660 29260 4172 29316
rect 4228 29260 4238 29316
rect 6850 29260 6860 29316
rect 6916 29260 8428 29316
rect 9538 29260 9548 29316
rect 9604 29260 11340 29316
rect 11396 29260 11406 29316
rect 13010 29260 13020 29316
rect 13076 29260 17724 29316
rect 17780 29260 17790 29316
rect 22530 29260 22540 29316
rect 22596 29260 26236 29316
rect 26292 29260 26302 29316
rect 30930 29260 30940 29316
rect 30996 29260 32172 29316
rect 32228 29260 32238 29316
rect 8372 29204 8428 29260
rect 3042 29148 3052 29204
rect 3108 29148 4396 29204
rect 4452 29148 4462 29204
rect 5170 29148 5180 29204
rect 5236 29148 6188 29204
rect 6244 29148 6254 29204
rect 8372 29148 10220 29204
rect 10276 29148 10286 29204
rect 16258 29148 16268 29204
rect 16324 29148 22876 29204
rect 22932 29148 22942 29204
rect 23650 29148 23660 29204
rect 23716 29148 27468 29204
rect 27524 29148 27534 29204
rect 4050 29036 4060 29092
rect 4116 29036 4956 29092
rect 5012 29036 5022 29092
rect 0 28980 800 29008
rect 5108 28980 5118 29036
rect 5174 28980 5222 29036
rect 5278 28980 5326 29036
rect 5382 28980 5392 29036
rect 12920 28980 12930 29036
rect 12986 28980 13034 29036
rect 13090 28980 13138 29036
rect 13194 28980 13204 29036
rect 20732 28980 20742 29036
rect 20798 28980 20846 29036
rect 20902 28980 20950 29036
rect 21006 28980 21016 29036
rect 28544 28980 28554 29036
rect 28610 28980 28658 29036
rect 28714 28980 28762 29036
rect 28818 28980 28828 29036
rect 33200 28980 34000 29008
rect 0 28924 980 28980
rect 7298 28924 7308 28980
rect 7364 28924 10332 28980
rect 10388 28924 10398 28980
rect 23314 28924 23324 28980
rect 23380 28924 26684 28980
rect 26740 28924 26750 28980
rect 31892 28924 34000 28980
rect 0 28896 800 28924
rect 924 28756 980 28924
rect 1362 28812 1372 28868
rect 1428 28812 10388 28868
rect 10546 28812 10556 28868
rect 10612 28812 17164 28868
rect 17220 28812 17230 28868
rect 20850 28812 20860 28868
rect 20916 28812 21308 28868
rect 21364 28812 21374 28868
rect 25890 28812 25900 28868
rect 25956 28812 29036 28868
rect 29092 28812 29102 28868
rect 10332 28756 10388 28812
rect 130 28700 140 28756
rect 196 28700 980 28756
rect 4050 28700 4060 28756
rect 4116 28700 7420 28756
rect 7476 28700 7486 28756
rect 8372 28700 9548 28756
rect 9604 28700 9614 28756
rect 10332 28700 11340 28756
rect 11396 28700 11406 28756
rect 8372 28644 8428 28700
rect 31892 28644 31948 28924
rect 33200 28896 34000 28924
rect 4806 28588 4844 28644
rect 4900 28588 4910 28644
rect 5618 28588 5628 28644
rect 5684 28588 6188 28644
rect 6244 28588 8092 28644
rect 8148 28588 8428 28644
rect 11554 28588 11564 28644
rect 11620 28588 13916 28644
rect 13972 28588 13982 28644
rect 16594 28588 16604 28644
rect 16660 28588 17948 28644
rect 18004 28588 18014 28644
rect 19730 28588 19740 28644
rect 19796 28588 22764 28644
rect 22820 28588 22830 28644
rect 23426 28588 23436 28644
rect 23492 28588 26236 28644
rect 26292 28588 26908 28644
rect 29026 28588 29036 28644
rect 29092 28588 31948 28644
rect 26852 28532 26908 28588
rect 8978 28476 8988 28532
rect 9044 28476 21308 28532
rect 21364 28476 21374 28532
rect 26852 28476 28588 28532
rect 28644 28476 28654 28532
rect 29138 28476 29148 28532
rect 29204 28476 31948 28532
rect 32004 28476 32014 28532
rect 4498 28364 4508 28420
rect 4564 28364 12684 28420
rect 12740 28364 12750 28420
rect 16482 28364 16492 28420
rect 16548 28364 19964 28420
rect 20020 28364 20030 28420
rect 31892 28364 32900 28420
rect 0 28308 800 28336
rect 31892 28308 31948 28364
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 5730 28252 5740 28308
rect 5796 28252 7980 28308
rect 8036 28252 8046 28308
rect 18834 28252 18844 28308
rect 18900 28252 21756 28308
rect 21812 28252 21822 28308
rect 29138 28252 29148 28308
rect 29204 28252 31948 28308
rect 32844 28308 32900 28364
rect 33200 28308 34000 28336
rect 32844 28252 34000 28308
rect 0 28224 800 28252
rect 9014 28196 9024 28252
rect 9080 28196 9128 28252
rect 9184 28196 9232 28252
rect 9288 28196 9298 28252
rect 16826 28196 16836 28252
rect 16892 28196 16940 28252
rect 16996 28196 17044 28252
rect 17100 28196 17110 28252
rect 24638 28196 24648 28252
rect 24704 28196 24752 28252
rect 24808 28196 24856 28252
rect 24912 28196 24922 28252
rect 32450 28196 32460 28252
rect 32516 28196 32564 28252
rect 32620 28196 32668 28252
rect 32724 28196 32734 28252
rect 33200 28224 34000 28252
rect 12114 28140 12124 28196
rect 12180 28140 15932 28196
rect 15988 28140 15998 28196
rect 20066 28140 20076 28196
rect 20132 28140 24332 28196
rect 24388 28140 24398 28196
rect 5954 28028 5964 28084
rect 6020 28028 9548 28084
rect 9604 28028 9614 28084
rect 12562 28028 12572 28084
rect 12628 28028 13692 28084
rect 13748 28028 13758 28084
rect 28914 28028 28924 28084
rect 28980 28028 31500 28084
rect 31556 28028 31566 28084
rect 2146 27916 2156 27972
rect 2212 27916 8764 27972
rect 8820 27916 8830 27972
rect 24098 27916 24108 27972
rect 24164 27916 27244 27972
rect 27300 27916 27310 27972
rect 3154 27804 3164 27860
rect 3220 27804 10108 27860
rect 10164 27804 10174 27860
rect 17154 27804 17164 27860
rect 17220 27804 19180 27860
rect 19236 27804 19246 27860
rect 21634 27804 21644 27860
rect 21700 27804 24444 27860
rect 24500 27804 24510 27860
rect 6066 27692 6076 27748
rect 6132 27692 12236 27748
rect 12292 27692 12302 27748
rect 13906 27692 13916 27748
rect 13972 27692 18732 27748
rect 18788 27692 18798 27748
rect 25218 27692 25228 27748
rect 25284 27692 26236 27748
rect 26292 27692 26302 27748
rect 0 27636 800 27664
rect 33200 27636 34000 27664
rect 0 27580 1764 27636
rect 3042 27580 3052 27636
rect 3108 27580 4396 27636
rect 4452 27580 4462 27636
rect 11778 27580 11788 27636
rect 11844 27580 13132 27636
rect 13188 27580 13198 27636
rect 29362 27580 29372 27636
rect 29428 27580 34000 27636
rect 0 27552 800 27580
rect 1708 27524 1764 27580
rect 33200 27552 34000 27580
rect 1708 27468 3388 27524
rect 3444 27468 3454 27524
rect 5108 27412 5118 27468
rect 5174 27412 5222 27468
rect 5278 27412 5326 27468
rect 5382 27412 5392 27468
rect 12920 27412 12930 27468
rect 12986 27412 13034 27468
rect 13090 27412 13138 27468
rect 13194 27412 13204 27468
rect 20732 27412 20742 27468
rect 20798 27412 20846 27468
rect 20902 27412 20950 27468
rect 21006 27412 21016 27468
rect 28544 27412 28554 27468
rect 28610 27412 28658 27468
rect 28714 27412 28762 27468
rect 28818 27412 28828 27468
rect 22194 27244 22204 27300
rect 22260 27244 30268 27300
rect 30324 27244 30334 27300
rect 2034 27132 2044 27188
rect 2100 27132 4508 27188
rect 4564 27132 4574 27188
rect 7522 27132 7532 27188
rect 7588 27132 13804 27188
rect 13860 27132 13870 27188
rect 2258 27020 2268 27076
rect 2324 27020 9772 27076
rect 9828 27020 9838 27076
rect 9996 27020 11788 27076
rect 11844 27020 11854 27076
rect 12450 27020 12460 27076
rect 12516 27020 13356 27076
rect 13412 27020 13422 27076
rect 14018 27020 14028 27076
rect 14084 27020 15596 27076
rect 15652 27020 15662 27076
rect 24994 27020 25004 27076
rect 25060 27020 31276 27076
rect 31332 27020 31342 27076
rect 31714 27020 31724 27076
rect 31780 27020 31948 27076
rect 0 26964 800 26992
rect 9996 26964 10052 27020
rect 31892 26964 31948 27020
rect 33200 26964 34000 26992
rect 0 26908 4620 26964
rect 4676 26908 4686 26964
rect 6514 26908 6524 26964
rect 6580 26908 10052 26964
rect 10210 26908 10220 26964
rect 10276 26908 14364 26964
rect 14420 26908 14430 26964
rect 16258 26908 16268 26964
rect 16324 26908 17276 26964
rect 17332 26908 18452 26964
rect 20290 26908 20300 26964
rect 20356 26908 21532 26964
rect 21588 26908 21598 26964
rect 21746 26908 21756 26964
rect 21812 26908 22988 26964
rect 23044 26908 23054 26964
rect 25778 26908 25788 26964
rect 25844 26908 28364 26964
rect 28420 26908 28430 26964
rect 29698 26908 29708 26964
rect 29764 26908 31164 26964
rect 31220 26908 31230 26964
rect 31892 26908 34000 26964
rect 0 26880 800 26908
rect 18396 26852 18452 26908
rect 33200 26880 34000 26908
rect 16370 26796 16380 26852
rect 16436 26796 18060 26852
rect 18116 26796 18126 26852
rect 18274 26796 18284 26852
rect 18340 26796 18452 26852
rect 20738 26796 20748 26852
rect 20804 26796 22204 26852
rect 22260 26796 24108 26852
rect 24164 26796 24174 26852
rect 9014 26628 9024 26684
rect 9080 26628 9128 26684
rect 9184 26628 9232 26684
rect 9288 26628 9298 26684
rect 16826 26628 16836 26684
rect 16892 26628 16940 26684
rect 16996 26628 17044 26684
rect 17100 26628 17110 26684
rect 24638 26628 24648 26684
rect 24704 26628 24752 26684
rect 24808 26628 24856 26684
rect 24912 26628 24922 26684
rect 32450 26628 32460 26684
rect 32516 26628 32564 26684
rect 32620 26628 32668 26684
rect 32724 26628 32734 26684
rect 28802 26572 28812 26628
rect 28868 26572 30044 26628
rect 30100 26572 30110 26628
rect 4162 26460 4172 26516
rect 4228 26460 11788 26516
rect 11844 26460 11854 26516
rect 3154 26348 3164 26404
rect 3220 26348 9100 26404
rect 9156 26348 9166 26404
rect 16370 26348 16380 26404
rect 16436 26348 17388 26404
rect 17444 26348 17454 26404
rect 21970 26348 21980 26404
rect 22036 26348 27244 26404
rect 27300 26348 27310 26404
rect 0 26292 800 26320
rect 33200 26292 34000 26320
rect 0 26236 3388 26292
rect 4050 26236 4060 26292
rect 4116 26236 5964 26292
rect 6020 26236 6030 26292
rect 13010 26236 13020 26292
rect 13076 26236 14028 26292
rect 14084 26236 14094 26292
rect 30044 26236 34000 26292
rect 0 26208 800 26236
rect 3332 26180 3388 26236
rect 30044 26180 30100 26236
rect 33200 26208 34000 26236
rect 3332 26124 4228 26180
rect 4172 26068 4228 26124
rect 4396 26124 5068 26180
rect 5124 26124 13692 26180
rect 13748 26124 13758 26180
rect 21074 26124 21084 26180
rect 21140 26124 26236 26180
rect 26292 26124 26302 26180
rect 29698 26124 29708 26180
rect 29764 26124 30100 26180
rect 2146 26012 2156 26068
rect 2212 26012 3388 26068
rect 4162 26012 4172 26068
rect 4228 26012 4238 26068
rect 3332 25956 3388 26012
rect 4396 25956 4452 26124
rect 3332 25900 4452 25956
rect 5108 25844 5118 25900
rect 5174 25844 5222 25900
rect 5278 25844 5326 25900
rect 5382 25844 5392 25900
rect 12920 25844 12930 25900
rect 12986 25844 13034 25900
rect 13090 25844 13138 25900
rect 13194 25844 13204 25900
rect 20732 25844 20742 25900
rect 20798 25844 20846 25900
rect 20902 25844 20950 25900
rect 21006 25844 21016 25900
rect 28544 25844 28554 25900
rect 28610 25844 28658 25900
rect 28714 25844 28762 25900
rect 28818 25844 28828 25900
rect 29250 25788 29260 25844
rect 29316 25788 30716 25844
rect 30772 25788 30782 25844
rect 2370 25676 2380 25732
rect 2436 25676 3556 25732
rect 3714 25676 3724 25732
rect 3780 25676 5516 25732
rect 5572 25676 5582 25732
rect 12898 25676 12908 25732
rect 12964 25676 14028 25732
rect 14084 25676 14588 25732
rect 14644 25676 16828 25732
rect 16884 25676 17612 25732
rect 17668 25676 17678 25732
rect 20066 25676 20076 25732
rect 20132 25676 24892 25732
rect 24948 25676 24958 25732
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 2930 25564 2940 25620
rect 2996 25564 3388 25620
rect 0 25536 800 25564
rect 3332 25284 3388 25564
rect 3500 25396 3556 25676
rect 33200 25620 34000 25648
rect 4722 25564 4732 25620
rect 4788 25564 6860 25620
rect 6916 25564 6926 25620
rect 17826 25564 17836 25620
rect 17892 25564 19292 25620
rect 19348 25564 19358 25620
rect 26674 25564 26684 25620
rect 26740 25564 30156 25620
rect 30212 25564 30222 25620
rect 32162 25564 32172 25620
rect 32228 25564 34000 25620
rect 33200 25536 34000 25564
rect 4162 25452 4172 25508
rect 4228 25452 11116 25508
rect 11172 25452 11182 25508
rect 11778 25452 11788 25508
rect 11844 25452 12460 25508
rect 12516 25452 12526 25508
rect 13794 25452 13804 25508
rect 13860 25452 15260 25508
rect 15316 25452 15326 25508
rect 3500 25340 10164 25396
rect 2594 25228 2604 25284
rect 2660 25228 2940 25284
rect 2996 25228 3006 25284
rect 3332 25228 4620 25284
rect 4676 25228 4732 25284
rect 4788 25228 4798 25284
rect 5730 25228 5740 25284
rect 5796 25228 6412 25284
rect 6468 25228 7756 25284
rect 7812 25228 8372 25284
rect 8316 25172 8372 25228
rect 10108 25172 10164 25340
rect 11330 25228 11340 25284
rect 11396 25228 13916 25284
rect 13972 25228 13982 25284
rect 21074 25228 21084 25284
rect 21140 25228 22316 25284
rect 22372 25228 22382 25284
rect 26562 25228 26572 25284
rect 26628 25228 27132 25284
rect 27188 25228 27198 25284
rect 27906 25228 27916 25284
rect 27972 25228 29036 25284
rect 29092 25228 29102 25284
rect 802 25116 812 25172
rect 868 25116 8092 25172
rect 8148 25116 8158 25172
rect 8316 25116 8540 25172
rect 8596 25116 8606 25172
rect 10108 25116 15148 25172
rect 9014 25060 9024 25116
rect 9080 25060 9128 25116
rect 9184 25060 9232 25116
rect 9288 25060 9298 25116
rect 2034 25004 2044 25060
rect 2100 25004 6300 25060
rect 6356 25004 6366 25060
rect 10770 25004 10780 25060
rect 10836 25004 12796 25060
rect 12852 25004 12862 25060
rect 0 24948 800 24976
rect 15092 24948 15148 25116
rect 16826 25060 16836 25116
rect 16892 25060 16940 25116
rect 16996 25060 17044 25116
rect 17100 25060 17110 25116
rect 24638 25060 24648 25116
rect 24704 25060 24752 25116
rect 24808 25060 24856 25116
rect 24912 25060 24922 25116
rect 32450 25060 32460 25116
rect 32516 25060 32564 25116
rect 32620 25060 32668 25116
rect 32724 25060 32734 25116
rect 0 24892 3388 24948
rect 7746 24892 7756 24948
rect 7812 24892 8204 24948
rect 8260 24892 8652 24948
rect 8708 24892 11676 24948
rect 11732 24892 11742 24948
rect 15092 24892 15484 24948
rect 15540 24892 15550 24948
rect 16594 24892 16604 24948
rect 16660 24892 19740 24948
rect 19796 24892 19806 24948
rect 31490 24892 31500 24948
rect 31556 24892 32284 24948
rect 32340 24892 32350 24948
rect 0 24864 800 24892
rect 3332 24612 3388 24892
rect 4946 24780 4956 24836
rect 5012 24780 5964 24836
rect 6020 24780 6030 24836
rect 7298 24780 7308 24836
rect 7364 24780 14812 24836
rect 14868 24780 14878 24836
rect 15092 24780 15260 24836
rect 15316 24780 15326 24836
rect 20514 24780 20524 24836
rect 20580 24780 23660 24836
rect 23716 24780 23726 24836
rect 23986 24780 23996 24836
rect 24052 24780 24332 24836
rect 24388 24780 28252 24836
rect 28308 24780 28318 24836
rect 15092 24724 15148 24780
rect 3490 24668 3500 24724
rect 3556 24668 4788 24724
rect 8530 24668 8540 24724
rect 8596 24668 8988 24724
rect 9044 24668 9884 24724
rect 9940 24668 10780 24724
rect 10836 24668 10846 24724
rect 11554 24668 11564 24724
rect 11620 24668 13244 24724
rect 13300 24668 13310 24724
rect 13468 24668 15148 24724
rect 17714 24668 17724 24724
rect 17780 24668 18396 24724
rect 18452 24668 18956 24724
rect 19012 24668 21532 24724
rect 21588 24668 21598 24724
rect 22194 24668 22204 24724
rect 22260 24668 23212 24724
rect 23268 24668 23278 24724
rect 4732 24612 4788 24668
rect 13468 24612 13524 24668
rect 1894 24556 1932 24612
rect 1988 24556 2940 24612
rect 2996 24556 3006 24612
rect 3332 24556 4676 24612
rect 4732 24556 9772 24612
rect 9828 24556 9838 24612
rect 10994 24556 11004 24612
rect 11060 24556 13524 24612
rect 14690 24556 14700 24612
rect 14756 24556 17612 24612
rect 17668 24556 17678 24612
rect 26562 24556 26572 24612
rect 26628 24556 28364 24612
rect 28420 24556 28430 24612
rect 4620 24500 4676 24556
rect 3042 24444 3052 24500
rect 3108 24444 4172 24500
rect 4228 24444 4238 24500
rect 4620 24444 15148 24500
rect 0 24276 800 24304
rect 5108 24276 5118 24332
rect 5174 24276 5222 24332
rect 5278 24276 5326 24332
rect 5382 24276 5392 24332
rect 12920 24276 12930 24332
rect 12986 24276 13034 24332
rect 13090 24276 13138 24332
rect 13194 24276 13204 24332
rect 0 24220 3948 24276
rect 4004 24220 4014 24276
rect 0 24192 800 24220
rect 9650 24108 9660 24164
rect 9716 24108 10220 24164
rect 10276 24108 11564 24164
rect 11620 24108 11630 24164
rect 15092 24052 15148 24444
rect 20732 24276 20742 24332
rect 20798 24276 20846 24332
rect 20902 24276 20950 24332
rect 21006 24276 21016 24332
rect 28544 24276 28554 24332
rect 28610 24276 28658 24332
rect 28714 24276 28762 24332
rect 28818 24276 28828 24332
rect 21186 24220 21196 24276
rect 21252 24220 27244 24276
rect 27300 24220 27310 24276
rect 20514 24108 20524 24164
rect 20580 24108 21644 24164
rect 21700 24108 22988 24164
rect 23044 24108 23996 24164
rect 24052 24108 24062 24164
rect 2034 23996 2044 24052
rect 2100 23996 4508 24052
rect 4564 23996 10668 24052
rect 10724 23996 10734 24052
rect 15092 23996 15260 24052
rect 15316 23996 15326 24052
rect 3714 23884 3724 23940
rect 3780 23884 4172 23940
rect 4228 23884 5068 23940
rect 5124 23884 6300 23940
rect 6356 23884 6366 23940
rect 12226 23884 12236 23940
rect 12292 23884 13916 23940
rect 13972 23884 13982 23940
rect 9090 23772 9100 23828
rect 9156 23772 10108 23828
rect 10164 23772 11340 23828
rect 11396 23772 12796 23828
rect 12852 23772 12862 23828
rect 20290 23772 20300 23828
rect 20356 23772 21308 23828
rect 21364 23772 21374 23828
rect 8306 23660 8316 23716
rect 8372 23660 9548 23716
rect 9604 23660 9614 23716
rect 0 23604 800 23632
rect 0 23548 3500 23604
rect 3556 23548 3566 23604
rect 9650 23548 9660 23604
rect 9716 23548 10332 23604
rect 10388 23548 10398 23604
rect 0 23520 800 23548
rect 9014 23492 9024 23548
rect 9080 23492 9128 23548
rect 9184 23492 9232 23548
rect 9288 23492 9298 23548
rect 16826 23492 16836 23548
rect 16892 23492 16940 23548
rect 16996 23492 17044 23548
rect 17100 23492 17110 23548
rect 24638 23492 24648 23548
rect 24704 23492 24752 23548
rect 24808 23492 24856 23548
rect 24912 23492 24922 23548
rect 32450 23492 32460 23548
rect 32516 23492 32564 23548
rect 32620 23492 32668 23548
rect 32724 23492 32734 23548
rect 9426 23436 9436 23492
rect 9492 23436 14140 23492
rect 14196 23436 14206 23492
rect 17714 23324 17724 23380
rect 17780 23324 27020 23380
rect 27076 23324 27086 23380
rect 16370 23212 16380 23268
rect 16436 23212 18060 23268
rect 18116 23212 18126 23268
rect 18722 23212 18732 23268
rect 18788 23212 20524 23268
rect 20580 23212 20590 23268
rect 4050 23100 4060 23156
rect 4116 23100 4956 23156
rect 5012 23100 5022 23156
rect 8082 23100 8092 23156
rect 8148 23100 10780 23156
rect 10836 23100 10846 23156
rect 16706 23100 16716 23156
rect 16772 23100 20860 23156
rect 20916 23100 25788 23156
rect 25844 23100 26684 23156
rect 26740 23100 26750 23156
rect 24434 22988 24444 23044
rect 24500 22988 25676 23044
rect 25732 22988 25742 23044
rect 0 22932 800 22960
rect 33200 22932 34000 22960
rect 0 22876 1820 22932
rect 1876 22876 1886 22932
rect 31490 22876 31500 22932
rect 31556 22876 34000 22932
rect 0 22848 800 22876
rect 33200 22848 34000 22876
rect 5108 22708 5118 22764
rect 5174 22708 5222 22764
rect 5278 22708 5326 22764
rect 5382 22708 5392 22764
rect 12920 22708 12930 22764
rect 12986 22708 13034 22764
rect 13090 22708 13138 22764
rect 13194 22708 13204 22764
rect 20732 22708 20742 22764
rect 20798 22708 20846 22764
rect 20902 22708 20950 22764
rect 21006 22708 21016 22764
rect 28544 22708 28554 22764
rect 28610 22708 28658 22764
rect 28714 22708 28762 22764
rect 28818 22708 28828 22764
rect 22978 22652 22988 22708
rect 23044 22652 26236 22708
rect 26292 22652 26302 22708
rect 2258 22540 2268 22596
rect 2324 22540 4172 22596
rect 4228 22540 4238 22596
rect 2146 22428 2156 22484
rect 2212 22428 2222 22484
rect 2482 22428 2492 22484
rect 2548 22428 2558 22484
rect 4610 22428 4620 22484
rect 4676 22428 5068 22484
rect 5124 22428 5628 22484
rect 5684 22428 8540 22484
rect 8596 22428 8606 22484
rect 28130 22428 28140 22484
rect 28196 22428 30156 22484
rect 30212 22428 30222 22484
rect 0 22260 800 22288
rect 2156 22260 2212 22428
rect 0 22204 2212 22260
rect 0 22176 800 22204
rect 2492 22148 2548 22428
rect 12786 22316 12796 22372
rect 12852 22316 13580 22372
rect 13636 22316 13916 22372
rect 13972 22316 15036 22372
rect 15092 22316 15102 22372
rect 22306 22316 22316 22372
rect 22372 22316 24668 22372
rect 24724 22316 25116 22372
rect 25172 22316 25182 22372
rect 11442 22204 11452 22260
rect 11508 22204 12572 22260
rect 12628 22204 12638 22260
rect 2146 22092 2156 22148
rect 2212 22092 2548 22148
rect 4162 22092 4172 22148
rect 4228 22092 4620 22148
rect 4676 22092 4686 22148
rect 4946 22092 4956 22148
rect 5012 22092 6524 22148
rect 6580 22092 6590 22148
rect 7074 22092 7084 22148
rect 7140 22092 12236 22148
rect 12292 22092 12302 22148
rect 16146 22092 16156 22148
rect 16212 22092 17164 22148
rect 17220 22092 18396 22148
rect 18452 22092 19964 22148
rect 20020 22092 20030 22148
rect 20626 22092 20636 22148
rect 20692 22092 25564 22148
rect 25620 22092 25630 22148
rect 2258 21980 2268 22036
rect 2324 21980 3388 22036
rect 3444 21980 3454 22036
rect 9014 21924 9024 21980
rect 9080 21924 9128 21980
rect 9184 21924 9232 21980
rect 9288 21924 9298 21980
rect 16826 21924 16836 21980
rect 16892 21924 16940 21980
rect 16996 21924 17044 21980
rect 17100 21924 17110 21980
rect 24638 21924 24648 21980
rect 24704 21924 24752 21980
rect 24808 21924 24856 21980
rect 24912 21924 24922 21980
rect 32450 21924 32460 21980
rect 32516 21924 32564 21980
rect 32620 21924 32668 21980
rect 32724 21924 32734 21980
rect 21970 21868 21980 21924
rect 22036 21868 23100 21924
rect 23156 21868 23166 21924
rect 25106 21868 25116 21924
rect 25172 21868 31164 21924
rect 31220 21868 31230 21924
rect 11554 21756 11564 21812
rect 11620 21756 12460 21812
rect 12516 21756 16268 21812
rect 16324 21756 16334 21812
rect 18050 21756 18060 21812
rect 18116 21756 26348 21812
rect 26404 21756 26414 21812
rect 26852 21756 30044 21812
rect 30100 21756 30110 21812
rect 2146 21644 2156 21700
rect 2212 21644 4620 21700
rect 4676 21644 4686 21700
rect 8754 21644 8764 21700
rect 8820 21644 11676 21700
rect 11732 21644 11742 21700
rect 0 21588 800 21616
rect 26852 21588 26908 21756
rect 0 21532 1764 21588
rect 3154 21532 3164 21588
rect 3220 21532 3892 21588
rect 4050 21532 4060 21588
rect 4116 21532 5964 21588
rect 6020 21532 6030 21588
rect 8530 21532 8540 21588
rect 8596 21532 9548 21588
rect 9604 21532 9614 21588
rect 10546 21532 10556 21588
rect 10612 21532 10622 21588
rect 18946 21532 18956 21588
rect 19012 21532 26908 21588
rect 0 21504 800 21532
rect 1708 21252 1764 21532
rect 3836 21476 3892 21532
rect 2594 21420 2604 21476
rect 2660 21420 3388 21476
rect 3836 21420 9100 21476
rect 9156 21420 9166 21476
rect 3332 21364 3388 21420
rect 10556 21364 10612 21532
rect 22194 21420 22204 21476
rect 22260 21420 22764 21476
rect 22820 21420 22830 21476
rect 28242 21420 28252 21476
rect 28308 21420 30044 21476
rect 30100 21420 30110 21476
rect 31490 21420 31500 21476
rect 31556 21420 31836 21476
rect 31892 21420 32172 21476
rect 32228 21420 32238 21476
rect 3332 21308 10612 21364
rect 12562 21308 12572 21364
rect 12628 21308 19516 21364
rect 19572 21308 19582 21364
rect 22642 21308 22652 21364
rect 22708 21308 23548 21364
rect 23604 21308 23614 21364
rect 1698 21196 1708 21252
rect 1764 21196 1774 21252
rect 5108 21140 5118 21196
rect 5174 21140 5222 21196
rect 5278 21140 5326 21196
rect 5382 21140 5392 21196
rect 12920 21140 12930 21196
rect 12986 21140 13034 21196
rect 13090 21140 13138 21196
rect 13194 21140 13204 21196
rect 20732 21140 20742 21196
rect 20798 21140 20846 21196
rect 20902 21140 20950 21196
rect 21006 21140 21016 21196
rect 28544 21140 28554 21196
rect 28610 21140 28658 21196
rect 28714 21140 28762 21196
rect 28818 21140 28828 21196
rect 3332 20972 4620 21028
rect 4676 20972 4686 21028
rect 10882 20972 10892 21028
rect 10948 20972 13804 21028
rect 13860 20972 13870 21028
rect 0 20916 800 20944
rect 0 20860 2156 20916
rect 2212 20860 2222 20916
rect 0 20832 800 20860
rect 3332 20804 3388 20972
rect 4722 20860 4732 20916
rect 4788 20860 6860 20916
rect 6916 20860 6926 20916
rect 13804 20860 17500 20916
rect 17556 20860 17566 20916
rect 21858 20860 21868 20916
rect 21924 20860 26684 20916
rect 26740 20860 26750 20916
rect 13804 20804 13860 20860
rect 2034 20748 2044 20804
rect 2100 20748 3388 20804
rect 4162 20748 4172 20804
rect 4228 20748 9100 20804
rect 9156 20748 9166 20804
rect 12002 20748 12012 20804
rect 12068 20748 13804 20804
rect 13860 20748 13870 20804
rect 14914 20748 14924 20804
rect 14980 20748 15148 20804
rect 15204 20748 19068 20804
rect 19124 20748 22204 20804
rect 22260 20748 22270 20804
rect 3042 20636 3052 20692
rect 3108 20636 8092 20692
rect 8148 20636 8158 20692
rect 12786 20636 12796 20692
rect 12852 20636 17948 20692
rect 18004 20636 18014 20692
rect 25778 20636 25788 20692
rect 25844 20636 26348 20692
rect 26404 20636 26414 20692
rect 29138 20636 29148 20692
rect 29204 20636 30268 20692
rect 30324 20636 30334 20692
rect 26114 20524 26124 20580
rect 26180 20524 31052 20580
rect 31108 20524 31118 20580
rect 9014 20356 9024 20412
rect 9080 20356 9128 20412
rect 9184 20356 9232 20412
rect 9288 20356 9298 20412
rect 16826 20356 16836 20412
rect 16892 20356 16940 20412
rect 16996 20356 17044 20412
rect 17100 20356 17110 20412
rect 24638 20356 24648 20412
rect 24704 20356 24752 20412
rect 24808 20356 24856 20412
rect 24912 20356 24922 20412
rect 32450 20356 32460 20412
rect 32516 20356 32564 20412
rect 32620 20356 32668 20412
rect 32724 20356 32734 20412
rect 0 20244 800 20272
rect 0 20188 4956 20244
rect 5012 20188 5022 20244
rect 23090 20188 23100 20244
rect 23156 20188 23436 20244
rect 23492 20188 23502 20244
rect 28466 20188 28476 20244
rect 28532 20188 31948 20244
rect 32004 20188 32014 20244
rect 0 20160 800 20188
rect 2370 20076 2380 20132
rect 2436 20076 5852 20132
rect 5908 20076 5918 20132
rect 15922 20076 15932 20132
rect 15988 20076 19404 20132
rect 19460 20076 19470 20132
rect 20290 20076 20300 20132
rect 20356 20076 22204 20132
rect 22260 20076 22270 20132
rect 4050 19964 4060 20020
rect 4116 19964 5964 20020
rect 6020 19964 6030 20020
rect 23538 19964 23548 20020
rect 23604 19964 25004 20020
rect 25060 19964 25564 20020
rect 25620 19964 25630 20020
rect 2818 19852 2828 19908
rect 2884 19852 9100 19908
rect 9156 19852 9166 19908
rect 17602 19852 17612 19908
rect 17668 19852 18396 19908
rect 18452 19852 18462 19908
rect 19058 19852 19068 19908
rect 19124 19852 21196 19908
rect 21252 19852 21262 19908
rect 21410 19852 21420 19908
rect 21476 19852 23548 19908
rect 23492 19796 23548 19852
rect 1586 19740 1596 19796
rect 1652 19740 2716 19796
rect 2772 19740 2782 19796
rect 8194 19740 8204 19796
rect 8260 19740 14476 19796
rect 14532 19740 14542 19796
rect 23492 19740 24332 19796
rect 24388 19740 25564 19796
rect 25620 19740 25630 19796
rect 0 19572 800 19600
rect 5108 19572 5118 19628
rect 5174 19572 5222 19628
rect 5278 19572 5326 19628
rect 5382 19572 5392 19628
rect 12920 19572 12930 19628
rect 12986 19572 13034 19628
rect 13090 19572 13138 19628
rect 13194 19572 13204 19628
rect 20732 19572 20742 19628
rect 20798 19572 20846 19628
rect 20902 19572 20950 19628
rect 21006 19572 21016 19628
rect 28544 19572 28554 19628
rect 28610 19572 28658 19628
rect 28714 19572 28762 19628
rect 28818 19572 28828 19628
rect 0 19516 3388 19572
rect 0 19488 800 19516
rect 3332 19460 3388 19516
rect 21420 19516 27356 19572
rect 27412 19516 27422 19572
rect 21420 19460 21476 19516
rect 3332 19404 16716 19460
rect 16772 19404 16782 19460
rect 19170 19404 19180 19460
rect 19236 19404 21476 19460
rect 24882 19404 24892 19460
rect 24948 19404 31500 19460
rect 31556 19404 31566 19460
rect 2034 19292 2044 19348
rect 2100 19292 4508 19348
rect 4564 19292 6412 19348
rect 6468 19292 9772 19348
rect 9828 19292 9838 19348
rect 11218 19292 11228 19348
rect 11284 19292 12908 19348
rect 12964 19292 13692 19348
rect 13748 19292 13758 19348
rect 26852 19292 30156 19348
rect 30212 19292 30222 19348
rect 9772 19236 9828 19292
rect 26852 19236 26908 19292
rect 4050 19180 4060 19236
rect 4116 19180 6076 19236
rect 6132 19180 6142 19236
rect 9772 19180 11452 19236
rect 11508 19180 11518 19236
rect 21858 19180 21868 19236
rect 21924 19180 26908 19236
rect 28690 19180 28700 19236
rect 28756 19180 29484 19236
rect 29540 19180 29550 19236
rect 20738 19068 20748 19124
rect 20804 19068 30940 19124
rect 30996 19068 31006 19124
rect 9014 18788 9024 18844
rect 9080 18788 9128 18844
rect 9184 18788 9232 18844
rect 9288 18788 9298 18844
rect 16826 18788 16836 18844
rect 16892 18788 16940 18844
rect 16996 18788 17044 18844
rect 17100 18788 17110 18844
rect 24638 18788 24648 18844
rect 24704 18788 24752 18844
rect 24808 18788 24856 18844
rect 24912 18788 24922 18844
rect 32450 18788 32460 18844
rect 32516 18788 32564 18844
rect 32620 18788 32668 18844
rect 32724 18788 32734 18844
rect 26852 18620 28140 18676
rect 28196 18620 28206 18676
rect 26852 18564 26908 18620
rect 16594 18508 16604 18564
rect 16660 18508 18060 18564
rect 18116 18508 18396 18564
rect 18452 18508 18462 18564
rect 26674 18508 26684 18564
rect 26740 18508 26908 18564
rect 2930 18396 2940 18452
rect 2996 18396 3500 18452
rect 3556 18396 3566 18452
rect 3714 18396 3724 18452
rect 3780 18396 5628 18452
rect 5684 18396 7644 18452
rect 7700 18396 8988 18452
rect 9044 18396 9054 18452
rect 11442 18396 11452 18452
rect 11508 18396 13020 18452
rect 13076 18396 13086 18452
rect 13906 18396 13916 18452
rect 13972 18396 15148 18452
rect 21186 18396 21196 18452
rect 21252 18396 22428 18452
rect 22484 18396 22494 18452
rect 29138 18396 29148 18452
rect 29204 18396 31276 18452
rect 31332 18396 32060 18452
rect 32116 18396 32126 18452
rect 8988 18340 9044 18396
rect 15092 18340 15148 18396
rect 4946 18284 4956 18340
rect 5012 18284 7868 18340
rect 7924 18284 7934 18340
rect 8988 18284 11676 18340
rect 11732 18284 11742 18340
rect 15092 18284 23212 18340
rect 23268 18284 23278 18340
rect 25554 18284 25564 18340
rect 25620 18284 26124 18340
rect 26180 18284 26460 18340
rect 26516 18284 27132 18340
rect 27188 18284 27198 18340
rect 27570 18284 27580 18340
rect 27636 18284 31948 18340
rect 32004 18284 32014 18340
rect 130 18172 140 18228
rect 196 18172 3388 18228
rect 3490 18172 3500 18228
rect 3556 18172 10836 18228
rect 10994 18172 11004 18228
rect 11060 18172 11788 18228
rect 11844 18172 11854 18228
rect 14354 18172 14364 18228
rect 14420 18172 16940 18228
rect 16996 18172 17006 18228
rect 22082 18172 22092 18228
rect 22148 18172 31164 18228
rect 31220 18172 31230 18228
rect 3332 18116 3388 18172
rect 10780 18116 10836 18172
rect 3332 18060 4956 18116
rect 5012 18060 5022 18116
rect 10780 18060 12012 18116
rect 12068 18060 12078 18116
rect 15092 18060 17612 18116
rect 17668 18060 18172 18116
rect 18228 18060 18238 18116
rect 23314 18060 23324 18116
rect 23380 18060 24556 18116
rect 24612 18060 25452 18116
rect 25508 18060 26572 18116
rect 26628 18060 26638 18116
rect 5108 18004 5118 18060
rect 5174 18004 5222 18060
rect 5278 18004 5326 18060
rect 5382 18004 5392 18060
rect 12920 18004 12930 18060
rect 12986 18004 13034 18060
rect 13090 18004 13138 18060
rect 13194 18004 13204 18060
rect 7410 17948 7420 18004
rect 7476 17948 7756 18004
rect 7812 17948 7822 18004
rect 15092 17892 15148 18060
rect 20732 18004 20742 18060
rect 20798 18004 20846 18060
rect 20902 18004 20950 18060
rect 21006 18004 21016 18060
rect 28544 18004 28554 18060
rect 28610 18004 28658 18060
rect 28714 18004 28762 18060
rect 28818 18004 28828 18060
rect 1932 17836 3052 17892
rect 3108 17836 4508 17892
rect 4564 17836 4574 17892
rect 4834 17836 4844 17892
rect 4900 17836 15148 17892
rect 23324 17836 30492 17892
rect 30548 17836 30558 17892
rect 1932 17556 1988 17836
rect 6962 17724 6972 17780
rect 7028 17724 7420 17780
rect 7476 17724 7644 17780
rect 7700 17724 7710 17780
rect 10210 17724 10220 17780
rect 10276 17724 12124 17780
rect 12180 17724 12190 17780
rect 18498 17724 18508 17780
rect 18564 17724 20748 17780
rect 20804 17724 20814 17780
rect 23324 17668 23380 17836
rect 25778 17724 25788 17780
rect 25844 17724 30156 17780
rect 30212 17724 30222 17780
rect 3938 17612 3948 17668
rect 4004 17612 8204 17668
rect 8260 17612 8270 17668
rect 15362 17612 15372 17668
rect 15428 17612 17164 17668
rect 17220 17612 17230 17668
rect 23314 17612 23324 17668
rect 23380 17612 23390 17668
rect 27122 17612 27132 17668
rect 27188 17612 27356 17668
rect 27412 17612 29260 17668
rect 29316 17612 32060 17668
rect 32116 17612 32126 17668
rect 1922 17500 1932 17556
rect 1988 17500 1998 17556
rect 3042 17500 3052 17556
rect 3108 17500 5404 17556
rect 5460 17500 5470 17556
rect 26338 17500 26348 17556
rect 26404 17500 31164 17556
rect 31220 17500 31230 17556
rect 17602 17388 17612 17444
rect 17668 17388 18732 17444
rect 18788 17388 18798 17444
rect 28578 17388 28588 17444
rect 28644 17388 29596 17444
rect 29652 17388 29662 17444
rect 9014 17220 9024 17276
rect 9080 17220 9128 17276
rect 9184 17220 9232 17276
rect 9288 17220 9298 17276
rect 16826 17220 16836 17276
rect 16892 17220 16940 17276
rect 16996 17220 17044 17276
rect 17100 17220 17110 17276
rect 24638 17220 24648 17276
rect 24704 17220 24752 17276
rect 24808 17220 24856 17276
rect 24912 17220 24922 17276
rect 32450 17220 32460 17276
rect 32516 17220 32564 17276
rect 32620 17220 32668 17276
rect 32724 17220 32734 17276
rect 10994 17164 11004 17220
rect 11060 17164 11564 17220
rect 11620 17164 12348 17220
rect 12404 17164 12908 17220
rect 12964 17164 13580 17220
rect 13636 17164 15484 17220
rect 15540 17164 15550 17220
rect 18946 17164 18956 17220
rect 19012 17164 22540 17220
rect 22596 17164 22606 17220
rect 8642 17052 8652 17108
rect 8708 17052 10668 17108
rect 10724 17052 10734 17108
rect 14354 17052 14364 17108
rect 14420 17052 15148 17108
rect 16370 17052 16380 17108
rect 16436 17052 19404 17108
rect 19460 17052 19470 17108
rect 23650 17052 23660 17108
rect 23716 17052 24332 17108
rect 24388 17052 26124 17108
rect 26180 17052 26190 17108
rect 26898 17052 26908 17108
rect 26964 17052 28028 17108
rect 28084 17052 28094 17108
rect 15092 16996 15148 17052
rect 6178 16940 6188 16996
rect 6244 16940 10892 16996
rect 10948 16940 10958 16996
rect 15092 16940 15260 16996
rect 15316 16940 15326 16996
rect 23314 16940 23324 16996
rect 23380 16940 23996 16996
rect 24052 16940 25900 16996
rect 25956 16940 25966 16996
rect 2818 16828 2828 16884
rect 2884 16828 3500 16884
rect 3556 16828 3566 16884
rect 7074 16828 7084 16884
rect 7140 16828 10332 16884
rect 10388 16828 10398 16884
rect 12562 16828 12572 16884
rect 12628 16828 15932 16884
rect 15988 16828 15998 16884
rect 16818 16828 16828 16884
rect 16884 16828 17500 16884
rect 17556 16828 17566 16884
rect 25330 16828 25340 16884
rect 25396 16828 29260 16884
rect 29316 16828 29326 16884
rect 6066 16716 6076 16772
rect 6132 16716 7756 16772
rect 7812 16716 7822 16772
rect 17826 16716 17836 16772
rect 17892 16716 22988 16772
rect 23044 16716 23054 16772
rect 23986 16716 23996 16772
rect 24052 16716 25564 16772
rect 25620 16716 25630 16772
rect 25778 16716 25788 16772
rect 25844 16716 30044 16772
rect 30100 16716 30110 16772
rect 14914 16604 14924 16660
rect 14980 16604 15820 16660
rect 15876 16604 15886 16660
rect 23090 16604 23100 16660
rect 23156 16604 30156 16660
rect 30212 16604 30222 16660
rect 5108 16436 5118 16492
rect 5174 16436 5222 16492
rect 5278 16436 5326 16492
rect 5382 16436 5392 16492
rect 12920 16436 12930 16492
rect 12986 16436 13034 16492
rect 13090 16436 13138 16492
rect 13194 16436 13204 16492
rect 20732 16436 20742 16492
rect 20798 16436 20846 16492
rect 20902 16436 20950 16492
rect 21006 16436 21016 16492
rect 28544 16436 28554 16492
rect 28610 16436 28658 16492
rect 28714 16436 28762 16492
rect 28818 16436 28828 16492
rect 28914 16380 28924 16436
rect 28980 16380 29372 16436
rect 29428 16380 29438 16436
rect 4722 16156 4732 16212
rect 4788 16156 5068 16212
rect 5124 16156 5964 16212
rect 6020 16156 7420 16212
rect 7476 16156 9772 16212
rect 9828 16156 9838 16212
rect 13010 16156 13020 16212
rect 13076 16156 14812 16212
rect 14868 16156 14878 16212
rect 22642 16156 22652 16212
rect 22708 16156 30156 16212
rect 30212 16156 30222 16212
rect 3938 16044 3948 16100
rect 4004 16044 11228 16100
rect 11284 16044 11294 16100
rect 18610 16044 18620 16100
rect 18676 16044 21420 16100
rect 21476 16044 21980 16100
rect 22036 16044 22046 16100
rect 24658 16044 24668 16100
rect 24724 16044 26908 16100
rect 26964 16044 26974 16100
rect 19618 15932 19628 15988
rect 19684 15932 20300 15988
rect 20356 15932 21308 15988
rect 21364 15932 23212 15988
rect 23268 15932 23278 15988
rect 24882 15932 24892 15988
rect 24948 15932 31164 15988
rect 31220 15932 31230 15988
rect 1250 15820 1260 15876
rect 1316 15820 2268 15876
rect 2324 15820 2334 15876
rect 6402 15820 6412 15876
rect 6468 15820 7308 15876
rect 7364 15820 7374 15876
rect 8978 15820 8988 15876
rect 9044 15820 9884 15876
rect 9940 15820 9950 15876
rect 23538 15820 23548 15876
rect 23604 15820 24108 15876
rect 24164 15820 24174 15876
rect 9014 15652 9024 15708
rect 9080 15652 9128 15708
rect 9184 15652 9232 15708
rect 9288 15652 9298 15708
rect 16826 15652 16836 15708
rect 16892 15652 16940 15708
rect 16996 15652 17044 15708
rect 17100 15652 17110 15708
rect 24638 15652 24648 15708
rect 24704 15652 24752 15708
rect 24808 15652 24856 15708
rect 24912 15652 24922 15708
rect 32450 15652 32460 15708
rect 32516 15652 32564 15708
rect 32620 15652 32668 15708
rect 32724 15652 32734 15708
rect 17714 15596 17724 15652
rect 17780 15596 24332 15652
rect 24388 15596 24398 15652
rect 25666 15596 25676 15652
rect 25732 15596 31052 15652
rect 31108 15596 31118 15652
rect 8978 15484 8988 15540
rect 9044 15484 9772 15540
rect 9828 15484 9838 15540
rect 15138 15484 15148 15540
rect 15204 15484 18284 15540
rect 18340 15484 18350 15540
rect 6626 15372 6636 15428
rect 6692 15372 8204 15428
rect 8260 15372 8270 15428
rect 18162 15372 18172 15428
rect 18228 15372 19628 15428
rect 19684 15372 19694 15428
rect 24658 15372 24668 15428
rect 24724 15372 26012 15428
rect 26068 15372 26078 15428
rect 3154 15260 3164 15316
rect 3220 15260 4620 15316
rect 4676 15260 4686 15316
rect 5618 15260 5628 15316
rect 5684 15260 5964 15316
rect 6020 15260 8540 15316
rect 8596 15260 11116 15316
rect 11172 15260 11182 15316
rect 16594 15148 16604 15204
rect 16660 15148 17500 15204
rect 17556 15148 17566 15204
rect 4722 15036 4732 15092
rect 4788 15036 17052 15092
rect 17108 15036 17118 15092
rect 22082 15036 22092 15092
rect 22148 15036 27916 15092
rect 27972 15036 27982 15092
rect 30706 15036 30716 15092
rect 30772 15036 31612 15092
rect 31668 15036 31678 15092
rect 8642 14924 8652 14980
rect 8708 14924 9660 14980
rect 9716 14924 9726 14980
rect 14690 14924 14700 14980
rect 14756 14924 20412 14980
rect 20468 14924 20478 14980
rect 21858 14924 21868 14980
rect 21924 14924 26796 14980
rect 26852 14924 26862 14980
rect 5108 14868 5118 14924
rect 5174 14868 5222 14924
rect 5278 14868 5326 14924
rect 5382 14868 5392 14924
rect 12920 14868 12930 14924
rect 12986 14868 13034 14924
rect 13090 14868 13138 14924
rect 13194 14868 13204 14924
rect 20732 14868 20742 14924
rect 20798 14868 20846 14924
rect 20902 14868 20950 14924
rect 21006 14868 21016 14924
rect 28544 14868 28554 14924
rect 28610 14868 28658 14924
rect 28714 14868 28762 14924
rect 28818 14868 28828 14924
rect 7970 14812 7980 14868
rect 8036 14812 9884 14868
rect 9940 14812 9950 14868
rect 3042 14700 3052 14756
rect 3108 14700 5628 14756
rect 5684 14700 5694 14756
rect 9426 14700 9436 14756
rect 9492 14700 17388 14756
rect 17444 14700 17454 14756
rect 4386 14588 4396 14644
rect 4452 14588 4732 14644
rect 4788 14588 4798 14644
rect 12450 14588 12460 14644
rect 12516 14588 16380 14644
rect 16436 14588 16446 14644
rect 24546 14588 24556 14644
rect 24612 14588 30156 14644
rect 30212 14588 30222 14644
rect 2482 14476 2492 14532
rect 2548 14476 3388 14532
rect 3714 14476 3724 14532
rect 3780 14476 8540 14532
rect 8596 14476 8606 14532
rect 9202 14476 9212 14532
rect 9268 14476 9996 14532
rect 10052 14476 12348 14532
rect 12404 14476 12414 14532
rect 3332 14420 3388 14476
rect 1586 14364 1596 14420
rect 1652 14364 2716 14420
rect 2772 14364 2782 14420
rect 3332 14364 20748 14420
rect 20804 14364 20814 14420
rect 21746 14364 21756 14420
rect 21812 14364 27244 14420
rect 27300 14364 27310 14420
rect 4610 14252 4620 14308
rect 4676 14252 4956 14308
rect 5012 14252 5022 14308
rect 10882 14252 10892 14308
rect 10948 14252 13020 14308
rect 13076 14252 13086 14308
rect 19170 14252 19180 14308
rect 19236 14252 20524 14308
rect 20580 14252 20590 14308
rect 29586 14252 29596 14308
rect 29652 14252 29820 14308
rect 29876 14252 30716 14308
rect 30772 14252 32060 14308
rect 32116 14252 32126 14308
rect 29362 14140 29372 14196
rect 29428 14140 30380 14196
rect 30436 14140 30446 14196
rect 9014 14084 9024 14140
rect 9080 14084 9128 14140
rect 9184 14084 9232 14140
rect 9288 14084 9298 14140
rect 16826 14084 16836 14140
rect 16892 14084 16940 14140
rect 16996 14084 17044 14140
rect 17100 14084 17110 14140
rect 24638 14084 24648 14140
rect 24704 14084 24752 14140
rect 24808 14084 24856 14140
rect 24912 14084 24922 14140
rect 32450 14084 32460 14140
rect 32516 14084 32564 14140
rect 32620 14084 32668 14140
rect 32724 14084 32734 14140
rect 4386 14028 4396 14084
rect 4452 14028 7252 14084
rect 28130 14028 28140 14084
rect 28196 14028 30156 14084
rect 30212 14028 30222 14084
rect 7196 13972 7252 14028
rect 2370 13916 2380 13972
rect 2436 13916 5740 13972
rect 5796 13916 5806 13972
rect 7196 13916 18060 13972
rect 18116 13916 18126 13972
rect 3332 13804 5404 13860
rect 5460 13804 5470 13860
rect 20738 13804 20748 13860
rect 20804 13804 21420 13860
rect 21476 13804 21486 13860
rect 3332 13524 3388 13804
rect 11890 13692 11900 13748
rect 11956 13692 13692 13748
rect 13748 13692 13758 13748
rect 14466 13692 14476 13748
rect 14532 13692 15260 13748
rect 15316 13692 16156 13748
rect 16212 13692 16604 13748
rect 16660 13692 16670 13748
rect 19058 13692 19068 13748
rect 19124 13692 22876 13748
rect 22932 13692 22942 13748
rect 4722 13580 4732 13636
rect 4788 13580 8652 13636
rect 8708 13580 8718 13636
rect 10098 13580 10108 13636
rect 10164 13580 11676 13636
rect 11732 13580 12796 13636
rect 12852 13580 12862 13636
rect 18274 13580 18284 13636
rect 18340 13580 18956 13636
rect 19012 13580 19022 13636
rect 22530 13580 22540 13636
rect 22596 13580 24668 13636
rect 24724 13580 25676 13636
rect 25732 13580 25742 13636
rect 26338 13580 26348 13636
rect 26404 13580 31276 13636
rect 31332 13580 31342 13636
rect 25676 13524 25732 13580
rect 3042 13468 3052 13524
rect 3108 13468 3388 13524
rect 5282 13468 5292 13524
rect 5348 13468 6804 13524
rect 25676 13468 27748 13524
rect 6748 13412 6804 13468
rect 27692 13412 27748 13468
rect 6748 13356 7420 13412
rect 7476 13356 7486 13412
rect 27692 13356 27804 13412
rect 27860 13356 27870 13412
rect 5108 13300 5118 13356
rect 5174 13300 5222 13356
rect 5278 13300 5326 13356
rect 5382 13300 5392 13356
rect 12920 13300 12930 13356
rect 12986 13300 13034 13356
rect 13090 13300 13138 13356
rect 13194 13300 13204 13356
rect 20732 13300 20742 13356
rect 20798 13300 20846 13356
rect 20902 13300 20950 13356
rect 21006 13300 21016 13356
rect 28544 13300 28554 13356
rect 28610 13300 28658 13356
rect 28714 13300 28762 13356
rect 28818 13300 28828 13356
rect 13682 13244 13692 13300
rect 13748 13244 15372 13300
rect 15428 13244 16492 13300
rect 16548 13244 16558 13300
rect 2034 13132 2044 13188
rect 2100 13132 17724 13188
rect 17780 13132 17790 13188
rect 21858 13132 21868 13188
rect 21924 13132 26460 13188
rect 26516 13132 26526 13188
rect 3826 13020 3836 13076
rect 3892 13020 4508 13076
rect 4564 13020 4574 13076
rect 4834 13020 4844 13076
rect 4900 13020 8092 13076
rect 8148 13020 8158 13076
rect 12450 13020 12460 13076
rect 12516 13020 13580 13076
rect 13636 13020 13646 13076
rect 17602 13020 17612 13076
rect 17668 13020 19292 13076
rect 19348 13020 19358 13076
rect 1698 12908 1708 12964
rect 1764 12908 2940 12964
rect 2996 12908 3006 12964
rect 6738 12908 6748 12964
rect 6804 12908 14588 12964
rect 14644 12908 14654 12964
rect 4946 12796 4956 12852
rect 5012 12796 12012 12852
rect 12068 12796 12078 12852
rect 12898 12684 12908 12740
rect 12964 12684 13692 12740
rect 13748 12684 13758 12740
rect 9014 12516 9024 12572
rect 9080 12516 9128 12572
rect 9184 12516 9232 12572
rect 9288 12516 9298 12572
rect 16826 12516 16836 12572
rect 16892 12516 16940 12572
rect 16996 12516 17044 12572
rect 17100 12516 17110 12572
rect 24638 12516 24648 12572
rect 24704 12516 24752 12572
rect 24808 12516 24856 12572
rect 24912 12516 24922 12572
rect 32450 12516 32460 12572
rect 32516 12516 32564 12572
rect 32620 12516 32668 12572
rect 32724 12516 32734 12572
rect 4050 12460 4060 12516
rect 4116 12460 8428 12516
rect 8484 12460 8494 12516
rect 2482 12348 2492 12404
rect 2548 12348 3276 12404
rect 3332 12348 3342 12404
rect 4386 12348 4396 12404
rect 4452 12348 5516 12404
rect 5572 12348 5582 12404
rect 7410 12348 7420 12404
rect 7476 12348 8988 12404
rect 9044 12348 9996 12404
rect 10052 12348 10062 12404
rect 7522 12236 7532 12292
rect 7588 12236 17388 12292
rect 17444 12236 17454 12292
rect 20178 12236 20188 12292
rect 20244 12236 23884 12292
rect 23940 12236 23950 12292
rect 11666 12124 11676 12180
rect 11732 12124 14364 12180
rect 14420 12124 15148 12180
rect 15204 12124 15214 12180
rect 27794 12124 27804 12180
rect 27860 12124 29148 12180
rect 29204 12124 29820 12180
rect 29876 12124 29886 12180
rect 4162 12012 4172 12068
rect 4228 12012 14924 12068
rect 14980 12012 16492 12068
rect 16548 12012 16558 12068
rect 6178 11900 6188 11956
rect 6244 11900 15260 11956
rect 15316 11900 15326 11956
rect 5108 11732 5118 11788
rect 5174 11732 5222 11788
rect 5278 11732 5326 11788
rect 5382 11732 5392 11788
rect 12920 11732 12930 11788
rect 12986 11732 13034 11788
rect 13090 11732 13138 11788
rect 13194 11732 13204 11788
rect 20732 11732 20742 11788
rect 20798 11732 20846 11788
rect 20902 11732 20950 11788
rect 21006 11732 21016 11788
rect 28544 11732 28554 11788
rect 28610 11732 28658 11788
rect 28714 11732 28762 11788
rect 28818 11732 28828 11788
rect 15092 11676 15372 11732
rect 15428 11676 18508 11732
rect 18564 11676 18574 11732
rect 21746 11676 21756 11732
rect 21812 11676 21822 11732
rect 2370 11564 2380 11620
rect 2436 11564 5740 11620
rect 5796 11564 5806 11620
rect 2258 11452 2268 11508
rect 2324 11452 3556 11508
rect 3500 11396 3556 11452
rect 3836 11452 14700 11508
rect 14756 11452 14766 11508
rect 3836 11396 3892 11452
rect 15092 11396 15148 11676
rect 21756 11508 21812 11676
rect 19170 11452 19180 11508
rect 19236 11452 21812 11508
rect 25218 11452 25228 11508
rect 25284 11452 26348 11508
rect 26404 11452 29260 11508
rect 29316 11452 29820 11508
rect 29876 11452 32060 11508
rect 32116 11452 32126 11508
rect 1922 11340 1932 11396
rect 1988 11340 3388 11396
rect 3500 11340 3892 11396
rect 4134 11340 4172 11396
rect 4228 11340 4238 11396
rect 9426 11340 9436 11396
rect 9492 11340 10892 11396
rect 10948 11340 12908 11396
rect 12964 11340 15148 11396
rect 18162 11340 18172 11396
rect 18228 11340 21196 11396
rect 21252 11340 21262 11396
rect 3332 11284 3388 11340
rect 3332 11228 4508 11284
rect 4564 11228 4574 11284
rect 21074 11228 21084 11284
rect 21140 11228 24388 11284
rect 25106 11228 25116 11284
rect 25172 11228 31164 11284
rect 31220 11228 31230 11284
rect 24332 11172 24388 11228
rect 13458 11116 13468 11172
rect 13524 11116 19180 11172
rect 19236 11116 19246 11172
rect 23090 11116 23100 11172
rect 23156 11116 24108 11172
rect 24164 11116 24174 11172
rect 24332 11116 30268 11172
rect 30324 11116 30334 11172
rect 26786 11004 26796 11060
rect 26852 11004 30156 11060
rect 30212 11004 30222 11060
rect 9014 10948 9024 11004
rect 9080 10948 9128 11004
rect 9184 10948 9232 11004
rect 9288 10948 9298 11004
rect 16826 10948 16836 11004
rect 16892 10948 16940 11004
rect 16996 10948 17044 11004
rect 17100 10948 17110 11004
rect 24638 10948 24648 11004
rect 24704 10948 24752 11004
rect 24808 10948 24856 11004
rect 24912 10948 24922 11004
rect 32450 10948 32460 11004
rect 32516 10948 32564 11004
rect 32620 10948 32668 11004
rect 32724 10948 32734 11004
rect 1932 10892 2604 10948
rect 2660 10892 2670 10948
rect 1932 10500 1988 10892
rect 4946 10780 4956 10836
rect 5012 10780 8428 10836
rect 8484 10780 10108 10836
rect 10164 10780 10174 10836
rect 10546 10780 10556 10836
rect 10612 10780 11676 10836
rect 11732 10780 11742 10836
rect 28242 10780 28252 10836
rect 28308 10780 30156 10836
rect 30212 10780 30222 10836
rect 10556 10724 10612 10780
rect 5954 10668 5964 10724
rect 6020 10668 6636 10724
rect 6692 10668 7308 10724
rect 7364 10668 8316 10724
rect 8372 10668 10612 10724
rect 19058 10668 19068 10724
rect 19124 10668 20972 10724
rect 21028 10668 21038 10724
rect 21634 10668 21644 10724
rect 21700 10668 23884 10724
rect 23940 10668 23950 10724
rect 29922 10668 29932 10724
rect 29988 10668 30604 10724
rect 30660 10668 32284 10724
rect 32340 10668 32350 10724
rect 18162 10556 18172 10612
rect 18228 10556 19404 10612
rect 19460 10556 20188 10612
rect 24434 10556 24444 10612
rect 24500 10556 30940 10612
rect 30996 10556 31006 10612
rect 20132 10500 20188 10556
rect 1922 10444 1932 10500
rect 1988 10444 1998 10500
rect 4498 10444 4508 10500
rect 4564 10444 15260 10500
rect 15316 10444 15326 10500
rect 20132 10444 20524 10500
rect 20580 10444 21868 10500
rect 21924 10444 21934 10500
rect 3042 10332 3052 10388
rect 3108 10332 5292 10388
rect 5348 10332 5358 10388
rect 10882 10332 10892 10388
rect 10948 10332 13468 10388
rect 13524 10332 13534 10388
rect 5108 10164 5118 10220
rect 5174 10164 5222 10220
rect 5278 10164 5326 10220
rect 5382 10164 5392 10220
rect 12920 10164 12930 10220
rect 12986 10164 13034 10220
rect 13090 10164 13138 10220
rect 13194 10164 13204 10220
rect 20732 10164 20742 10220
rect 20798 10164 20846 10220
rect 20902 10164 20950 10220
rect 21006 10164 21016 10220
rect 28544 10164 28554 10220
rect 28610 10164 28658 10220
rect 28714 10164 28762 10220
rect 28818 10164 28828 10220
rect 30034 10108 30044 10164
rect 30100 10108 30110 10164
rect 30044 10052 30100 10108
rect 1474 9996 1484 10052
rect 1540 9996 2716 10052
rect 2772 9996 2782 10052
rect 21522 9996 21532 10052
rect 21588 9996 25508 10052
rect 28354 9996 28364 10052
rect 28420 9996 29148 10052
rect 29204 9996 29214 10052
rect 30044 9996 32172 10052
rect 32228 9996 32238 10052
rect 25452 9828 25508 9996
rect 25666 9884 25676 9940
rect 25732 9884 30044 9940
rect 30100 9884 30110 9940
rect 8306 9772 8316 9828
rect 8372 9772 10892 9828
rect 10948 9772 10958 9828
rect 11330 9772 11340 9828
rect 11396 9772 18956 9828
rect 19012 9772 19404 9828
rect 19460 9772 19470 9828
rect 20738 9772 20748 9828
rect 20804 9772 21532 9828
rect 21588 9772 21598 9828
rect 25452 9772 31724 9828
rect 31780 9772 31790 9828
rect 3826 9660 3836 9716
rect 3892 9660 14028 9716
rect 14084 9660 14812 9716
rect 14868 9660 14878 9716
rect 24994 9660 25004 9716
rect 25060 9660 31164 9716
rect 31220 9660 31230 9716
rect 1810 9548 1820 9604
rect 1876 9548 4620 9604
rect 4676 9548 4686 9604
rect 5058 9548 5068 9604
rect 5124 9548 5964 9604
rect 6020 9548 6030 9604
rect 6626 9548 6636 9604
rect 6692 9548 8316 9604
rect 8372 9548 8382 9604
rect 12450 9548 12460 9604
rect 12516 9548 13580 9604
rect 13636 9548 13646 9604
rect 17714 9548 17724 9604
rect 17780 9548 19180 9604
rect 19236 9548 19246 9604
rect 21634 9548 21644 9604
rect 21700 9548 25564 9604
rect 25620 9548 25630 9604
rect 25778 9548 25788 9604
rect 25844 9548 27468 9604
rect 27524 9548 27534 9604
rect 27346 9436 27356 9492
rect 27412 9436 28588 9492
rect 28644 9436 28654 9492
rect 9014 9380 9024 9436
rect 9080 9380 9128 9436
rect 9184 9380 9232 9436
rect 9288 9380 9298 9436
rect 16826 9380 16836 9436
rect 16892 9380 16940 9436
rect 16996 9380 17044 9436
rect 17100 9380 17110 9436
rect 24638 9380 24648 9436
rect 24704 9380 24752 9436
rect 24808 9380 24856 9436
rect 24912 9380 24922 9436
rect 32450 9380 32460 9436
rect 32516 9380 32564 9436
rect 32620 9380 32668 9436
rect 32724 9380 32734 9436
rect 2034 9324 2044 9380
rect 2100 9324 5852 9380
rect 5908 9324 5918 9380
rect 10770 9324 10780 9380
rect 10836 9324 16268 9380
rect 16324 9324 16334 9380
rect 3938 9212 3948 9268
rect 4004 9212 5516 9268
rect 5572 9212 5582 9268
rect 10434 9212 10444 9268
rect 10500 9212 11228 9268
rect 11284 9212 13468 9268
rect 13524 9212 14252 9268
rect 14308 9212 14318 9268
rect 21522 9212 21532 9268
rect 21588 9212 22316 9268
rect 22372 9212 22876 9268
rect 22932 9212 25228 9268
rect 25284 9212 25294 9268
rect 1922 9100 1932 9156
rect 1988 9100 9548 9156
rect 9604 9100 9614 9156
rect 14802 9100 14812 9156
rect 14868 9100 16156 9156
rect 16212 9100 16222 9156
rect 24210 9100 24220 9156
rect 24276 9100 24286 9156
rect 8530 8988 8540 9044
rect 8596 8988 15484 9044
rect 15540 8988 15550 9044
rect 18946 8988 18956 9044
rect 19012 8988 19022 9044
rect 19170 8988 19180 9044
rect 19236 8988 21420 9044
rect 21476 8988 21486 9044
rect 18956 8932 19012 8988
rect 24220 8932 24276 9100
rect 10658 8876 10668 8932
rect 10724 8876 13244 8932
rect 13300 8876 13310 8932
rect 13794 8876 13804 8932
rect 13860 8876 16492 8932
rect 16548 8876 16558 8932
rect 18956 8876 23212 8932
rect 23268 8876 23278 8932
rect 23436 8876 24276 8932
rect 13244 8820 13300 8876
rect 23436 8820 23492 8876
rect 1810 8764 1820 8820
rect 1876 8764 2828 8820
rect 2884 8764 2894 8820
rect 13244 8764 15148 8820
rect 19282 8764 19292 8820
rect 19348 8764 23492 8820
rect 24322 8764 24332 8820
rect 24388 8764 25340 8820
rect 25396 8764 25406 8820
rect 28130 8764 28140 8820
rect 28196 8764 30156 8820
rect 30212 8764 30222 8820
rect 5108 8596 5118 8652
rect 5174 8596 5222 8652
rect 5278 8596 5326 8652
rect 5382 8596 5392 8652
rect 12920 8596 12930 8652
rect 12986 8596 13034 8652
rect 13090 8596 13138 8652
rect 13194 8596 13204 8652
rect 15092 8484 15148 8764
rect 22978 8652 22988 8708
rect 23044 8652 26348 8708
rect 26404 8652 27356 8708
rect 27412 8652 27422 8708
rect 20732 8596 20742 8652
rect 20798 8596 20846 8652
rect 20902 8596 20950 8652
rect 21006 8596 21016 8652
rect 28544 8596 28554 8652
rect 28610 8596 28658 8652
rect 28714 8596 28762 8652
rect 28818 8596 28828 8652
rect 15092 8428 15260 8484
rect 15316 8428 15820 8484
rect 15876 8428 15886 8484
rect 28018 8428 28028 8484
rect 28084 8428 28700 8484
rect 28756 8428 29708 8484
rect 29764 8428 29774 8484
rect 1586 8316 1596 8372
rect 1652 8316 3276 8372
rect 3332 8316 3342 8372
rect 14242 8316 14252 8372
rect 14308 8316 15036 8372
rect 15092 8316 15102 8372
rect 8754 8204 8764 8260
rect 8820 8204 17500 8260
rect 17556 8204 17566 8260
rect 18386 8204 18396 8260
rect 18452 8204 21196 8260
rect 21252 8204 23548 8260
rect 23604 8204 23614 8260
rect 9090 8092 9100 8148
rect 9156 8092 12236 8148
rect 12292 8092 12302 8148
rect 16930 8092 16940 8148
rect 16996 8092 19404 8148
rect 19460 8092 19470 8148
rect 27122 8092 27132 8148
rect 27188 8092 31164 8148
rect 31220 8092 31230 8148
rect 33200 8064 34000 8176
rect 8642 7980 8652 8036
rect 8708 7980 20524 8036
rect 20580 7980 20590 8036
rect 25890 7980 25900 8036
rect 25956 7980 29260 8036
rect 29316 7980 29326 8036
rect 9762 7868 9772 7924
rect 9828 7868 9838 7924
rect 9986 7868 9996 7924
rect 10052 7868 11228 7924
rect 11284 7868 11294 7924
rect 9014 7812 9024 7868
rect 9080 7812 9128 7868
rect 9184 7812 9232 7868
rect 9288 7812 9298 7868
rect 9772 7700 9828 7868
rect 16826 7812 16836 7868
rect 16892 7812 16940 7868
rect 16996 7812 17044 7868
rect 17100 7812 17110 7868
rect 24638 7812 24648 7868
rect 24704 7812 24752 7868
rect 24808 7812 24856 7868
rect 24912 7812 24922 7868
rect 32450 7812 32460 7868
rect 32516 7812 32564 7868
rect 32620 7812 32668 7868
rect 32724 7812 32734 7868
rect 28354 7756 28364 7812
rect 28420 7756 30156 7812
rect 30212 7756 30222 7812
rect 2034 7644 2044 7700
rect 2100 7644 9828 7700
rect 15810 7644 15820 7700
rect 15876 7644 16828 7700
rect 16884 7644 17948 7700
rect 18004 7644 20748 7700
rect 20804 7644 20814 7700
rect 15922 7532 15932 7588
rect 15988 7532 26292 7588
rect 15026 7420 15036 7476
rect 15092 7420 17500 7476
rect 17556 7420 17566 7476
rect 18722 7420 18732 7476
rect 18788 7420 24332 7476
rect 24388 7420 24398 7476
rect 26236 7364 26292 7532
rect 33200 7476 34000 7504
rect 31826 7420 31836 7476
rect 31892 7420 34000 7476
rect 33200 7392 34000 7420
rect 3490 7308 3500 7364
rect 3556 7308 6748 7364
rect 6804 7308 6814 7364
rect 16258 7308 16268 7364
rect 16324 7308 18396 7364
rect 18452 7308 18462 7364
rect 21970 7308 21980 7364
rect 22036 7308 24108 7364
rect 24164 7308 24174 7364
rect 26226 7308 26236 7364
rect 26292 7308 26302 7364
rect 5394 7196 5404 7252
rect 5460 7196 6636 7252
rect 6692 7196 6702 7252
rect 16706 7196 16716 7252
rect 16772 7196 20076 7252
rect 20132 7196 20142 7252
rect 14018 7084 14028 7140
rect 14084 7084 15372 7140
rect 15428 7084 15438 7140
rect 5108 7028 5118 7084
rect 5174 7028 5222 7084
rect 5278 7028 5326 7084
rect 5382 7028 5392 7084
rect 12920 7028 12930 7084
rect 12986 7028 13034 7084
rect 13090 7028 13138 7084
rect 13194 7028 13204 7084
rect 20732 7028 20742 7084
rect 20798 7028 20846 7084
rect 20902 7028 20950 7084
rect 21006 7028 21016 7084
rect 28544 7028 28554 7084
rect 28610 7028 28658 7084
rect 28714 7028 28762 7084
rect 28818 7028 28828 7084
rect 4610 6860 4620 6916
rect 4676 6860 11340 6916
rect 11396 6860 11406 6916
rect 28466 6860 28476 6916
rect 28532 6860 29036 6916
rect 29092 6860 29102 6916
rect 0 6804 800 6832
rect 33200 6804 34000 6832
rect 0 6748 3836 6804
rect 3892 6748 3902 6804
rect 5058 6748 5068 6804
rect 5124 6748 5404 6804
rect 5460 6748 6300 6804
rect 6356 6748 7588 6804
rect 17826 6748 17836 6804
rect 17892 6748 19180 6804
rect 19236 6748 19246 6804
rect 21970 6748 21980 6804
rect 22036 6748 23100 6804
rect 23156 6748 23166 6804
rect 23986 6748 23996 6804
rect 24052 6748 25900 6804
rect 25956 6748 25966 6804
rect 28588 6748 34000 6804
rect 0 6720 800 6748
rect 7532 6692 7588 6748
rect 3378 6636 3388 6692
rect 3444 6636 3482 6692
rect 4050 6636 4060 6692
rect 4116 6636 6860 6692
rect 6916 6636 6926 6692
rect 7522 6636 7532 6692
rect 7588 6636 7598 6692
rect 10322 6636 10332 6692
rect 10388 6636 10780 6692
rect 10836 6636 11676 6692
rect 11732 6636 11742 6692
rect 16034 6636 16044 6692
rect 16100 6636 18844 6692
rect 18900 6636 19516 6692
rect 19572 6636 20300 6692
rect 20356 6636 20366 6692
rect 3602 6524 3612 6580
rect 3668 6524 5628 6580
rect 5684 6524 5694 6580
rect 10658 6524 10668 6580
rect 10724 6524 14700 6580
rect 14756 6524 14766 6580
rect 15026 6524 15036 6580
rect 15092 6524 16380 6580
rect 16436 6524 16446 6580
rect 18162 6524 18172 6580
rect 18228 6524 20188 6580
rect 20244 6524 20254 6580
rect 21522 6524 21532 6580
rect 21588 6524 22316 6580
rect 22372 6524 22382 6580
rect 25106 6524 25116 6580
rect 25172 6524 26908 6580
rect 26964 6524 26974 6580
rect 28588 6468 28644 6748
rect 33200 6720 34000 6748
rect 29362 6636 29372 6692
rect 29428 6636 31164 6692
rect 31220 6636 31230 6692
rect 1250 6412 1260 6468
rect 1316 6412 9772 6468
rect 9828 6412 9838 6468
rect 15138 6412 15148 6468
rect 15204 6412 16044 6468
rect 16100 6412 16110 6468
rect 17490 6412 17500 6468
rect 17556 6412 18284 6468
rect 18340 6412 28644 6468
rect 3042 6300 3052 6356
rect 3108 6300 4060 6356
rect 4116 6300 4126 6356
rect 17826 6300 17836 6356
rect 17892 6300 18620 6356
rect 18676 6300 18686 6356
rect 9014 6244 9024 6300
rect 9080 6244 9128 6300
rect 9184 6244 9232 6300
rect 9288 6244 9298 6300
rect 16826 6244 16836 6300
rect 16892 6244 16940 6300
rect 16996 6244 17044 6300
rect 17100 6244 17110 6300
rect 24638 6244 24648 6300
rect 24704 6244 24752 6300
rect 24808 6244 24856 6300
rect 24912 6244 24922 6300
rect 32450 6244 32460 6300
rect 32516 6244 32564 6300
rect 32620 6244 32668 6300
rect 32724 6244 32734 6300
rect 1810 6188 1820 6244
rect 1876 6188 4172 6244
rect 4228 6188 4508 6244
rect 4564 6188 4574 6244
rect 0 6132 800 6160
rect 33200 6132 34000 6160
rect 0 6076 3388 6132
rect 7410 6076 7420 6132
rect 7476 6076 8092 6132
rect 8148 6076 8158 6132
rect 9538 6076 9548 6132
rect 9604 6076 10444 6132
rect 10500 6076 10510 6132
rect 27346 6076 27356 6132
rect 27412 6076 34000 6132
rect 0 6048 800 6076
rect 3332 6020 3388 6076
rect 33200 6048 34000 6076
rect 3332 5964 13468 6020
rect 13524 5964 14476 6020
rect 14532 5964 14542 6020
rect 16146 5964 16156 6020
rect 16212 5964 17388 6020
rect 17444 5964 17454 6020
rect 20962 5964 20972 6020
rect 21028 5964 22316 6020
rect 22372 5964 22382 6020
rect 24994 5964 25004 6020
rect 25060 5964 25788 6020
rect 25844 5964 25854 6020
rect 2258 5852 2268 5908
rect 2324 5852 5628 5908
rect 5684 5852 5694 5908
rect 7186 5852 7196 5908
rect 7252 5852 7262 5908
rect 7522 5852 7532 5908
rect 7588 5852 8316 5908
rect 8372 5852 8382 5908
rect 13906 5852 13916 5908
rect 13972 5852 15148 5908
rect 15204 5852 15214 5908
rect 29922 5852 29932 5908
rect 29988 5852 31052 5908
rect 31108 5852 31118 5908
rect 7196 5796 7252 5852
rect 3378 5740 3388 5796
rect 3444 5740 3948 5796
rect 4004 5740 4014 5796
rect 4834 5740 4844 5796
rect 4900 5740 6356 5796
rect 7196 5740 18060 5796
rect 18116 5740 18126 5796
rect 6300 5684 6356 5740
rect 3826 5628 3836 5684
rect 3892 5628 6076 5684
rect 6132 5628 6142 5684
rect 6300 5628 21308 5684
rect 21364 5628 21374 5684
rect 22418 5628 22428 5684
rect 22484 5628 29036 5684
rect 29092 5628 29102 5684
rect 7186 5516 7196 5572
rect 7252 5516 8092 5572
rect 8148 5516 8158 5572
rect 0 5460 800 5488
rect 5108 5460 5118 5516
rect 5174 5460 5222 5516
rect 5278 5460 5326 5516
rect 5382 5460 5392 5516
rect 12920 5460 12930 5516
rect 12986 5460 13034 5516
rect 13090 5460 13138 5516
rect 13194 5460 13204 5516
rect 20732 5460 20742 5516
rect 20798 5460 20846 5516
rect 20902 5460 20950 5516
rect 21006 5460 21016 5516
rect 28544 5460 28554 5516
rect 28610 5460 28658 5516
rect 28714 5460 28762 5516
rect 28818 5460 28828 5516
rect 33200 5460 34000 5488
rect 0 5404 1932 5460
rect 1988 5404 1998 5460
rect 6402 5404 6412 5460
rect 6468 5404 12572 5460
rect 12628 5404 12638 5460
rect 21746 5404 21756 5460
rect 21812 5404 26236 5460
rect 26292 5404 26302 5460
rect 31892 5404 34000 5460
rect 0 5376 800 5404
rect 31892 5348 31948 5404
rect 33200 5376 34000 5404
rect 2930 5292 2940 5348
rect 2996 5292 3388 5348
rect 9426 5292 9436 5348
rect 9492 5292 20300 5348
rect 20356 5292 20366 5348
rect 21186 5292 21196 5348
rect 21252 5292 21980 5348
rect 22036 5292 22046 5348
rect 23762 5292 23772 5348
rect 23828 5292 31948 5348
rect 3332 5236 3388 5292
rect 3332 5180 17164 5236
rect 17220 5180 17230 5236
rect 20402 5180 20412 5236
rect 20468 5180 24332 5236
rect 24388 5180 25620 5236
rect 27570 5180 27580 5236
rect 27636 5180 31388 5236
rect 31444 5180 31454 5236
rect 25564 5124 25620 5180
rect 3332 5068 10108 5124
rect 10164 5068 10174 5124
rect 12562 5068 12572 5124
rect 12628 5068 13916 5124
rect 13972 5068 13982 5124
rect 17266 5068 17276 5124
rect 17332 5068 17724 5124
rect 17780 5068 19852 5124
rect 19908 5068 22092 5124
rect 22148 5068 22540 5124
rect 22596 5068 24668 5124
rect 24724 5068 24734 5124
rect 25564 5068 30044 5124
rect 30100 5068 30110 5124
rect 0 4788 800 4816
rect 3332 4788 3388 5068
rect 6290 4956 6300 5012
rect 6356 4956 8764 5012
rect 8820 4956 8830 5012
rect 16594 4956 16604 5012
rect 16660 4956 17164 5012
rect 17220 4956 26124 5012
rect 26180 4956 26190 5012
rect 26562 4956 26572 5012
rect 26628 4956 28140 5012
rect 28196 4956 28206 5012
rect 5058 4844 5068 4900
rect 5124 4844 6748 4900
rect 6804 4844 6814 4900
rect 8194 4844 8204 4900
rect 8260 4844 10108 4900
rect 10164 4844 10174 4900
rect 14130 4844 14140 4900
rect 14196 4844 15484 4900
rect 15540 4844 15550 4900
rect 20738 4844 20748 4900
rect 20804 4844 22764 4900
rect 22820 4844 22830 4900
rect 25330 4844 25340 4900
rect 25396 4844 32900 4900
rect 32844 4788 32900 4844
rect 33200 4788 34000 4816
rect 0 4732 3388 4788
rect 5730 4732 5740 4788
rect 5796 4732 7532 4788
rect 7588 4732 7598 4788
rect 27122 4732 27132 4788
rect 27188 4732 31164 4788
rect 31220 4732 31230 4788
rect 32844 4732 34000 4788
rect 0 4704 800 4732
rect 9014 4676 9024 4732
rect 9080 4676 9128 4732
rect 9184 4676 9232 4732
rect 9288 4676 9298 4732
rect 16826 4676 16836 4732
rect 16892 4676 16940 4732
rect 16996 4676 17044 4732
rect 17100 4676 17110 4732
rect 24638 4676 24648 4732
rect 24704 4676 24752 4732
rect 24808 4676 24856 4732
rect 24912 4676 24922 4732
rect 32450 4676 32460 4732
rect 32516 4676 32564 4732
rect 32620 4676 32668 4732
rect 32724 4676 32734 4732
rect 33200 4704 34000 4732
rect 9436 4620 14588 4676
rect 14644 4620 14654 4676
rect 9436 4564 9492 4620
rect 4722 4508 4732 4564
rect 4788 4508 9492 4564
rect 9650 4508 9660 4564
rect 9716 4508 18956 4564
rect 19012 4508 19022 4564
rect 26786 4508 26796 4564
rect 26852 4508 27468 4564
rect 27524 4508 27534 4564
rect 27682 4508 27692 4564
rect 27748 4508 28700 4564
rect 28756 4508 28766 4564
rect 4610 4396 4620 4452
rect 4676 4396 5740 4452
rect 5796 4396 5806 4452
rect 16258 4396 16268 4452
rect 16324 4396 19404 4452
rect 19460 4396 19470 4452
rect 20132 4396 28980 4452
rect 20132 4340 20188 4396
rect 12786 4284 12796 4340
rect 12852 4284 14700 4340
rect 14756 4284 14766 4340
rect 18498 4284 18508 4340
rect 18564 4284 20188 4340
rect 20290 4284 20300 4340
rect 20356 4284 23548 4340
rect 23604 4284 23614 4340
rect 15138 4172 15148 4228
rect 15204 4172 18396 4228
rect 18452 4172 18462 4228
rect 20178 4172 20188 4228
rect 20244 4172 21308 4228
rect 21364 4172 24108 4228
rect 24164 4172 24668 4228
rect 24724 4172 24734 4228
rect 0 4116 800 4144
rect 0 4060 4172 4116
rect 4228 4060 4238 4116
rect 13234 4060 13244 4116
rect 13300 4060 14812 4116
rect 14868 4060 14878 4116
rect 24210 4060 24220 4116
rect 24276 4060 27580 4116
rect 27636 4060 27646 4116
rect 0 4032 800 4060
rect 15092 3948 19628 4004
rect 19684 3948 19694 4004
rect 5108 3892 5118 3948
rect 5174 3892 5222 3948
rect 5278 3892 5326 3948
rect 5382 3892 5392 3948
rect 12920 3892 12930 3948
rect 12986 3892 13034 3948
rect 13090 3892 13138 3948
rect 13194 3892 13204 3948
rect 15092 3780 15148 3948
rect 20732 3892 20742 3948
rect 20798 3892 20846 3948
rect 20902 3892 20950 3948
rect 21006 3892 21016 3948
rect 28544 3892 28554 3948
rect 28610 3892 28658 3948
rect 28714 3892 28762 3948
rect 28818 3892 28828 3948
rect 23426 3836 23436 3892
rect 23492 3836 28252 3892
rect 28308 3836 28318 3892
rect 28924 3780 28980 4396
rect 29810 4284 29820 4340
rect 29876 4284 31612 4340
rect 31668 4284 31678 4340
rect 33200 4116 34000 4144
rect 32274 4060 32284 4116
rect 32340 4060 34000 4116
rect 33200 4032 34000 4060
rect 2370 3724 2380 3780
rect 2436 3724 5068 3780
rect 5124 3724 15148 3780
rect 18610 3724 18620 3780
rect 18676 3724 28588 3780
rect 28644 3724 28654 3780
rect 28802 3724 28812 3780
rect 28868 3724 28980 3780
rect 4582 3612 4620 3668
rect 4676 3612 4686 3668
rect 17714 3612 17724 3668
rect 17780 3612 18396 3668
rect 18452 3612 18462 3668
rect 24994 3612 25004 3668
rect 25060 3612 26012 3668
rect 26068 3612 26078 3668
rect 29026 3612 29036 3668
rect 29092 3612 31948 3668
rect 1372 3500 4508 3556
rect 4564 3500 4574 3556
rect 6066 3500 6076 3556
rect 6132 3500 12124 3556
rect 12180 3500 13356 3556
rect 13412 3500 13422 3556
rect 16818 3500 16828 3556
rect 16884 3500 19852 3556
rect 19908 3500 19918 3556
rect 22194 3500 22204 3556
rect 22260 3500 24220 3556
rect 24276 3500 25116 3556
rect 25172 3500 25182 3556
rect 0 3444 800 3472
rect 1372 3444 1428 3500
rect 31892 3444 31948 3612
rect 33200 3444 34000 3472
rect 0 3388 1428 3444
rect 1586 3388 1596 3444
rect 1652 3388 2604 3444
rect 2660 3388 2670 3444
rect 8642 3388 8652 3444
rect 8708 3388 13132 3444
rect 13188 3388 13198 3444
rect 14242 3388 14252 3444
rect 14308 3388 15820 3444
rect 15876 3388 15886 3444
rect 22418 3388 22428 3444
rect 22484 3388 25228 3444
rect 25284 3388 25294 3444
rect 25442 3388 25452 3444
rect 25508 3388 26908 3444
rect 26964 3388 26974 3444
rect 31892 3388 34000 3444
rect 0 3360 800 3388
rect 33200 3360 34000 3388
rect 4162 3276 4172 3332
rect 4228 3276 12348 3332
rect 12404 3276 12414 3332
rect 22866 3276 22876 3332
rect 22932 3276 24556 3332
rect 24612 3276 24622 3332
rect 9014 3108 9024 3164
rect 9080 3108 9128 3164
rect 9184 3108 9232 3164
rect 9288 3108 9298 3164
rect 16826 3108 16836 3164
rect 16892 3108 16940 3164
rect 16996 3108 17044 3164
rect 17100 3108 17110 3164
rect 24638 3108 24648 3164
rect 24704 3108 24752 3164
rect 24808 3108 24856 3164
rect 24912 3108 24922 3164
rect 32450 3108 32460 3164
rect 32516 3108 32564 3164
rect 32620 3108 32668 3164
rect 32724 3108 32734 3164
rect 0 2772 800 2800
rect 33200 2772 34000 2800
rect 0 2716 12236 2772
rect 12292 2716 12302 2772
rect 32162 2716 32172 2772
rect 32228 2716 34000 2772
rect 0 2688 800 2716
rect 33200 2688 34000 2716
rect 0 2100 800 2128
rect 33200 2100 34000 2128
rect 0 2044 3500 2100
rect 3556 2044 3566 2100
rect 28802 2044 28812 2100
rect 28868 2044 34000 2100
rect 0 2016 800 2044
rect 33200 2016 34000 2044
rect 33200 1428 34000 1456
rect 30146 1372 30156 1428
rect 30212 1372 34000 1428
rect 33200 1344 34000 1372
rect 33200 756 34000 784
rect 32050 700 32060 756
rect 32116 700 34000 756
rect 33200 672 34000 700
rect 33200 0 34000 112
<< via3 >>
rect 5118 30548 5174 30604
rect 5222 30548 5278 30604
rect 5326 30548 5382 30604
rect 12930 30548 12986 30604
rect 13034 30548 13090 30604
rect 13138 30548 13194 30604
rect 20742 30548 20798 30604
rect 20846 30548 20902 30604
rect 20950 30548 21006 30604
rect 28554 30548 28610 30604
rect 28658 30548 28714 30604
rect 28762 30548 28818 30604
rect 9024 29764 9080 29820
rect 9128 29764 9184 29820
rect 9232 29764 9288 29820
rect 16836 29764 16892 29820
rect 16940 29764 16996 29820
rect 17044 29764 17100 29820
rect 24648 29764 24704 29820
rect 24752 29764 24808 29820
rect 24856 29764 24912 29820
rect 32460 29764 32516 29820
rect 32564 29764 32620 29820
rect 32668 29764 32724 29820
rect 4956 29036 5012 29092
rect 5118 28980 5174 29036
rect 5222 28980 5278 29036
rect 5326 28980 5382 29036
rect 12930 28980 12986 29036
rect 13034 28980 13090 29036
rect 13138 28980 13194 29036
rect 20742 28980 20798 29036
rect 20846 28980 20902 29036
rect 20950 28980 21006 29036
rect 28554 28980 28610 29036
rect 28658 28980 28714 29036
rect 28762 28980 28818 29036
rect 4844 28588 4900 28644
rect 9024 28196 9080 28252
rect 9128 28196 9184 28252
rect 9232 28196 9288 28252
rect 16836 28196 16892 28252
rect 16940 28196 16996 28252
rect 17044 28196 17100 28252
rect 24648 28196 24704 28252
rect 24752 28196 24808 28252
rect 24856 28196 24912 28252
rect 32460 28196 32516 28252
rect 32564 28196 32620 28252
rect 32668 28196 32724 28252
rect 3388 27468 3444 27524
rect 5118 27412 5174 27468
rect 5222 27412 5278 27468
rect 5326 27412 5382 27468
rect 12930 27412 12986 27468
rect 13034 27412 13090 27468
rect 13138 27412 13194 27468
rect 20742 27412 20798 27468
rect 20846 27412 20902 27468
rect 20950 27412 21006 27468
rect 28554 27412 28610 27468
rect 28658 27412 28714 27468
rect 28762 27412 28818 27468
rect 4620 26908 4676 26964
rect 9024 26628 9080 26684
rect 9128 26628 9184 26684
rect 9232 26628 9288 26684
rect 16836 26628 16892 26684
rect 16940 26628 16996 26684
rect 17044 26628 17100 26684
rect 24648 26628 24704 26684
rect 24752 26628 24808 26684
rect 24856 26628 24912 26684
rect 32460 26628 32516 26684
rect 32564 26628 32620 26684
rect 32668 26628 32724 26684
rect 4172 26012 4228 26068
rect 5118 25844 5174 25900
rect 5222 25844 5278 25900
rect 5326 25844 5382 25900
rect 12930 25844 12986 25900
rect 13034 25844 13090 25900
rect 13138 25844 13194 25900
rect 20742 25844 20798 25900
rect 20846 25844 20902 25900
rect 20950 25844 21006 25900
rect 28554 25844 28610 25900
rect 28658 25844 28714 25900
rect 28762 25844 28818 25900
rect 4732 25228 4788 25284
rect 9024 25060 9080 25116
rect 9128 25060 9184 25116
rect 9232 25060 9288 25116
rect 16836 25060 16892 25116
rect 16940 25060 16996 25116
rect 17044 25060 17100 25116
rect 24648 25060 24704 25116
rect 24752 25060 24808 25116
rect 24856 25060 24912 25116
rect 32460 25060 32516 25116
rect 32564 25060 32620 25116
rect 32668 25060 32724 25116
rect 1932 24556 1988 24612
rect 5118 24276 5174 24332
rect 5222 24276 5278 24332
rect 5326 24276 5382 24332
rect 12930 24276 12986 24332
rect 13034 24276 13090 24332
rect 13138 24276 13194 24332
rect 20742 24276 20798 24332
rect 20846 24276 20902 24332
rect 20950 24276 21006 24332
rect 28554 24276 28610 24332
rect 28658 24276 28714 24332
rect 28762 24276 28818 24332
rect 9024 23492 9080 23548
rect 9128 23492 9184 23548
rect 9232 23492 9288 23548
rect 16836 23492 16892 23548
rect 16940 23492 16996 23548
rect 17044 23492 17100 23548
rect 24648 23492 24704 23548
rect 24752 23492 24808 23548
rect 24856 23492 24912 23548
rect 32460 23492 32516 23548
rect 32564 23492 32620 23548
rect 32668 23492 32724 23548
rect 5118 22708 5174 22764
rect 5222 22708 5278 22764
rect 5326 22708 5382 22764
rect 12930 22708 12986 22764
rect 13034 22708 13090 22764
rect 13138 22708 13194 22764
rect 20742 22708 20798 22764
rect 20846 22708 20902 22764
rect 20950 22708 21006 22764
rect 28554 22708 28610 22764
rect 28658 22708 28714 22764
rect 28762 22708 28818 22764
rect 9024 21924 9080 21980
rect 9128 21924 9184 21980
rect 9232 21924 9288 21980
rect 16836 21924 16892 21980
rect 16940 21924 16996 21980
rect 17044 21924 17100 21980
rect 24648 21924 24704 21980
rect 24752 21924 24808 21980
rect 24856 21924 24912 21980
rect 32460 21924 32516 21980
rect 32564 21924 32620 21980
rect 32668 21924 32724 21980
rect 5118 21140 5174 21196
rect 5222 21140 5278 21196
rect 5326 21140 5382 21196
rect 12930 21140 12986 21196
rect 13034 21140 13090 21196
rect 13138 21140 13194 21196
rect 20742 21140 20798 21196
rect 20846 21140 20902 21196
rect 20950 21140 21006 21196
rect 28554 21140 28610 21196
rect 28658 21140 28714 21196
rect 28762 21140 28818 21196
rect 9024 20356 9080 20412
rect 9128 20356 9184 20412
rect 9232 20356 9288 20412
rect 16836 20356 16892 20412
rect 16940 20356 16996 20412
rect 17044 20356 17100 20412
rect 24648 20356 24704 20412
rect 24752 20356 24808 20412
rect 24856 20356 24912 20412
rect 32460 20356 32516 20412
rect 32564 20356 32620 20412
rect 32668 20356 32724 20412
rect 5118 19572 5174 19628
rect 5222 19572 5278 19628
rect 5326 19572 5382 19628
rect 12930 19572 12986 19628
rect 13034 19572 13090 19628
rect 13138 19572 13194 19628
rect 20742 19572 20798 19628
rect 20846 19572 20902 19628
rect 20950 19572 21006 19628
rect 28554 19572 28610 19628
rect 28658 19572 28714 19628
rect 28762 19572 28818 19628
rect 9024 18788 9080 18844
rect 9128 18788 9184 18844
rect 9232 18788 9288 18844
rect 16836 18788 16892 18844
rect 16940 18788 16996 18844
rect 17044 18788 17100 18844
rect 24648 18788 24704 18844
rect 24752 18788 24808 18844
rect 24856 18788 24912 18844
rect 32460 18788 32516 18844
rect 32564 18788 32620 18844
rect 32668 18788 32724 18844
rect 3500 18396 3556 18452
rect 3500 18172 3556 18228
rect 5118 18004 5174 18060
rect 5222 18004 5278 18060
rect 5326 18004 5382 18060
rect 12930 18004 12986 18060
rect 13034 18004 13090 18060
rect 13138 18004 13194 18060
rect 20742 18004 20798 18060
rect 20846 18004 20902 18060
rect 20950 18004 21006 18060
rect 28554 18004 28610 18060
rect 28658 18004 28714 18060
rect 28762 18004 28818 18060
rect 4844 17836 4900 17892
rect 9024 17220 9080 17276
rect 9128 17220 9184 17276
rect 9232 17220 9288 17276
rect 16836 17220 16892 17276
rect 16940 17220 16996 17276
rect 17044 17220 17100 17276
rect 24648 17220 24704 17276
rect 24752 17220 24808 17276
rect 24856 17220 24912 17276
rect 32460 17220 32516 17276
rect 32564 17220 32620 17276
rect 32668 17220 32724 17276
rect 5118 16436 5174 16492
rect 5222 16436 5278 16492
rect 5326 16436 5382 16492
rect 12930 16436 12986 16492
rect 13034 16436 13090 16492
rect 13138 16436 13194 16492
rect 20742 16436 20798 16492
rect 20846 16436 20902 16492
rect 20950 16436 21006 16492
rect 28554 16436 28610 16492
rect 28658 16436 28714 16492
rect 28762 16436 28818 16492
rect 9024 15652 9080 15708
rect 9128 15652 9184 15708
rect 9232 15652 9288 15708
rect 16836 15652 16892 15708
rect 16940 15652 16996 15708
rect 17044 15652 17100 15708
rect 24648 15652 24704 15708
rect 24752 15652 24808 15708
rect 24856 15652 24912 15708
rect 32460 15652 32516 15708
rect 32564 15652 32620 15708
rect 32668 15652 32724 15708
rect 4732 15036 4788 15092
rect 5118 14868 5174 14924
rect 5222 14868 5278 14924
rect 5326 14868 5382 14924
rect 12930 14868 12986 14924
rect 13034 14868 13090 14924
rect 13138 14868 13194 14924
rect 20742 14868 20798 14924
rect 20846 14868 20902 14924
rect 20950 14868 21006 14924
rect 28554 14868 28610 14924
rect 28658 14868 28714 14924
rect 28762 14868 28818 14924
rect 9024 14084 9080 14140
rect 9128 14084 9184 14140
rect 9232 14084 9288 14140
rect 16836 14084 16892 14140
rect 16940 14084 16996 14140
rect 17044 14084 17100 14140
rect 24648 14084 24704 14140
rect 24752 14084 24808 14140
rect 24856 14084 24912 14140
rect 32460 14084 32516 14140
rect 32564 14084 32620 14140
rect 32668 14084 32724 14140
rect 5118 13300 5174 13356
rect 5222 13300 5278 13356
rect 5326 13300 5382 13356
rect 12930 13300 12986 13356
rect 13034 13300 13090 13356
rect 13138 13300 13194 13356
rect 20742 13300 20798 13356
rect 20846 13300 20902 13356
rect 20950 13300 21006 13356
rect 28554 13300 28610 13356
rect 28658 13300 28714 13356
rect 28762 13300 28818 13356
rect 9024 12516 9080 12572
rect 9128 12516 9184 12572
rect 9232 12516 9288 12572
rect 16836 12516 16892 12572
rect 16940 12516 16996 12572
rect 17044 12516 17100 12572
rect 24648 12516 24704 12572
rect 24752 12516 24808 12572
rect 24856 12516 24912 12572
rect 32460 12516 32516 12572
rect 32564 12516 32620 12572
rect 32668 12516 32724 12572
rect 4172 12012 4228 12068
rect 5118 11732 5174 11788
rect 5222 11732 5278 11788
rect 5326 11732 5382 11788
rect 12930 11732 12986 11788
rect 13034 11732 13090 11788
rect 13138 11732 13194 11788
rect 20742 11732 20798 11788
rect 20846 11732 20902 11788
rect 20950 11732 21006 11788
rect 28554 11732 28610 11788
rect 28658 11732 28714 11788
rect 28762 11732 28818 11788
rect 4172 11340 4228 11396
rect 9024 10948 9080 11004
rect 9128 10948 9184 11004
rect 9232 10948 9288 11004
rect 16836 10948 16892 11004
rect 16940 10948 16996 11004
rect 17044 10948 17100 11004
rect 24648 10948 24704 11004
rect 24752 10948 24808 11004
rect 24856 10948 24912 11004
rect 32460 10948 32516 11004
rect 32564 10948 32620 11004
rect 32668 10948 32724 11004
rect 4956 10780 5012 10836
rect 5118 10164 5174 10220
rect 5222 10164 5278 10220
rect 5326 10164 5382 10220
rect 12930 10164 12986 10220
rect 13034 10164 13090 10220
rect 13138 10164 13194 10220
rect 20742 10164 20798 10220
rect 20846 10164 20902 10220
rect 20950 10164 21006 10220
rect 28554 10164 28610 10220
rect 28658 10164 28714 10220
rect 28762 10164 28818 10220
rect 9024 9380 9080 9436
rect 9128 9380 9184 9436
rect 9232 9380 9288 9436
rect 16836 9380 16892 9436
rect 16940 9380 16996 9436
rect 17044 9380 17100 9436
rect 24648 9380 24704 9436
rect 24752 9380 24808 9436
rect 24856 9380 24912 9436
rect 32460 9380 32516 9436
rect 32564 9380 32620 9436
rect 32668 9380 32724 9436
rect 1932 9100 1988 9156
rect 5118 8596 5174 8652
rect 5222 8596 5278 8652
rect 5326 8596 5382 8652
rect 12930 8596 12986 8652
rect 13034 8596 13090 8652
rect 13138 8596 13194 8652
rect 20742 8596 20798 8652
rect 20846 8596 20902 8652
rect 20950 8596 21006 8652
rect 28554 8596 28610 8652
rect 28658 8596 28714 8652
rect 28762 8596 28818 8652
rect 9024 7812 9080 7868
rect 9128 7812 9184 7868
rect 9232 7812 9288 7868
rect 16836 7812 16892 7868
rect 16940 7812 16996 7868
rect 17044 7812 17100 7868
rect 24648 7812 24704 7868
rect 24752 7812 24808 7868
rect 24856 7812 24912 7868
rect 32460 7812 32516 7868
rect 32564 7812 32620 7868
rect 32668 7812 32724 7868
rect 5118 7028 5174 7084
rect 5222 7028 5278 7084
rect 5326 7028 5382 7084
rect 12930 7028 12986 7084
rect 13034 7028 13090 7084
rect 13138 7028 13194 7084
rect 20742 7028 20798 7084
rect 20846 7028 20902 7084
rect 20950 7028 21006 7084
rect 28554 7028 28610 7084
rect 28658 7028 28714 7084
rect 28762 7028 28818 7084
rect 3388 6636 3444 6692
rect 9024 6244 9080 6300
rect 9128 6244 9184 6300
rect 9232 6244 9288 6300
rect 16836 6244 16892 6300
rect 16940 6244 16996 6300
rect 17044 6244 17100 6300
rect 24648 6244 24704 6300
rect 24752 6244 24808 6300
rect 24856 6244 24912 6300
rect 32460 6244 32516 6300
rect 32564 6244 32620 6300
rect 32668 6244 32724 6300
rect 4172 6188 4228 6244
rect 5118 5460 5174 5516
rect 5222 5460 5278 5516
rect 5326 5460 5382 5516
rect 12930 5460 12986 5516
rect 13034 5460 13090 5516
rect 13138 5460 13194 5516
rect 20742 5460 20798 5516
rect 20846 5460 20902 5516
rect 20950 5460 21006 5516
rect 28554 5460 28610 5516
rect 28658 5460 28714 5516
rect 28762 5460 28818 5516
rect 9024 4676 9080 4732
rect 9128 4676 9184 4732
rect 9232 4676 9288 4732
rect 16836 4676 16892 4732
rect 16940 4676 16996 4732
rect 17044 4676 17100 4732
rect 24648 4676 24704 4732
rect 24752 4676 24808 4732
rect 24856 4676 24912 4732
rect 32460 4676 32516 4732
rect 32564 4676 32620 4732
rect 32668 4676 32724 4732
rect 4620 4396 4676 4452
rect 5118 3892 5174 3948
rect 5222 3892 5278 3948
rect 5326 3892 5382 3948
rect 12930 3892 12986 3948
rect 13034 3892 13090 3948
rect 13138 3892 13194 3948
rect 20742 3892 20798 3948
rect 20846 3892 20902 3948
rect 20950 3892 21006 3948
rect 28554 3892 28610 3948
rect 28658 3892 28714 3948
rect 28762 3892 28818 3948
rect 4620 3612 4676 3668
rect 9024 3108 9080 3164
rect 9128 3108 9184 3164
rect 9232 3108 9288 3164
rect 16836 3108 16892 3164
rect 16940 3108 16996 3164
rect 17044 3108 17100 3164
rect 24648 3108 24704 3164
rect 24752 3108 24808 3164
rect 24856 3108 24912 3164
rect 32460 3108 32516 3164
rect 32564 3108 32620 3164
rect 32668 3108 32724 3164
<< metal4 >>
rect 5090 30604 5410 30636
rect 5090 30548 5118 30604
rect 5174 30548 5222 30604
rect 5278 30548 5326 30604
rect 5382 30548 5410 30604
rect 4956 29092 5012 29102
rect 4844 28644 4900 28654
rect 3388 27524 3444 27534
rect 1932 24612 1988 24622
rect 1932 9156 1988 24556
rect 1932 9090 1988 9100
rect 3388 6692 3444 27468
rect 4620 26964 4676 26974
rect 4172 26068 4228 26078
rect 3500 18452 3556 18462
rect 3500 18228 3556 18396
rect 3500 18162 3556 18172
rect 4172 12068 4228 26012
rect 4172 12002 4228 12012
rect 3388 6626 3444 6636
rect 4172 11396 4228 11406
rect 4172 6244 4228 11340
rect 4172 6178 4228 6188
rect 4620 4452 4676 26908
rect 4732 25284 4788 25294
rect 4732 15092 4788 25228
rect 4844 17892 4900 28588
rect 4844 17826 4900 17836
rect 4732 15026 4788 15036
rect 4956 10836 5012 29036
rect 4956 10770 5012 10780
rect 5090 29036 5410 30548
rect 5090 28980 5118 29036
rect 5174 28980 5222 29036
rect 5278 28980 5326 29036
rect 5382 28980 5410 29036
rect 5090 27468 5410 28980
rect 5090 27412 5118 27468
rect 5174 27412 5222 27468
rect 5278 27412 5326 27468
rect 5382 27412 5410 27468
rect 5090 25900 5410 27412
rect 5090 25844 5118 25900
rect 5174 25844 5222 25900
rect 5278 25844 5326 25900
rect 5382 25844 5410 25900
rect 5090 24332 5410 25844
rect 5090 24276 5118 24332
rect 5174 24276 5222 24332
rect 5278 24276 5326 24332
rect 5382 24276 5410 24332
rect 5090 22764 5410 24276
rect 5090 22708 5118 22764
rect 5174 22708 5222 22764
rect 5278 22708 5326 22764
rect 5382 22708 5410 22764
rect 5090 21196 5410 22708
rect 5090 21140 5118 21196
rect 5174 21140 5222 21196
rect 5278 21140 5326 21196
rect 5382 21140 5410 21196
rect 5090 19628 5410 21140
rect 5090 19572 5118 19628
rect 5174 19572 5222 19628
rect 5278 19572 5326 19628
rect 5382 19572 5410 19628
rect 5090 18060 5410 19572
rect 5090 18004 5118 18060
rect 5174 18004 5222 18060
rect 5278 18004 5326 18060
rect 5382 18004 5410 18060
rect 5090 16492 5410 18004
rect 5090 16436 5118 16492
rect 5174 16436 5222 16492
rect 5278 16436 5326 16492
rect 5382 16436 5410 16492
rect 5090 14924 5410 16436
rect 5090 14868 5118 14924
rect 5174 14868 5222 14924
rect 5278 14868 5326 14924
rect 5382 14868 5410 14924
rect 5090 13356 5410 14868
rect 5090 13300 5118 13356
rect 5174 13300 5222 13356
rect 5278 13300 5326 13356
rect 5382 13300 5410 13356
rect 5090 11788 5410 13300
rect 5090 11732 5118 11788
rect 5174 11732 5222 11788
rect 5278 11732 5326 11788
rect 5382 11732 5410 11788
rect 4620 3668 4676 4396
rect 4620 3602 4676 3612
rect 5090 10220 5410 11732
rect 5090 10164 5118 10220
rect 5174 10164 5222 10220
rect 5278 10164 5326 10220
rect 5382 10164 5410 10220
rect 5090 8652 5410 10164
rect 5090 8596 5118 8652
rect 5174 8596 5222 8652
rect 5278 8596 5326 8652
rect 5382 8596 5410 8652
rect 5090 7084 5410 8596
rect 5090 7028 5118 7084
rect 5174 7028 5222 7084
rect 5278 7028 5326 7084
rect 5382 7028 5410 7084
rect 5090 5516 5410 7028
rect 5090 5460 5118 5516
rect 5174 5460 5222 5516
rect 5278 5460 5326 5516
rect 5382 5460 5410 5516
rect 5090 3948 5410 5460
rect 5090 3892 5118 3948
rect 5174 3892 5222 3948
rect 5278 3892 5326 3948
rect 5382 3892 5410 3948
rect 5090 3076 5410 3892
rect 8996 29820 9316 30636
rect 8996 29764 9024 29820
rect 9080 29764 9128 29820
rect 9184 29764 9232 29820
rect 9288 29764 9316 29820
rect 8996 28252 9316 29764
rect 8996 28196 9024 28252
rect 9080 28196 9128 28252
rect 9184 28196 9232 28252
rect 9288 28196 9316 28252
rect 8996 26684 9316 28196
rect 8996 26628 9024 26684
rect 9080 26628 9128 26684
rect 9184 26628 9232 26684
rect 9288 26628 9316 26684
rect 8996 25116 9316 26628
rect 8996 25060 9024 25116
rect 9080 25060 9128 25116
rect 9184 25060 9232 25116
rect 9288 25060 9316 25116
rect 8996 23548 9316 25060
rect 8996 23492 9024 23548
rect 9080 23492 9128 23548
rect 9184 23492 9232 23548
rect 9288 23492 9316 23548
rect 8996 21980 9316 23492
rect 8996 21924 9024 21980
rect 9080 21924 9128 21980
rect 9184 21924 9232 21980
rect 9288 21924 9316 21980
rect 8996 20412 9316 21924
rect 8996 20356 9024 20412
rect 9080 20356 9128 20412
rect 9184 20356 9232 20412
rect 9288 20356 9316 20412
rect 8996 18844 9316 20356
rect 8996 18788 9024 18844
rect 9080 18788 9128 18844
rect 9184 18788 9232 18844
rect 9288 18788 9316 18844
rect 8996 17276 9316 18788
rect 8996 17220 9024 17276
rect 9080 17220 9128 17276
rect 9184 17220 9232 17276
rect 9288 17220 9316 17276
rect 8996 15708 9316 17220
rect 8996 15652 9024 15708
rect 9080 15652 9128 15708
rect 9184 15652 9232 15708
rect 9288 15652 9316 15708
rect 8996 14140 9316 15652
rect 8996 14084 9024 14140
rect 9080 14084 9128 14140
rect 9184 14084 9232 14140
rect 9288 14084 9316 14140
rect 8996 12572 9316 14084
rect 8996 12516 9024 12572
rect 9080 12516 9128 12572
rect 9184 12516 9232 12572
rect 9288 12516 9316 12572
rect 8996 11004 9316 12516
rect 8996 10948 9024 11004
rect 9080 10948 9128 11004
rect 9184 10948 9232 11004
rect 9288 10948 9316 11004
rect 8996 9436 9316 10948
rect 8996 9380 9024 9436
rect 9080 9380 9128 9436
rect 9184 9380 9232 9436
rect 9288 9380 9316 9436
rect 8996 7868 9316 9380
rect 8996 7812 9024 7868
rect 9080 7812 9128 7868
rect 9184 7812 9232 7868
rect 9288 7812 9316 7868
rect 8996 6300 9316 7812
rect 8996 6244 9024 6300
rect 9080 6244 9128 6300
rect 9184 6244 9232 6300
rect 9288 6244 9316 6300
rect 8996 4732 9316 6244
rect 8996 4676 9024 4732
rect 9080 4676 9128 4732
rect 9184 4676 9232 4732
rect 9288 4676 9316 4732
rect 8996 3164 9316 4676
rect 8996 3108 9024 3164
rect 9080 3108 9128 3164
rect 9184 3108 9232 3164
rect 9288 3108 9316 3164
rect 8996 3076 9316 3108
rect 12902 30604 13222 30636
rect 12902 30548 12930 30604
rect 12986 30548 13034 30604
rect 13090 30548 13138 30604
rect 13194 30548 13222 30604
rect 12902 29036 13222 30548
rect 12902 28980 12930 29036
rect 12986 28980 13034 29036
rect 13090 28980 13138 29036
rect 13194 28980 13222 29036
rect 12902 27468 13222 28980
rect 12902 27412 12930 27468
rect 12986 27412 13034 27468
rect 13090 27412 13138 27468
rect 13194 27412 13222 27468
rect 12902 25900 13222 27412
rect 12902 25844 12930 25900
rect 12986 25844 13034 25900
rect 13090 25844 13138 25900
rect 13194 25844 13222 25900
rect 12902 24332 13222 25844
rect 12902 24276 12930 24332
rect 12986 24276 13034 24332
rect 13090 24276 13138 24332
rect 13194 24276 13222 24332
rect 12902 22764 13222 24276
rect 12902 22708 12930 22764
rect 12986 22708 13034 22764
rect 13090 22708 13138 22764
rect 13194 22708 13222 22764
rect 12902 21196 13222 22708
rect 12902 21140 12930 21196
rect 12986 21140 13034 21196
rect 13090 21140 13138 21196
rect 13194 21140 13222 21196
rect 12902 19628 13222 21140
rect 12902 19572 12930 19628
rect 12986 19572 13034 19628
rect 13090 19572 13138 19628
rect 13194 19572 13222 19628
rect 12902 18060 13222 19572
rect 12902 18004 12930 18060
rect 12986 18004 13034 18060
rect 13090 18004 13138 18060
rect 13194 18004 13222 18060
rect 12902 16492 13222 18004
rect 12902 16436 12930 16492
rect 12986 16436 13034 16492
rect 13090 16436 13138 16492
rect 13194 16436 13222 16492
rect 12902 14924 13222 16436
rect 12902 14868 12930 14924
rect 12986 14868 13034 14924
rect 13090 14868 13138 14924
rect 13194 14868 13222 14924
rect 12902 13356 13222 14868
rect 12902 13300 12930 13356
rect 12986 13300 13034 13356
rect 13090 13300 13138 13356
rect 13194 13300 13222 13356
rect 12902 11788 13222 13300
rect 12902 11732 12930 11788
rect 12986 11732 13034 11788
rect 13090 11732 13138 11788
rect 13194 11732 13222 11788
rect 12902 10220 13222 11732
rect 12902 10164 12930 10220
rect 12986 10164 13034 10220
rect 13090 10164 13138 10220
rect 13194 10164 13222 10220
rect 12902 8652 13222 10164
rect 12902 8596 12930 8652
rect 12986 8596 13034 8652
rect 13090 8596 13138 8652
rect 13194 8596 13222 8652
rect 12902 7084 13222 8596
rect 12902 7028 12930 7084
rect 12986 7028 13034 7084
rect 13090 7028 13138 7084
rect 13194 7028 13222 7084
rect 12902 5516 13222 7028
rect 12902 5460 12930 5516
rect 12986 5460 13034 5516
rect 13090 5460 13138 5516
rect 13194 5460 13222 5516
rect 12902 3948 13222 5460
rect 12902 3892 12930 3948
rect 12986 3892 13034 3948
rect 13090 3892 13138 3948
rect 13194 3892 13222 3948
rect 12902 3076 13222 3892
rect 16808 29820 17128 30636
rect 16808 29764 16836 29820
rect 16892 29764 16940 29820
rect 16996 29764 17044 29820
rect 17100 29764 17128 29820
rect 16808 28252 17128 29764
rect 16808 28196 16836 28252
rect 16892 28196 16940 28252
rect 16996 28196 17044 28252
rect 17100 28196 17128 28252
rect 16808 26684 17128 28196
rect 16808 26628 16836 26684
rect 16892 26628 16940 26684
rect 16996 26628 17044 26684
rect 17100 26628 17128 26684
rect 16808 25116 17128 26628
rect 16808 25060 16836 25116
rect 16892 25060 16940 25116
rect 16996 25060 17044 25116
rect 17100 25060 17128 25116
rect 16808 23548 17128 25060
rect 16808 23492 16836 23548
rect 16892 23492 16940 23548
rect 16996 23492 17044 23548
rect 17100 23492 17128 23548
rect 16808 21980 17128 23492
rect 16808 21924 16836 21980
rect 16892 21924 16940 21980
rect 16996 21924 17044 21980
rect 17100 21924 17128 21980
rect 16808 20412 17128 21924
rect 16808 20356 16836 20412
rect 16892 20356 16940 20412
rect 16996 20356 17044 20412
rect 17100 20356 17128 20412
rect 16808 18844 17128 20356
rect 16808 18788 16836 18844
rect 16892 18788 16940 18844
rect 16996 18788 17044 18844
rect 17100 18788 17128 18844
rect 16808 17276 17128 18788
rect 16808 17220 16836 17276
rect 16892 17220 16940 17276
rect 16996 17220 17044 17276
rect 17100 17220 17128 17276
rect 16808 15708 17128 17220
rect 16808 15652 16836 15708
rect 16892 15652 16940 15708
rect 16996 15652 17044 15708
rect 17100 15652 17128 15708
rect 16808 14140 17128 15652
rect 16808 14084 16836 14140
rect 16892 14084 16940 14140
rect 16996 14084 17044 14140
rect 17100 14084 17128 14140
rect 16808 12572 17128 14084
rect 16808 12516 16836 12572
rect 16892 12516 16940 12572
rect 16996 12516 17044 12572
rect 17100 12516 17128 12572
rect 16808 11004 17128 12516
rect 16808 10948 16836 11004
rect 16892 10948 16940 11004
rect 16996 10948 17044 11004
rect 17100 10948 17128 11004
rect 16808 9436 17128 10948
rect 16808 9380 16836 9436
rect 16892 9380 16940 9436
rect 16996 9380 17044 9436
rect 17100 9380 17128 9436
rect 16808 7868 17128 9380
rect 16808 7812 16836 7868
rect 16892 7812 16940 7868
rect 16996 7812 17044 7868
rect 17100 7812 17128 7868
rect 16808 6300 17128 7812
rect 16808 6244 16836 6300
rect 16892 6244 16940 6300
rect 16996 6244 17044 6300
rect 17100 6244 17128 6300
rect 16808 4732 17128 6244
rect 16808 4676 16836 4732
rect 16892 4676 16940 4732
rect 16996 4676 17044 4732
rect 17100 4676 17128 4732
rect 16808 3164 17128 4676
rect 16808 3108 16836 3164
rect 16892 3108 16940 3164
rect 16996 3108 17044 3164
rect 17100 3108 17128 3164
rect 16808 3076 17128 3108
rect 20714 30604 21034 30636
rect 20714 30548 20742 30604
rect 20798 30548 20846 30604
rect 20902 30548 20950 30604
rect 21006 30548 21034 30604
rect 20714 29036 21034 30548
rect 20714 28980 20742 29036
rect 20798 28980 20846 29036
rect 20902 28980 20950 29036
rect 21006 28980 21034 29036
rect 20714 27468 21034 28980
rect 20714 27412 20742 27468
rect 20798 27412 20846 27468
rect 20902 27412 20950 27468
rect 21006 27412 21034 27468
rect 20714 25900 21034 27412
rect 20714 25844 20742 25900
rect 20798 25844 20846 25900
rect 20902 25844 20950 25900
rect 21006 25844 21034 25900
rect 20714 24332 21034 25844
rect 20714 24276 20742 24332
rect 20798 24276 20846 24332
rect 20902 24276 20950 24332
rect 21006 24276 21034 24332
rect 20714 22764 21034 24276
rect 20714 22708 20742 22764
rect 20798 22708 20846 22764
rect 20902 22708 20950 22764
rect 21006 22708 21034 22764
rect 20714 21196 21034 22708
rect 20714 21140 20742 21196
rect 20798 21140 20846 21196
rect 20902 21140 20950 21196
rect 21006 21140 21034 21196
rect 20714 19628 21034 21140
rect 20714 19572 20742 19628
rect 20798 19572 20846 19628
rect 20902 19572 20950 19628
rect 21006 19572 21034 19628
rect 20714 18060 21034 19572
rect 20714 18004 20742 18060
rect 20798 18004 20846 18060
rect 20902 18004 20950 18060
rect 21006 18004 21034 18060
rect 20714 16492 21034 18004
rect 20714 16436 20742 16492
rect 20798 16436 20846 16492
rect 20902 16436 20950 16492
rect 21006 16436 21034 16492
rect 20714 14924 21034 16436
rect 20714 14868 20742 14924
rect 20798 14868 20846 14924
rect 20902 14868 20950 14924
rect 21006 14868 21034 14924
rect 20714 13356 21034 14868
rect 20714 13300 20742 13356
rect 20798 13300 20846 13356
rect 20902 13300 20950 13356
rect 21006 13300 21034 13356
rect 20714 11788 21034 13300
rect 20714 11732 20742 11788
rect 20798 11732 20846 11788
rect 20902 11732 20950 11788
rect 21006 11732 21034 11788
rect 20714 10220 21034 11732
rect 20714 10164 20742 10220
rect 20798 10164 20846 10220
rect 20902 10164 20950 10220
rect 21006 10164 21034 10220
rect 20714 8652 21034 10164
rect 20714 8596 20742 8652
rect 20798 8596 20846 8652
rect 20902 8596 20950 8652
rect 21006 8596 21034 8652
rect 20714 7084 21034 8596
rect 20714 7028 20742 7084
rect 20798 7028 20846 7084
rect 20902 7028 20950 7084
rect 21006 7028 21034 7084
rect 20714 5516 21034 7028
rect 20714 5460 20742 5516
rect 20798 5460 20846 5516
rect 20902 5460 20950 5516
rect 21006 5460 21034 5516
rect 20714 3948 21034 5460
rect 20714 3892 20742 3948
rect 20798 3892 20846 3948
rect 20902 3892 20950 3948
rect 21006 3892 21034 3948
rect 20714 3076 21034 3892
rect 24620 29820 24940 30636
rect 24620 29764 24648 29820
rect 24704 29764 24752 29820
rect 24808 29764 24856 29820
rect 24912 29764 24940 29820
rect 24620 28252 24940 29764
rect 24620 28196 24648 28252
rect 24704 28196 24752 28252
rect 24808 28196 24856 28252
rect 24912 28196 24940 28252
rect 24620 26684 24940 28196
rect 24620 26628 24648 26684
rect 24704 26628 24752 26684
rect 24808 26628 24856 26684
rect 24912 26628 24940 26684
rect 24620 25116 24940 26628
rect 24620 25060 24648 25116
rect 24704 25060 24752 25116
rect 24808 25060 24856 25116
rect 24912 25060 24940 25116
rect 24620 23548 24940 25060
rect 24620 23492 24648 23548
rect 24704 23492 24752 23548
rect 24808 23492 24856 23548
rect 24912 23492 24940 23548
rect 24620 21980 24940 23492
rect 24620 21924 24648 21980
rect 24704 21924 24752 21980
rect 24808 21924 24856 21980
rect 24912 21924 24940 21980
rect 24620 20412 24940 21924
rect 24620 20356 24648 20412
rect 24704 20356 24752 20412
rect 24808 20356 24856 20412
rect 24912 20356 24940 20412
rect 24620 18844 24940 20356
rect 24620 18788 24648 18844
rect 24704 18788 24752 18844
rect 24808 18788 24856 18844
rect 24912 18788 24940 18844
rect 24620 17276 24940 18788
rect 24620 17220 24648 17276
rect 24704 17220 24752 17276
rect 24808 17220 24856 17276
rect 24912 17220 24940 17276
rect 24620 15708 24940 17220
rect 24620 15652 24648 15708
rect 24704 15652 24752 15708
rect 24808 15652 24856 15708
rect 24912 15652 24940 15708
rect 24620 14140 24940 15652
rect 24620 14084 24648 14140
rect 24704 14084 24752 14140
rect 24808 14084 24856 14140
rect 24912 14084 24940 14140
rect 24620 12572 24940 14084
rect 24620 12516 24648 12572
rect 24704 12516 24752 12572
rect 24808 12516 24856 12572
rect 24912 12516 24940 12572
rect 24620 11004 24940 12516
rect 24620 10948 24648 11004
rect 24704 10948 24752 11004
rect 24808 10948 24856 11004
rect 24912 10948 24940 11004
rect 24620 9436 24940 10948
rect 24620 9380 24648 9436
rect 24704 9380 24752 9436
rect 24808 9380 24856 9436
rect 24912 9380 24940 9436
rect 24620 7868 24940 9380
rect 24620 7812 24648 7868
rect 24704 7812 24752 7868
rect 24808 7812 24856 7868
rect 24912 7812 24940 7868
rect 24620 6300 24940 7812
rect 24620 6244 24648 6300
rect 24704 6244 24752 6300
rect 24808 6244 24856 6300
rect 24912 6244 24940 6300
rect 24620 4732 24940 6244
rect 24620 4676 24648 4732
rect 24704 4676 24752 4732
rect 24808 4676 24856 4732
rect 24912 4676 24940 4732
rect 24620 3164 24940 4676
rect 24620 3108 24648 3164
rect 24704 3108 24752 3164
rect 24808 3108 24856 3164
rect 24912 3108 24940 3164
rect 24620 3076 24940 3108
rect 28526 30604 28846 30636
rect 28526 30548 28554 30604
rect 28610 30548 28658 30604
rect 28714 30548 28762 30604
rect 28818 30548 28846 30604
rect 28526 29036 28846 30548
rect 28526 28980 28554 29036
rect 28610 28980 28658 29036
rect 28714 28980 28762 29036
rect 28818 28980 28846 29036
rect 28526 27468 28846 28980
rect 28526 27412 28554 27468
rect 28610 27412 28658 27468
rect 28714 27412 28762 27468
rect 28818 27412 28846 27468
rect 28526 25900 28846 27412
rect 28526 25844 28554 25900
rect 28610 25844 28658 25900
rect 28714 25844 28762 25900
rect 28818 25844 28846 25900
rect 28526 24332 28846 25844
rect 28526 24276 28554 24332
rect 28610 24276 28658 24332
rect 28714 24276 28762 24332
rect 28818 24276 28846 24332
rect 28526 22764 28846 24276
rect 28526 22708 28554 22764
rect 28610 22708 28658 22764
rect 28714 22708 28762 22764
rect 28818 22708 28846 22764
rect 28526 21196 28846 22708
rect 28526 21140 28554 21196
rect 28610 21140 28658 21196
rect 28714 21140 28762 21196
rect 28818 21140 28846 21196
rect 28526 19628 28846 21140
rect 28526 19572 28554 19628
rect 28610 19572 28658 19628
rect 28714 19572 28762 19628
rect 28818 19572 28846 19628
rect 28526 18060 28846 19572
rect 28526 18004 28554 18060
rect 28610 18004 28658 18060
rect 28714 18004 28762 18060
rect 28818 18004 28846 18060
rect 28526 16492 28846 18004
rect 28526 16436 28554 16492
rect 28610 16436 28658 16492
rect 28714 16436 28762 16492
rect 28818 16436 28846 16492
rect 28526 14924 28846 16436
rect 28526 14868 28554 14924
rect 28610 14868 28658 14924
rect 28714 14868 28762 14924
rect 28818 14868 28846 14924
rect 28526 13356 28846 14868
rect 28526 13300 28554 13356
rect 28610 13300 28658 13356
rect 28714 13300 28762 13356
rect 28818 13300 28846 13356
rect 28526 11788 28846 13300
rect 28526 11732 28554 11788
rect 28610 11732 28658 11788
rect 28714 11732 28762 11788
rect 28818 11732 28846 11788
rect 28526 10220 28846 11732
rect 28526 10164 28554 10220
rect 28610 10164 28658 10220
rect 28714 10164 28762 10220
rect 28818 10164 28846 10220
rect 28526 8652 28846 10164
rect 28526 8596 28554 8652
rect 28610 8596 28658 8652
rect 28714 8596 28762 8652
rect 28818 8596 28846 8652
rect 28526 7084 28846 8596
rect 28526 7028 28554 7084
rect 28610 7028 28658 7084
rect 28714 7028 28762 7084
rect 28818 7028 28846 7084
rect 28526 5516 28846 7028
rect 28526 5460 28554 5516
rect 28610 5460 28658 5516
rect 28714 5460 28762 5516
rect 28818 5460 28846 5516
rect 28526 3948 28846 5460
rect 28526 3892 28554 3948
rect 28610 3892 28658 3948
rect 28714 3892 28762 3948
rect 28818 3892 28846 3948
rect 28526 3076 28846 3892
rect 32432 29820 32752 30636
rect 32432 29764 32460 29820
rect 32516 29764 32564 29820
rect 32620 29764 32668 29820
rect 32724 29764 32752 29820
rect 32432 28252 32752 29764
rect 32432 28196 32460 28252
rect 32516 28196 32564 28252
rect 32620 28196 32668 28252
rect 32724 28196 32752 28252
rect 32432 26684 32752 28196
rect 32432 26628 32460 26684
rect 32516 26628 32564 26684
rect 32620 26628 32668 26684
rect 32724 26628 32752 26684
rect 32432 25116 32752 26628
rect 32432 25060 32460 25116
rect 32516 25060 32564 25116
rect 32620 25060 32668 25116
rect 32724 25060 32752 25116
rect 32432 23548 32752 25060
rect 32432 23492 32460 23548
rect 32516 23492 32564 23548
rect 32620 23492 32668 23548
rect 32724 23492 32752 23548
rect 32432 21980 32752 23492
rect 32432 21924 32460 21980
rect 32516 21924 32564 21980
rect 32620 21924 32668 21980
rect 32724 21924 32752 21980
rect 32432 20412 32752 21924
rect 32432 20356 32460 20412
rect 32516 20356 32564 20412
rect 32620 20356 32668 20412
rect 32724 20356 32752 20412
rect 32432 18844 32752 20356
rect 32432 18788 32460 18844
rect 32516 18788 32564 18844
rect 32620 18788 32668 18844
rect 32724 18788 32752 18844
rect 32432 17276 32752 18788
rect 32432 17220 32460 17276
rect 32516 17220 32564 17276
rect 32620 17220 32668 17276
rect 32724 17220 32752 17276
rect 32432 15708 32752 17220
rect 32432 15652 32460 15708
rect 32516 15652 32564 15708
rect 32620 15652 32668 15708
rect 32724 15652 32752 15708
rect 32432 14140 32752 15652
rect 32432 14084 32460 14140
rect 32516 14084 32564 14140
rect 32620 14084 32668 14140
rect 32724 14084 32752 14140
rect 32432 12572 32752 14084
rect 32432 12516 32460 12572
rect 32516 12516 32564 12572
rect 32620 12516 32668 12572
rect 32724 12516 32752 12572
rect 32432 11004 32752 12516
rect 32432 10948 32460 11004
rect 32516 10948 32564 11004
rect 32620 10948 32668 11004
rect 32724 10948 32752 11004
rect 32432 9436 32752 10948
rect 32432 9380 32460 9436
rect 32516 9380 32564 9436
rect 32620 9380 32668 9436
rect 32724 9380 32752 9436
rect 32432 7868 32752 9380
rect 32432 7812 32460 7868
rect 32516 7812 32564 7868
rect 32620 7812 32668 7868
rect 32724 7812 32752 7868
rect 32432 6300 32752 7812
rect 32432 6244 32460 6300
rect 32516 6244 32564 6300
rect 32620 6244 32668 6300
rect 32724 6244 32752 6300
rect 32432 4732 32752 6244
rect 32432 4676 32460 4732
rect 32516 4676 32564 4732
rect 32620 4676 32668 4732
rect 32724 4676 32752 4732
rect 32432 3164 32752 4676
rect 32432 3108 32460 3164
rect 32516 3108 32564 3164
rect 32620 3108 32668 3164
rect 32724 3108 32752 3164
rect 32432 3076 32752 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14560 0 1 20384
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _120_
timestamp 1698431365
transform 1 0 10752 0 -1 10976
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _122_
timestamp 1698431365
transform -1 0 14448 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _123_
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _124_
timestamp 1698431365
transform -1 0 6608 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _125_
timestamp 1698431365
transform 1 0 20048 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _126_
timestamp 1698431365
transform 1 0 21168 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _127_
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _128_
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _129_
timestamp 1698431365
transform -1 0 16688 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _130_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _131_
timestamp 1698431365
transform 1 0 8400 0 1 10976
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _132_
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _133_
timestamp 1698431365
transform 1 0 7056 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _134_
timestamp 1698431365
transform 1 0 5600 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _135_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _136_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _137_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _138_
timestamp 1698431365
transform -1 0 6944 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _139_
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _140_
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _141_
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _142_
timestamp 1698431365
transform -1 0 13664 0 -1 12544
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _143_
timestamp 1698431365
transform 1 0 21728 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _144_
timestamp 1698431365
transform -1 0 20048 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _145_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _146_
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _147_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _148_
timestamp 1698431365
transform -1 0 15568 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _149_
timestamp 1698431365
transform -1 0 14448 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _150_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _151_
timestamp 1698431365
transform -1 0 20720 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _152_
timestamp 1698431365
transform -1 0 18368 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _153_
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _154_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _155_
timestamp 1698431365
transform -1 0 28000 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _156_
timestamp 1698431365
transform 1 0 27216 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _157_
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _158_
timestamp 1698431365
transform -1 0 31248 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _159_
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _160_
timestamp 1698431365
transform 1 0 31248 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _161_
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _162_
timestamp 1698431365
transform -1 0 26208 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _163_
timestamp 1698431365
transform -1 0 23408 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _166_
timestamp 1698431365
transform -1 0 25760 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _167_
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _168_
timestamp 1698431365
transform -1 0 22512 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _169_
timestamp 1698431365
transform -1 0 20608 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _170_
timestamp 1698431365
transform -1 0 18368 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _171_
timestamp 1698431365
transform -1 0 24864 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _172_
timestamp 1698431365
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _173_
timestamp 1698431365
transform -1 0 20048 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _174_
timestamp 1698431365
transform -1 0 19936 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _175_
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _176_
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _177_
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _178_
timestamp 1698431365
transform -1 0 32032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _179_
timestamp 1698431365
transform -1 0 32368 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _180_
timestamp 1698431365
transform -1 0 32368 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _181_
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _182_
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _183_
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _184_
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _185_
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _186_
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _187_
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _188_
timestamp 1698431365
transform -1 0 26880 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _189_
timestamp 1698431365
transform 1 0 21728 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _190_
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _191_
timestamp 1698431365
transform 1 0 27888 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _192_
timestamp 1698431365
transform 1 0 27888 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _193_
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _194_
timestamp 1698431365
transform -1 0 18592 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _195_
timestamp 1698431365
transform -1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _196_
timestamp 1698431365
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _197_
timestamp 1698431365
transform -1 0 15120 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _198_
timestamp 1698431365
transform -1 0 11200 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _199_
timestamp 1698431365
transform -1 0 6384 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _200_
timestamp 1698431365
transform 1 0 1792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _201_
timestamp 1698431365
transform 1 0 1792 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _202_
timestamp 1698431365
transform -1 0 11424 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _203_
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _204_
timestamp 1698431365
transform -1 0 12656 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _205_
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _206_
timestamp 1698431365
transform -1 0 16464 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _207_
timestamp 1698431365
transform -1 0 15792 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _208_
timestamp 1698431365
transform -1 0 24752 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _209_
timestamp 1698431365
transform 1 0 27216 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _210_
timestamp 1698431365
transform 1 0 21280 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _211_
timestamp 1698431365
transform -1 0 27216 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _212_
timestamp 1698431365
transform -1 0 21840 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _213_
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _214_
timestamp 1698431365
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _215_
timestamp 1698431365
transform -1 0 24080 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _216_
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _217_
timestamp 1698431365
transform -1 0 20496 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _218_
timestamp 1698431365
transform -1 0 18592 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _219_
timestamp 1698431365
transform 1 0 13440 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _220_
timestamp 1698431365
transform -1 0 14224 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _221_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _222_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _223_
timestamp 1698431365
transform -1 0 12992 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _224_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _225_
timestamp 1698431365
transform -1 0 10080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _226_
timestamp 1698431365
transform 1 0 3472 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _227_
timestamp 1698431365
transform -1 0 2464 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _228_
timestamp 1698431365
transform -1 0 7952 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _229_
timestamp 1698431365
transform -1 0 6496 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _230_
timestamp 1698431365
transform -1 0 10080 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _231_
timestamp 1698431365
transform -1 0 8848 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _232_
timestamp 1698431365
transform -1 0 14000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _233_
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _234_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _235_
timestamp 1698431365
transform 1 0 14896 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _236_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _237_
timestamp 1698431365
transform 1 0 12544 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _238_
timestamp 1698431365
transform 1 0 10416 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _239_
timestamp 1698431365
transform -1 0 11984 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _240_
timestamp 1698431365
transform 1 0 6272 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _241_
timestamp 1698431365
transform -1 0 7840 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _242_
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _243_
timestamp 1698431365
transform -1 0 5376 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _244_
timestamp 1698431365
transform 1 0 13104 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _245_
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _246_
timestamp 1698431365
transform -1 0 11984 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _247_
timestamp 1698431365
transform -1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _248_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _249_
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _250_
timestamp 1698431365
transform -1 0 5376 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _251_
timestamp 1698431365
transform -1 0 5376 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _252_
timestamp 1698431365
transform 1 0 5376 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _253_
timestamp 1698431365
transform 1 0 4368 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _254_
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _255_
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _256_
timestamp 1698431365
transform -1 0 23856 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _257_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _258_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _259_
timestamp 1698431365
transform 1 0 18256 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _260_
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _261_
timestamp 1698431365
transform 1 0 13216 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _262_
timestamp 1698431365
transform 1 0 11088 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _263_
timestamp 1698431365
transform 1 0 9296 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _264_
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _265_
timestamp 1698431365
transform 1 0 15232 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _266_
timestamp 1698431365
transform -1 0 32144 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _267_
timestamp 1698431365
transform -1 0 31920 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _268_
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _269_
timestamp 1698431365
transform 1 0 23408 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _270_
timestamp 1698431365
transform 1 0 27776 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _271_
timestamp 1698431365
transform 1 0 24976 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _272_
timestamp 1698431365
transform 1 0 28224 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _273_
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _274_
timestamp 1698431365
transform -1 0 28896 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _275_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _276_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _277_
timestamp 1698431365
transform 1 0 21952 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _278_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _279_
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _280_
timestamp 1698431365
transform 1 0 16464 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _281_
timestamp 1698431365
transform 1 0 15456 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _282_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _283_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _284_
timestamp 1698431365
transform 1 0 16576 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _285_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _286_
timestamp 1698431365
transform -1 0 28784 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _287_
timestamp 1698431365
transform -1 0 30128 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _288_
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _289_
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _290_
timestamp 1698431365
transform 1 0 28560 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _291_
timestamp 1698431365
transform -1 0 31360 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _292_
timestamp 1698431365
transform 1 0 24976 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _293_
timestamp 1698431365
transform 1 0 22624 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _294_
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _295_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _296_
timestamp 1698431365
transform -1 0 28896 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _297_
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _298_
timestamp 1698431365
transform -1 0 24976 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _299_
timestamp 1698431365
transform 1 0 18256 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _300_
timestamp 1698431365
transform -1 0 28672 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _301_
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _302_
timestamp 1698431365
transform 1 0 15904 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _303_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _304_
timestamp 1698431365
transform -1 0 23520 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _305_
timestamp 1698431365
transform 1 0 17136 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _306_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _307_
timestamp 1698431365
transform -1 0 5376 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _308_
timestamp 1698431365
transform -1 0 5376 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _309_
timestamp 1698431365
transform -1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _310_
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _311_
timestamp 1698431365
transform 1 0 3472 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _312_
timestamp 1698431365
transform -1 0 13216 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _313_
timestamp 1698431365
transform 1 0 7616 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _314_
timestamp 1698431365
transform -1 0 15568 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _315_
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _316_
timestamp 1698431365
transform -1 0 26544 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _317_
timestamp 1698431365
transform -1 0 25984 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _318_
timestamp 1698431365
transform 1 0 20384 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _319_
timestamp 1698431365
transform 1 0 18256 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _320_
timestamp 1698431365
transform 1 0 16016 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _321_
timestamp 1698431365
transform 1 0 13216 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _322_
timestamp 1698431365
transform -1 0 23184 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _323_
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _324_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _325_
timestamp 1698431365
transform 1 0 13216 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _326_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _327_
timestamp 1698431365
transform -1 0 12544 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _328_
timestamp 1698431365
transform 1 0 11536 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _329_
timestamp 1698431365
transform 1 0 9296 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _330_
timestamp 1698431365
transform -1 0 11872 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _331_
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _332_
timestamp 1698431365
transform -1 0 8176 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _333_
timestamp 1698431365
transform -1 0 8176 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _334_
timestamp 1698431365
transform 1 0 4368 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _335_
timestamp 1698431365
transform -1 0 7952 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _336_
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _337_
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _338_
timestamp 1698431365
transform 1 0 10192 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _339_
timestamp 1698431365
transform 1 0 8512 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _340_
timestamp 1698431365
transform -1 0 18256 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _341_
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _368_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _369_
timestamp 1698431365
transform 1 0 17584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _370_
timestamp 1698431365
transform -1 0 15120 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _371_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _372_
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _373_
timestamp 1698431365
transform 1 0 12320 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _375_
timestamp 1698431365
transform -1 0 10864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _376_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _377_
timestamp 1698431365
transform -1 0 17920 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _378_
timestamp 1698431365
transform 1 0 24192 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _379_
timestamp 1698431365
transform 1 0 1792 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_
timestamp 1698431365
transform 1 0 1904 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1698431365
transform 1 0 1792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _382_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1698431365
transform -1 0 26544 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _384_
timestamp 1698431365
transform -1 0 2464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1698431365
transform 1 0 22624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1698431365
transform -1 0 10080 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1698431365
transform -1 0 17920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1698431365
transform -1 0 6048 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1698431365
transform -1 0 16800 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _391_
timestamp 1698431365
transform -1 0 8848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1698431365
transform 1 0 1792 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _393_
timestamp 1698431365
transform 1 0 21392 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1698431365
transform -1 0 17920 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _395_
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1698431365
transform -1 0 10080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1698431365
transform -1 0 12656 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1698431365
transform 1 0 21280 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _400_
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1698431365
transform 1 0 9744 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1698431365
transform -1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1698431365
transform 1 0 12320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1698431365
transform -1 0 14112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__I
timestamp 1698431365
transform -1 0 6384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__I
timestamp 1698431365
transform 1 0 18816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1698431365
transform 1 0 15344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__I
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1698431365
transform 1 0 12768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1698431365
transform 1 0 6944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__I
timestamp 1698431365
transform -1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__I
timestamp 1698431365
transform -1 0 7056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__I
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I
timestamp 1698431365
transform 1 0 14336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__I
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I
timestamp 1698431365
transform 1 0 24640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__I
timestamp 1698431365
transform -1 0 17808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1698431365
transform 1 0 21840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1698431365
transform 1 0 22288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1698431365
transform -1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__I
timestamp 1698431365
transform 1 0 19376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__I
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__I
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__I
timestamp 1698431365
transform 1 0 27552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__I
timestamp 1698431365
transform 1 0 29792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__I
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__I
timestamp 1698431365
transform 1 0 32032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1698431365
transform 1 0 27552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__I
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__I
timestamp 1698431365
transform 1 0 22736 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1698431365
transform -1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1698431365
transform -1 0 26208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1698431365
transform 1 0 32032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1698431365
transform 1 0 31472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1698431365
transform 1 0 32032 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1698431365
transform 1 0 28112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__I
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I
timestamp 1698431365
transform 1 0 6384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I
timestamp 1698431365
transform -1 0 2016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__I
timestamp 1698431365
transform 1 0 16240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I
timestamp 1698431365
transform 1 0 25312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I
timestamp 1698431365
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__I
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__I
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__I
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I
timestamp 1698431365
transform 1 0 8512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__I
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I
timestamp 1698431365
transform 1 0 4144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I
timestamp 1698431365
transform -1 0 4704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__I
timestamp 1698431365
transform 1 0 5712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__I
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I
timestamp 1698431365
transform -1 0 11424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__I
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__I
timestamp 1698431365
transform 1 0 11984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I
timestamp 1698431365
transform 1 0 17472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__I
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698431365
transform 1 0 18032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698431365
transform -1 0 14672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698431365
transform 1 0 14896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698431365
transform 1 0 11872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698431365
transform 1 0 5040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__RN
timestamp 1698431365
transform -1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698431365
transform 1 0 10304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698431365
transform -1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__RN
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698431365
transform 1 0 16128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698431365
transform 1 0 12320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698431365
transform 1 0 9968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698431365
transform 1 0 4592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698431365
transform 1 0 8400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698431365
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698431365
transform 1 0 14672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698431365
transform 1 0 10752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__CLK
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__CLK
timestamp 1698431365
transform 1 0 29792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__CLK
timestamp 1698431365
transform -1 0 30016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__CLK
timestamp 1698431365
transform 1 0 29680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__CLK
timestamp 1698431365
transform 1 0 32032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__CLK
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__CLK
timestamp 1698431365
transform 1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__CLK
timestamp 1698431365
transform 1 0 29792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__CLK
timestamp 1698431365
transform 1 0 29568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__CLK
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__CLK
timestamp 1698431365
transform 1 0 14448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__CLK
timestamp 1698431365
transform -1 0 20832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__CLK
timestamp 1698431365
transform 1 0 29232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__CLK
timestamp 1698431365
transform 1 0 29792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__CLK
timestamp 1698431365
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__CLK
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__CLK
timestamp 1698431365
transform 1 0 19936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__CLK
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__CLK
timestamp 1698431365
transform 1 0 22176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__CLK
timestamp 1698431365
transform 1 0 7392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__CLK
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__CLK
timestamp 1698431365
transform 1 0 4592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__CLK
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__CLK
timestamp 1698431365
transform -1 0 7056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__CLK
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__CLK
timestamp 1698431365
transform 1 0 11648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__CLK
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__CLK
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__CLK
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__CLK
timestamp 1698431365
transform -1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__CLK
timestamp 1698431365
transform 1 0 12432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__CLK
timestamp 1698431365
transform 1 0 9520 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__CLK
timestamp 1698431365
transform 1 0 6160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__CLK
timestamp 1698431365
transform -1 0 11424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__CLK
timestamp 1698431365
transform 1 0 7952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__CLK
timestamp 1698431365
transform 1 0 8624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__CLK
timestamp 1698431365
transform 1 0 18480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__I
timestamp 1698431365
transform -1 0 21056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__I
timestamp 1698431365
transform 1 0 5040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__I
timestamp 1698431365
transform -1 0 4704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__I
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_prog_clk_I
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_prog_clk_I
timestamp 1698431365
transform -1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_prog_clk_I
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_prog_clk_I
timestamp 1698431365
transform 1 0 12432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_prog_clk_I
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_prog_clk_I
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_prog_clk_I
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_prog_clk_I
timestamp 1698431365
transform 1 0 25760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_prog_clk_I
timestamp 1698431365
transform -1 0 25536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 14112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 29232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 12208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 23408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 14000 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 17136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 3920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 4592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 19040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 17808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 10080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 26208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 18256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 24416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 22400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 10192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1698431365
transform 1 0 3808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1698431365
transform -1 0 7056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1698431365
transform 1 0 32144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698431365
transform -1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698431365
transform -1 0 2016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output62_I
timestamp 1698431365
transform 1 0 4144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1698431365
transform -1 0 4816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output70_I
timestamp 1698431365
transform -1 0 2016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1698431365
transform -1 0 12432 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1698431365
transform -1 0 16464 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1698431365
transform -1 0 27664 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_8 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_27
timestamp 1698431365
transform 1 0 4368 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_30
timestamp 1698431365
transform 1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_42
timestamp 1698431365
transform 1 0 6048 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_88 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_92
timestamp 1698431365
transform 1 0 11648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_94
timestamp 1698431365
transform 1 0 11872 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_110
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_114
timestamp 1698431365
transform 1 0 14112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_116
timestamp 1698431365
transform 1 0 14336 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_140
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_143
timestamp 1698431365
transform 1 0 17360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_163
timestamp 1698431365
transform 1 0 19600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_182
timestamp 1698431365
transform 1 0 21728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_200
timestamp 1698431365
transform 1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_214
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_225
timestamp 1698431365
transform 1 0 26544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_227
timestamp 1698431365
transform 1 0 26768 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_246 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_276
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_42
timestamp 1698431365
transform 1 0 6048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_44
timestamp 1698431365
transform 1 0 6272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_61
timestamp 1698431365
transform 1 0 8176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_65
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_74
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_91
timestamp 1698431365
transform 1 0 11536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_93
timestamp 1698431365
transform 1 0 11760 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_96
timestamp 1698431365
transform 1 0 12096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698431365
transform 1 0 17472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_147
timestamp 1698431365
transform 1 0 17808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_187
timestamp 1698431365
transform 1 0 22288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_189
timestamp 1698431365
transform 1 0 22512 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_225
timestamp 1698431365
transform 1 0 26544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_4
timestamp 1698431365
transform 1 0 1792 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_21
timestamp 1698431365
transform 1 0 3696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_25
timestamp 1698431365
transform 1 0 4144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_47
timestamp 1698431365
transform 1 0 6608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_202
timestamp 1698431365
transform 1 0 23968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_206
timestamp 1698431365
transform 1 0 24416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_236
timestamp 1698431365
transform 1 0 27776 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_251
timestamp 1698431365
transform 1 0 29456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_253
timestamp 1698431365
transform 1 0 29680 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_272
timestamp 1698431365
transform 1 0 31808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_276
timestamp 1698431365
transform 1 0 32256 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_22
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_78
timestamp 1698431365
transform 1 0 10080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_80
timestamp 1698431365
transform 1 0 10304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_115
timestamp 1698431365
transform 1 0 14224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_119
timestamp 1698431365
transform 1 0 14672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_123
timestamp 1698431365
transform 1 0 15120 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_176
timestamp 1698431365
transform 1 0 21056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_178
timestamp 1698431365
transform 1 0 21280 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_201
timestamp 1698431365
transform 1 0 23856 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_232
timestamp 1698431365
transform 1 0 27328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_236
timestamp 1698431365
transform 1 0 27776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_240
timestamp 1698431365
transform 1 0 28224 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 2240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_26
timestamp 1698431365
transform 1 0 4256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_30
timestamp 1698431365
transform 1 0 4704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_43
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_78
timestamp 1698431365
transform 1 0 10080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_82
timestamp 1698431365
transform 1 0 10528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_86
timestamp 1698431365
transform 1 0 10976 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_113
timestamp 1698431365
transform 1 0 14000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_117
timestamp 1698431365
transform 1 0 14448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_121
timestamp 1698431365
transform 1 0 14896 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_141
timestamp 1698431365
transform 1 0 17136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_149
timestamp 1698431365
transform 1 0 18032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_153
timestamp 1698431365
transform 1 0 18480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_184
timestamp 1698431365
transform 1 0 21952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_188
timestamp 1698431365
transform 1 0 22400 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_192
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_209
timestamp 1698431365
transform 1 0 24752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_276
timestamp 1698431365
transform 1 0 32256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_10
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_86
timestamp 1698431365
transform 1 0 10976 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_121
timestamp 1698431365
transform 1 0 14896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_125
timestamp 1698431365
transform 1 0 15344 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_203
timestamp 1698431365
transform 1 0 24080 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_237
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_239
timestamp 1698431365
transform 1 0 28112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_274
timestamp 1698431365
transform 1 0 32032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_30
timestamp 1698431365
transform 1 0 4704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_251
timestamp 1698431365
transform 1 0 29456 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_276
timestamp 1698431365
transform 1 0 32256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_78
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_82
timestamp 1698431365
transform 1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_86
timestamp 1698431365
transform 1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_185
timestamp 1698431365
transform 1 0 22064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_189
timestamp 1698431365
transform 1 0 22512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_191
timestamp 1698431365
transform 1 0 22736 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_232
timestamp 1698431365
transform 1 0 27328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_26
timestamp 1698431365
transform 1 0 4256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_39
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_164
timestamp 1698431365
transform 1 0 19712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_253
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_272
timestamp 1698431365
transform 1 0 31808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_274
timestamp 1698431365
transform 1 0 32032 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_152
timestamp 1698431365
transform 1 0 18368 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_160
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_163
timestamp 1698431365
transform 1 0 19600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_181
timestamp 1698431365
transform 1 0 21616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_185
timestamp 1698431365
transform 1 0 22064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_189
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_214
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_255
timestamp 1698431365
transform 1 0 29904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_273
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_30
timestamp 1698431365
transform 1 0 4704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_51
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_55
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_161
timestamp 1698431365
transform 1 0 19376 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_272
timestamp 1698431365
transform 1 0 31808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_276
timestamp 1698431365
transform 1 0 32256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_42
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_44
timestamp 1698431365
transform 1 0 6272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_61
timestamp 1698431365
transform 1 0 8176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_65
timestamp 1698431365
transform 1 0 8624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_110
timestamp 1698431365
transform 1 0 13664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_114
timestamp 1698431365
transform 1 0 14112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_118
timestamp 1698431365
transform 1 0 14560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_182
timestamp 1698431365
transform 1 0 21728 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_207
timestamp 1698431365
transform 1 0 24528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_246
timestamp 1698431365
transform 1 0 28896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_250
timestamp 1698431365
transform 1 0 29344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_254
timestamp 1698431365
transform 1 0 29792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_256
timestamp 1698431365
transform 1 0 30016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_16
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_48
timestamp 1698431365
transform 1 0 6720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_52
timestamp 1698431365
transform 1 0 7168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_56
timestamp 1698431365
transform 1 0 7616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_58
timestamp 1698431365
transform 1 0 7840 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_75
timestamp 1698431365
transform 1 0 9744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_79
timestamp 1698431365
transform 1 0 10192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_96
timestamp 1698431365
transform 1 0 12096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_98
timestamp 1698431365
transform 1 0 12320 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_127
timestamp 1698431365
transform 1 0 15568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_152
timestamp 1698431365
transform 1 0 18368 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_155
timestamp 1698431365
transform 1 0 18704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_263
timestamp 1698431365
transform 1 0 30800 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_271
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_275
timestamp 1698431365
transform 1 0 32144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_100
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_154
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_197
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_272
timestamp 1698431365
transform 1 0 31808 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_28
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_218
timestamp 1698431365
transform 1 0 25760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_226
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_253
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_272
timestamp 1698431365
transform 1 0 31808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_276
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_36
timestamp 1698431365
transform 1 0 5376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_38
timestamp 1698431365
transform 1 0 5600 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_63
timestamp 1698431365
transform 1 0 8400 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_90
timestamp 1698431365
transform 1 0 11424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_92
timestamp 1698431365
transform 1 0 11648 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_186
timestamp 1698431365
transform 1 0 22176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_218
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_222
timestamp 1698431365
transform 1 0 26208 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_47
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_125
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_251
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_253
timestamp 1698431365
transform 1 0 29680 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_272
timestamp 1698431365
transform 1 0 31808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_276
timestamp 1698431365
transform 1 0 32256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_135
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_250
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_254
timestamp 1698431365
transform 1 0 29792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_51
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_90
timestamp 1698431365
transform 1 0 11424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_94
timestamp 1698431365
transform 1 0 11872 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_131
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_135
timestamp 1698431365
transform 1 0 16464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_170
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_189
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_234
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_255
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_272
timestamp 1698431365
transform 1 0 31808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_276
timestamp 1698431365
transform 1 0 32256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_16
timestamp 1698431365
transform 1 0 3136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_148
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_186
timestamp 1698431365
transform 1 0 22176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_274
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_71
timestamp 1698431365
transform 1 0 9296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_96
timestamp 1698431365
transform 1 0 12096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_98
timestamp 1698431365
transform 1 0 12320 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_151
timestamp 1698431365
transform 1 0 18256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_167
timestamp 1698431365
transform 1 0 20048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_272
timestamp 1698431365
transform 1 0 31808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_276
timestamp 1698431365
transform 1 0 32256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_94
timestamp 1698431365
transform 1 0 11872 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_131
timestamp 1698431365
transform 1 0 16016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_171
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_173
timestamp 1698431365
transform 1 0 20720 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_192
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_250
timestamp 1698431365
transform 1 0 29344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_258
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_275
timestamp 1698431365
transform 1 0 32144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_30
timestamp 1698431365
transform 1 0 4704 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_47
timestamp 1698431365
transform 1 0 6608 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_113
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_117
timestamp 1698431365
transform 1 0 14448 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_156
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_160
timestamp 1698431365
transform 1 0 19264 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_228
timestamp 1698431365
transform 1 0 26880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_230
timestamp 1698431365
transform 1 0 27104 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_267
timestamp 1698431365
transform 1 0 31248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_271
timestamp 1698431365
transform 1 0 31696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_275
timestamp 1698431365
transform 1 0 32144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_4
timestamp 1698431365
transform 1 0 1792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_27
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_31
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_35
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_185
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_189
timestamp 1698431365
transform 1 0 22512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_193
timestamp 1698431365
transform 1 0 22960 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_246
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_254
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_30
timestamp 1698431365
transform 1 0 4704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_127
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_129
timestamp 1698431365
transform 1 0 15792 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_164
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_255
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_272
timestamp 1698431365
transform 1 0 31808 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_276
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_22
timestamp 1698431365
transform 1 0 3808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_24
timestamp 1698431365
transform 1 0 4032 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_78
timestamp 1698431365
transform 1 0 10080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_262
timestamp 1698431365
transform 1 0 30688 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_39
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_62
timestamp 1698431365
transform 1 0 8288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_64
timestamp 1698431365
transform 1 0 8512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_67
timestamp 1698431365
transform 1 0 8848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_276
timestamp 1698431365
transform 1 0 32256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_16
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_63
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_82
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_86
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_90
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_137
timestamp 1698431365
transform 1 0 16688 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_154
timestamp 1698431365
transform 1 0 18592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_163
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_59
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_122
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_126
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_150
timestamp 1698431365
transform 1 0 18144 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_158
timestamp 1698431365
transform 1 0 19040 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_184
timestamp 1698431365
transform 1 0 21952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_188
timestamp 1698431365
transform 1 0 22400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_209
timestamp 1698431365
transform 1 0 24752 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_272
timestamp 1698431365
transform 1 0 31808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_4
timestamp 1698431365
transform 1 0 1792 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_27
timestamp 1698431365
transform 1 0 4368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_31
timestamp 1698431365
transform 1 0 4816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_35
timestamp 1698431365
transform 1 0 5264 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_74
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_97
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_103
timestamp 1698431365
transform 1 0 12880 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_148
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_201
timestamp 1698431365
transform 1 0 23856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_237
timestamp 1698431365
transform 1 0 27888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_30
timestamp 1698431365
transform 1 0 4704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_57
timestamp 1698431365
transform 1 0 7728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_61
timestamp 1698431365
transform 1 0 8176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_63
timestamp 1698431365
transform 1 0 8400 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_125
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_129
timestamp 1698431365
transform 1 0 15792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_183
timestamp 1698431365
transform 1 0 21840 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_252
timestamp 1698431365
transform 1 0 29568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_260
timestamp 1698431365
transform 1 0 30464 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_61
timestamp 1698431365
transform 1 0 8176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_63
timestamp 1698431365
transform 1 0 8400 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_26
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_71
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_75
timestamp 1698431365
transform 1 0 9744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_79
timestamp 1698431365
transform 1 0 10192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_87
timestamp 1698431365
transform 1 0 11088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_187
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_239
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_276
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_23
timestamp 1698431365
transform 1 0 3920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_61
timestamp 1698431365
transform 1 0 8176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_63
timestamp 1698431365
transform 1 0 8400 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_86
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_106 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_122
timestamp 1698431365
transform 1 0 15008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_152
timestamp 1698431365
transform 1 0 18368 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_237
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_241
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_245
timestamp 1698431365
transform 1 0 28784 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_262
timestamp 1698431365
transform 1 0 30688 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_273
timestamp 1698431365
transform 1 0 31920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_20
timestamp 1698431365
transform 1 0 3584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_36
timestamp 1698431365
transform 1 0 5376 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_43
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_47
timestamp 1698431365
transform 1 0 6608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_51
timestamp 1698431365
transform 1 0 7056 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_70
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_93
timestamp 1698431365
transform 1 0 11760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_119
timestamp 1698431365
transform 1 0 14672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_138
timestamp 1698431365
transform 1 0 16800 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_146
timestamp 1698431365
transform 1 0 17696 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_169
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_203
timestamp 1698431365
transform 1 0 24080 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_206
timestamp 1698431365
transform 1 0 24416 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_221
timestamp 1698431365
transform 1 0 26096 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_237
timestamp 1698431365
transform 1 0 27888 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_240
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_274
timestamp 1698431365
transform 1 0 32032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_276
timestamp 1698431365
transform 1 0 32256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform 1 0 11424 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 19600 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 31696 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform 1 0 2576 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform -1 0 31808 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 4368 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 16464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 18144 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 20048 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 30688 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform -1 0 31808 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 27888 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform 1 0 7504 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 32144 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 20832 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform -1 0 27888 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform 1 0 9744 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 13216 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 24528 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 21616 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold26
timestamp 1698431365
transform 1 0 6384 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform -1 0 32368 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold30
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 24752 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 24528 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold34
timestamp 1698431365
transform -1 0 31808 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform -1 0 28560 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform 1 0 2576 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 31696 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 20048 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold42
timestamp 1698431365
transform 1 0 10304 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform -1 0 23408 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold46
timestamp 1698431365
transform -1 0 12880 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform -1 0 8176 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform -1 0 20048 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold50
timestamp 1698431365
transform 1 0 25984 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform -1 0 27888 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform -1 0 22848 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold54
timestamp 1698431365
transform -1 0 3696 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform 1 0 10416 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold58
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform -1 0 31808 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold62
timestamp 1698431365
transform 1 0 25984 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 27888 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform -1 0 16464 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 27552 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold67
timestamp 1698431365
transform -1 0 31808 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold68
timestamp 1698431365
transform 1 0 6384 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold69
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold70
timestamp 1698431365
transform -1 0 31920 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold71
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold72
timestamp 1698431365
transform -1 0 19600 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold73
timestamp 1698431365
transform -1 0 18144 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold74
timestamp 1698431365
transform -1 0 31808 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold75
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold76
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold77
timestamp 1698431365
transform -1 0 8176 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold78
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold79
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold80
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold81
timestamp 1698431365
transform 1 0 9968 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold82
timestamp 1698431365
transform 1 0 6496 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold83
timestamp 1698431365
transform -1 0 8960 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold84
timestamp 1698431365
transform 1 0 22064 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold85
timestamp 1698431365
transform -1 0 31808 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold86
timestamp 1698431365
transform -1 0 31808 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold87
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold88
timestamp 1698431365
transform -1 0 20384 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold89
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold90
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold91
timestamp 1698431365
transform -1 0 16576 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold92
timestamp 1698431365
transform -1 0 17136 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold93
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold94
timestamp 1698431365
transform -1 0 8512 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold95
timestamp 1698431365
transform -1 0 31808 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold96
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold97
timestamp 1698431365
transform -1 0 31808 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold98
timestamp 1698431365
transform -1 0 31808 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold99
timestamp 1698431365
transform -1 0 9744 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold100
timestamp 1698431365
transform -1 0 31808 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold101
timestamp 1698431365
transform 1 0 2352 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold102
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold103
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold104
timestamp 1698431365
transform -1 0 31808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold105
timestamp 1698431365
transform -1 0 31808 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 15120 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1792 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 26096 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 9968 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 13664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 21952 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 23072 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 13776 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 16352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 32256 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 16800 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 23520 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 1904 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 19712 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 18256 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 8176 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 1792 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 30800 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 20272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 17360 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 6048 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 21280 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 17920 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 18592 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 2464 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32368 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output39
timestamp 1698431365
transform -1 0 7056 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output40
timestamp 1698431365
transform 1 0 24976 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42
timestamp 1698431365
transform -1 0 3136 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform 1 0 30800 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform -1 0 5152 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform -1 0 7504 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform 1 0 30800 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output49
timestamp 1698431365
transform -1 0 28112 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output50
timestamp 1698431365
transform -1 0 7056 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output51
timestamp 1698431365
transform 1 0 22848 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698431365
transform 1 0 2800 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform -1 0 25984 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output54
timestamp 1698431365
transform -1 0 10528 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output55
timestamp 1698431365
transform 1 0 3136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output56
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output57 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3136 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform 1 0 22624 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output60
timestamp 1698431365
transform -1 0 8176 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698431365
transform -1 0 10976 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output62
timestamp 1698431365
transform -1 0 2800 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output63
timestamp 1698431365
transform 1 0 27216 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output64
timestamp 1698431365
transform -1 0 3136 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform 1 0 23296 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output68
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output69
timestamp 1698431365
transform -1 0 3136 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output70
timestamp 1698431365
transform -1 0 3136 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output71
timestamp 1698431365
transform -1 0 14896 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_35 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_36
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 32592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_37
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 32592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_38
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 32592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_39
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 32592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_40
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 32592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_41
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 32592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_42
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 32592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_43
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 32592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 32592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 32592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 32592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 32592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 32592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 32592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 32592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 32592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 32592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 32592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 32592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 32592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 32592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 32592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 32592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 32592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 32592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 32592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 32592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 32592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 32592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 32592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 32592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 32592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 32592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__73
timestamp 1698431365
transform -1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__74
timestamp 1698431365
transform 1 0 31920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__75
timestamp 1698431365
transform -1 0 9856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__76
timestamp 1698431365
transform -1 0 32256 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__77
timestamp 1698431365
transform 1 0 4816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__78
timestamp 1698431365
transform 1 0 31808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__79
timestamp 1698431365
transform 1 0 26544 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__80
timestamp 1698431365
transform -1 0 12992 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__81
timestamp 1698431365
transform -1 0 12992 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__82
timestamp 1698431365
transform 1 0 29120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__83
timestamp 1698431365
transform -1 0 6832 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__84
timestamp 1698431365
transform -1 0 7056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__85
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__86
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__87
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__88
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__89
timestamp 1698431365
transform -1 0 19376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__90
timestamp 1698431365
transform 1 0 31920 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__91
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__92
timestamp 1698431365
transform 1 0 31808 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__93
timestamp 1698431365
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__94
timestamp 1698431365
transform -1 0 8400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__95
timestamp 1698431365
transform 1 0 3136 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__96
timestamp 1698431365
transform -1 0 12320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  sb_0__1__97
timestamp 1698431365
transform -1 0 24864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_71
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_72
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_73
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_74
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_75
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_76
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_77
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_78
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_79
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_80
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_81
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_82
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_83
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_84
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_85
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_86
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_87
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_88
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_89
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_90
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_91
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_92
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_93
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_94
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_95
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_96
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_97
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_98
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_99
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_100
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_101
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_102
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_103
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_104
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_105
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_113
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_114
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_115
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_116
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_117
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_118
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_119
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_120
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_121
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_122
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_123
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_124
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_125
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_126
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_127
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_128
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_129
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_130
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_131
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_132
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_133
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_134
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_135
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_136
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_137
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_138
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_139
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_140
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_141
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_142
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_143
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_144
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_145
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_146
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_147
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_148
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_149
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_150
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_151
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_152
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_153
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_154
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_155
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_156
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_157
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_158
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_159
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_160
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_161
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_162
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_163
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_164
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_165
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_166
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_167
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_168
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_169
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_170
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_171
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_172
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_173
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_174
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_175
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_176
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_177
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_178
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_179
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_180
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_181
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_182
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_183
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_184
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_185
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_186
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_187
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_188
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_189
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_190
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_191
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_192
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_193
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_194
timestamp 1698431365
transform 1 0 8960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_195
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_196
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_197
timestamp 1698431365
transform 1 0 20384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_198
timestamp 1698431365
transform 1 0 24192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_199
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_200
timestamp 1698431365
transform 1 0 31808 0 1 29792
box -86 -86 310 870
<< labels >>
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 1 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 2 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 3 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 4 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 5 nsew signal input
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 ccff_head
port 6 nsew signal input
flabel metal3 s 33200 22848 34000 22960 0 FreeSans 448 0 0 0 ccff_tail
port 7 nsew signal tristate
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 chanx_right_in[0]
port 8 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 chanx_right_in[10]
port 9 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 chanx_right_in[11]
port 10 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 chanx_right_in[12]
port 11 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 chanx_right_in[13]
port 12 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 chanx_right_in[14]
port 13 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 chanx_right_in[15]
port 14 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 chanx_right_in[16]
port 15 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 chanx_right_in[17]
port 16 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 chanx_right_in[18]
port 17 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 chanx_right_in[19]
port 18 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 chanx_right_in[1]
port 19 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 chanx_right_in[2]
port 20 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 chanx_right_in[3]
port 21 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 chanx_right_in[4]
port 22 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 chanx_right_in[5]
port 23 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 chanx_right_in[6]
port 24 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 chanx_right_in[7]
port 25 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 chanx_right_in[8]
port 26 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 chanx_right_in[9]
port 27 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 chanx_right_out[0]
port 28 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 chanx_right_out[10]
port 29 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 chanx_right_out[11]
port 30 nsew signal tristate
flabel metal2 s 8736 33200 8848 34000 0 FreeSans 448 90 0 0 chanx_right_out[12]
port 31 nsew signal tristate
flabel metal3 s 0 2016 800 2128 0 FreeSans 448 0 0 0 chanx_right_out[13]
port 32 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 chanx_right_out[14]
port 33 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 chanx_right_out[15]
port 34 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 chanx_right_out[16]
port 35 nsew signal tristate
flabel metal2 s 24864 33200 24976 34000 0 FreeSans 448 90 0 0 chanx_right_out[17]
port 36 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 chanx_right_out[18]
port 37 nsew signal tristate
flabel metal3 s 33200 27552 34000 27664 0 FreeSans 448 0 0 0 chanx_right_out[19]
port 38 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 chanx_right_out[1]
port 39 nsew signal tristate
flabel metal2 s 9408 33200 9520 34000 0 FreeSans 448 90 0 0 chanx_right_out[2]
port 40 nsew signal tristate
flabel metal2 s 672 33200 784 34000 0 FreeSans 448 90 0 0 chanx_right_out[3]
port 41 nsew signal tristate
flabel metal3 s 33200 31584 34000 31696 0 FreeSans 448 0 0 0 chanx_right_out[4]
port 42 nsew signal tristate
flabel metal3 s 33200 672 34000 784 0 FreeSans 448 0 0 0 chanx_right_out[5]
port 43 nsew signal tristate
flabel metal2 s 8064 33200 8176 34000 0 FreeSans 448 90 0 0 chanx_right_out[6]
port 44 nsew signal tristate
flabel metal3 s 33200 25536 34000 25648 0 FreeSans 448 0 0 0 chanx_right_out[7]
port 45 nsew signal tristate
flabel metal2 s 18816 33200 18928 34000 0 FreeSans 448 90 0 0 chanx_right_out[8]
port 46 nsew signal tristate
flabel metal2 s 28224 33200 28336 34000 0 FreeSans 448 90 0 0 chanx_right_out[9]
port 47 nsew signal tristate
flabel metal2 s 12768 33200 12880 34000 0 FreeSans 448 90 0 0 chany_bottom_in[0]
port 48 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 chany_bottom_in[10]
port 49 nsew signal input
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 chany_bottom_in[11]
port 50 nsew signal input
flabel metal2 s 15456 33200 15568 34000 0 FreeSans 448 90 0 0 chany_bottom_in[12]
port 51 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 chany_bottom_in[13]
port 52 nsew signal input
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 chany_bottom_in[14]
port 53 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 chany_bottom_in[15]
port 54 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 chany_bottom_in[16]
port 55 nsew signal input
flabel metal3 s 33200 30912 34000 31024 0 FreeSans 448 0 0 0 chany_bottom_in[17]
port 56 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 chany_bottom_in[18]
port 57 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 chany_bottom_in[19]
port 58 nsew signal input
flabel metal2 s 16128 33200 16240 34000 0 FreeSans 448 90 0 0 chany_bottom_in[1]
port 59 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 chany_bottom_in[2]
port 60 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 chany_bottom_in[3]
port 61 nsew signal input
flabel metal3 s 33200 28224 34000 28336 0 FreeSans 448 0 0 0 chany_bottom_in[4]
port 62 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 chany_bottom_in[5]
port 63 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 chany_bottom_in[6]
port 64 nsew signal input
flabel metal2 s 25536 33200 25648 34000 0 FreeSans 448 90 0 0 chany_bottom_in[7]
port 65 nsew signal input
flabel metal2 s 2016 33200 2128 34000 0 FreeSans 448 90 0 0 chany_bottom_in[8]
port 66 nsew signal input
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 chany_bottom_in[9]
port 67 nsew signal input
flabel metal3 s 0 2688 800 2800 0 FreeSans 448 0 0 0 chany_bottom_out[0]
port 68 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 chany_bottom_out[10]
port 69 nsew signal tristate
flabel metal3 s 33200 7392 34000 7504 0 FreeSans 448 0 0 0 chany_bottom_out[11]
port 70 nsew signal tristate
flabel metal3 s 33200 4032 34000 4144 0 FreeSans 448 0 0 0 chany_bottom_out[12]
port 71 nsew signal tristate
flabel metal2 s 6720 33200 6832 34000 0 FreeSans 448 90 0 0 chany_bottom_out[13]
port 72 nsew signal tristate
flabel metal2 s 26880 33200 26992 34000 0 FreeSans 448 90 0 0 chany_bottom_out[14]
port 73 nsew signal tristate
flabel metal2 s 10080 33200 10192 34000 0 FreeSans 448 90 0 0 chany_bottom_out[15]
port 74 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 chany_bottom_out[16]
port 75 nsew signal tristate
flabel metal3 s 33200 26880 34000 26992 0 FreeSans 448 0 0 0 chany_bottom_out[17]
port 76 nsew signal tristate
flabel metal2 s 16800 33200 16912 34000 0 FreeSans 448 90 0 0 chany_bottom_out[18]
port 77 nsew signal tristate
flabel metal3 s 33200 6048 34000 6160 0 FreeSans 448 0 0 0 chany_bottom_out[19]
port 78 nsew signal tristate
flabel metal2 s 5376 33200 5488 34000 0 FreeSans 448 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal3 s 33200 5376 34000 5488 0 FreeSans 448 0 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 6048 33200 6160 34000 0 FreeSans 448 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal3 s 33200 4704 34000 4816 0 FreeSans 448 0 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal2 s 3360 33200 3472 34000 0 FreeSans 448 90 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal2 s 27552 33200 27664 34000 0 FreeSans 448 90 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 12096 33200 12208 34000 0 FreeSans 448 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal2 s 2688 33200 2800 34000 0 FreeSans 448 90 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal3 s 33200 2016 34000 2128 0 FreeSans 448 0 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal2 s 4032 33200 4144 34000 0 FreeSans 448 90 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal2 s 26208 33200 26320 34000 0 FreeSans 448 90 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal2 s 10752 33200 10864 34000 0 FreeSans 448 90 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal3 s 33200 26208 34000 26320 0 FreeSans 448 0 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 18144 33200 18256 34000 0 FreeSans 448 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal3 s 33200 6720 34000 6832 0 FreeSans 448 0 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 chany_top_in[19]
port 98 nsew signal input
flabel metal3 s 33200 1344 34000 1456 0 FreeSans 448 0 0 0 chany_top_in[1]
port 99 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 chany_top_in[2]
port 100 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 chany_top_in[3]
port 101 nsew signal input
flabel metal3 s 33200 3360 34000 3472 0 FreeSans 448 0 0 0 chany_top_in[4]
port 102 nsew signal input
flabel metal2 s 4704 33200 4816 34000 0 FreeSans 448 90 0 0 chany_top_in[5]
port 103 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 chany_top_in[6]
port 104 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 chany_top_in[7]
port 105 nsew signal input
flabel metal2 s 11424 33200 11536 34000 0 FreeSans 448 90 0 0 chany_top_in[8]
port 106 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 chany_top_in[9]
port 107 nsew signal input
flabel metal2 s 28896 33200 29008 34000 0 FreeSans 448 90 0 0 chany_top_out[0]
port 108 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 chany_top_out[10]
port 109 nsew signal tristate
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 chany_top_out[11]
port 110 nsew signal tristate
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 chany_top_out[12]
port 111 nsew signal tristate
flabel metal2 s 14784 33200 14896 34000 0 FreeSans 448 90 0 0 chany_top_out[13]
port 112 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 chany_top_out[14]
port 113 nsew signal tristate
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 chany_top_out[15]
port 114 nsew signal tristate
flabel metal3 s 33200 30240 34000 30352 0 FreeSans 448 0 0 0 chany_top_out[16]
port 115 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 chany_top_out[17]
port 116 nsew signal tristate
flabel metal3 s 33200 29568 34000 29680 0 FreeSans 448 0 0 0 chany_top_out[18]
port 117 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 chany_top_out[19]
port 118 nsew signal tristate
flabel metal2 s 14112 33200 14224 34000 0 FreeSans 448 90 0 0 chany_top_out[1]
port 119 nsew signal tristate
flabel metal2 s 17472 33200 17584 34000 0 FreeSans 448 90 0 0 chany_top_out[2]
port 120 nsew signal tristate
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 chany_top_out[3]
port 121 nsew signal tristate
flabel metal2 s 7392 33200 7504 34000 0 FreeSans 448 90 0 0 chany_top_out[4]
port 122 nsew signal tristate
flabel metal3 s 33200 28896 34000 29008 0 FreeSans 448 0 0 0 chany_top_out[5]
port 123 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 chany_top_out[6]
port 124 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 chany_top_out[7]
port 125 nsew signal tristate
flabel metal3 s 33200 2688 34000 2800 0 FreeSans 448 0 0 0 chany_top_out[8]
port 126 nsew signal tristate
flabel metal2 s 1344 33200 1456 34000 0 FreeSans 448 90 0 0 chany_top_out[9]
port 127 nsew signal tristate
flabel metal2 s 13440 33200 13552 34000 0 FreeSans 448 90 0 0 pReset
port 128 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 prog_clk
port 129 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 130 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 131 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 132 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 133 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 137 nsew signal input
flabel metal3 s 33200 8064 34000 8176 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 138 nsew signal input
flabel metal3 s 33200 0 34000 112 0 FreeSans 448 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 139 nsew signal input
flabel metal4 s 5090 3076 5410 30636 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 12902 3076 13222 30636 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 20714 3076 21034 30636 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 28526 3076 28846 30636 0 FreeSans 1280 90 0 0 vdd
port 140 nsew power bidirectional
flabel metal4 s 8996 3076 9316 30636 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
flabel metal4 s 16808 3076 17128 30636 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
flabel metal4 s 24620 3076 24940 30636 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
flabel metal4 s 32432 3076 32752 30636 0 FreeSans 1280 90 0 0 vss
port 141 nsew ground bidirectional
rlabel metal1 16968 30576 16968 30576 0 vdd
rlabel via1 17048 29792 17048 29792 0 vss
rlabel metal2 17416 5488 17416 5488 0 _000_
rlabel metal2 15512 4704 15512 4704 0 _001_
rlabel metal2 12824 5656 12824 5656 0 _002_
rlabel metal2 8792 4928 8792 4928 0 _003_
rlabel metal2 20328 4928 20328 4928 0 _004_
rlabel metal2 21336 5096 21336 5096 0 _005_
rlabel metal2 20552 5880 20552 5880 0 _006_
rlabel metal2 19656 5992 19656 5992 0 _007_
rlabel metal2 16072 14560 16072 14560 0 _008_
rlabel metal2 12488 13664 12488 13664 0 _009_
rlabel metal3 9464 15848 9464 15848 0 _010_
rlabel metal3 6888 15848 6888 15848 0 _011_
rlabel metal2 6216 13440 6216 13440 0 _012_
rlabel metal2 4760 12208 4760 12208 0 _013_
rlabel metal2 2408 11928 2408 11928 0 _014_
rlabel metal3 4088 13944 4088 13944 0 _015_
rlabel metal2 8344 9408 8344 9408 0 _016_
rlabel metal2 7448 6888 7448 6888 0 _017_
rlabel metal2 4536 9856 4536 9856 0 _018_
rlabel metal2 6216 11368 6216 11368 0 _019_
rlabel metal2 20888 7392 20888 7392 0 _020_
rlabel metal2 19768 5656 19768 5656 0 _021_
rlabel metal3 24864 8792 24864 8792 0 _022_
rlabel metal2 21224 9408 21224 9408 0 _023_
rlabel metal2 21448 9296 21448 9296 0 _024_
rlabel metal2 14840 8736 14840 8736 0 _025_
rlabel metal2 14168 7840 14168 7840 0 _026_
rlabel metal2 12488 8792 12488 8792 0 _027_
rlabel metal2 20440 11928 20440 11928 0 _028_
rlabel metal2 18144 9688 18144 9688 0 _029_
rlabel metal3 28784 10024 28784 10024 0 _030_
rlabel metal2 27720 4144 27720 4144 0 _031_
rlabel metal3 26656 9576 26656 9576 0 _032_
rlabel metal2 26488 9408 26488 9408 0 _033_
rlabel metal2 30856 12208 30856 12208 0 _034_
rlabel metal2 27944 11984 27944 11984 0 _035_
rlabel metal2 31136 7672 31136 7672 0 _036_
rlabel metal2 28504 6720 28504 6720 0 _037_
rlabel metal2 25928 12936 25928 12936 0 _038_
rlabel metal2 23128 10584 23128 10584 0 _039_
rlabel metal3 27496 17080 27496 17080 0 _040_
rlabel metal2 25144 14700 25144 14700 0 _041_
rlabel metal2 23576 15624 23576 15624 0 _042_
rlabel metal2 21560 16240 21560 16240 0 _043_
rlabel metal2 19880 14280 19880 14280 0 _044_
rlabel metal2 18088 15680 18088 15680 0 _045_
rlabel metal2 24360 18760 24360 18760 0 _046_
rlabel metal2 21336 18144 21336 18144 0 _047_
rlabel metal2 19544 18312 19544 18312 0 _048_
rlabel metal2 19432 16632 19432 16632 0 _049_
rlabel metal2 25592 16296 25592 16296 0 _050_
rlabel metal2 24696 16408 24696 16408 0 _051_
rlabel metal2 31472 18424 31472 18424 0 _052_
rlabel metal2 28504 20160 28504 20160 0 _053_
rlabel metal2 31808 16968 31808 16968 0 _054_
rlabel metal3 26796 18536 26796 18536 0 _055_
rlabel metal2 27384 18760 27384 18760 0 _056_
rlabel metal2 25704 17864 25704 17864 0 _057_
rlabel metal3 30240 28056 30240 28056 0 _058_
rlabel metal2 20552 21504 20552 21504 0 _059_
rlabel metal2 25704 22400 25704 22400 0 _060_
rlabel metal2 25704 20552 25704 20552 0 _061_
rlabel metal2 22120 21504 22120 21504 0 _062_
rlabel metal2 21168 21784 21168 21784 0 _063_
rlabel metal2 28392 27328 28392 27328 0 _064_
rlabel metal2 26600 24136 26600 24136 0 _065_
rlabel metal2 18984 22568 18984 22568 0 _066_
rlabel metal3 17248 23240 17248 23240 0 _067_
rlabel metal3 22120 24808 22120 24808 0 _068_
rlabel metal2 20328 23744 20328 23744 0 _069_
rlabel metal2 10696 17024 10696 17024 0 _070_
rlabel metal2 5880 21168 5880 21168 0 _071_
rlabel metal2 2128 15512 2128 15512 0 _072_
rlabel metal2 2296 17304 2296 17304 0 _073_
rlabel metal2 10920 16184 10920 16184 0 _074_
rlabel metal2 6272 15400 6272 15400 0 _075_
rlabel metal3 11200 17752 11200 17752 0 _076_
rlabel metal2 9912 18256 9912 18256 0 _077_
rlabel metal2 12600 16184 12600 16184 0 _078_
rlabel metal3 15204 16968 15204 16968 0 _079_
rlabel metal2 27496 29568 27496 29568 0 _080_
rlabel metal3 22400 26936 22400 26936 0 _081_
rlabel metal2 23352 28504 23352 28504 0 _082_
rlabel metal2 21336 26712 21336 26712 0 _083_
rlabel metal2 18984 25872 18984 25872 0 _084_
rlabel metal2 16408 26432 16408 26432 0 _085_
rlabel metal2 20216 29848 20216 29848 0 _086_
rlabel metal2 24360 28056 24360 28056 0 _087_
rlabel metal2 19992 27776 19992 27776 0 _088_
rlabel metal3 17248 26824 17248 26824 0 _089_
rlabel metal2 13720 27608 13720 27608 0 _090_
rlabel metal2 5992 29064 5992 29064 0 _091_
rlabel metal2 14728 24752 14728 24752 0 _092_
rlabel metal2 12544 23688 12544 23688 0 _093_
rlabel metal2 8904 25088 8904 25088 0 _094_
rlabel metal2 9576 23464 9576 23464 0 _095_
rlabel metal2 5376 27944 5376 27944 0 _096_
rlabel metal2 6272 29176 6272 29176 0 _097_
rlabel metal2 7448 24360 7448 24360 0 _098_
rlabel metal2 5992 24416 5992 24416 0 _099_
rlabel metal2 8568 21672 8568 21672 0 _100_
rlabel metal2 8456 21616 8456 21616 0 _101_
rlabel metal2 13440 20664 13440 20664 0 _102_
rlabel metal2 11480 21448 11480 21448 0 _103_
rlabel metal2 15288 19264 15288 19264 0 _104_
rlabel metal2 15400 21224 15400 21224 0 _105_
rlabel metal2 15176 24192 15176 24192 0 _106_
rlabel metal2 15344 7672 15344 7672 0 _107_
rlabel metal2 20216 4928 20216 4928 0 _108_
rlabel metal2 15176 11368 15176 11368 0 _109_
rlabel metal3 23408 5096 23408 5096 0 _110_
rlabel metal2 27552 6104 27552 6104 0 _111_
rlabel metal2 19656 15736 19656 15736 0 _112_
rlabel metal2 28168 29736 28168 29736 0 _113_
rlabel metal2 28168 27496 28168 27496 0 _114_
rlabel metal2 2072 19264 2072 19264 0 _115_
rlabel metal2 26936 29904 26936 29904 0 _116_
rlabel metal2 5656 29960 5656 29960 0 _117_
rlabel metal2 14840 9744 14840 9744 0 ccff_head
rlabel metal2 31528 22960 31528 22960 0 ccff_tail
rlabel metal2 24920 1190 24920 1190 0 chanx_right_out[15]
rlabel metal3 1302 30296 1302 30296 0 chanx_right_out[16]
rlabel metal3 25424 29960 25424 29960 0 chanx_right_out[17]
rlabel metal3 560 28728 560 28728 0 chanx_right_out[18]
rlabel metal2 4536 27776 4536 27776 0 chany_bottom_in[0]
rlabel metal2 25816 7000 25816 7000 0 chany_bottom_in[10]
rlabel metal3 2366 29624 2366 29624 0 chany_bottom_in[11]
rlabel metal3 10920 30072 10920 30072 0 chany_bottom_in[12]
rlabel metal3 9128 3528 9128 3528 0 chany_bottom_in[13]
rlabel metal3 2058 6104 2058 6104 0 chany_bottom_in[14]
rlabel metal3 23688 3528 23688 3528 0 chany_bottom_in[15]
rlabel metal2 3976 22008 3976 22008 0 chany_bottom_in[16]
rlabel metal2 29904 30968 29904 30968 0 chany_bottom_in[17]
rlabel metal3 1246 21560 1246 21560 0 chany_bottom_in[18]
rlabel metal3 13832 30184 13832 30184 0 chany_bottom_in[1]
rlabel metal2 26264 1638 26264 1638 0 chany_bottom_in[2]
rlabel metal3 1246 27608 1246 27608 0 chany_bottom_in[3]
rlabel metal3 30072 10080 30072 10080 0 chany_bottom_in[4]
rlabel metal2 16520 12096 16520 12096 0 chany_bottom_in[5]
rlabel metal2 1848 8232 1848 8232 0 chany_bottom_in[6]
rlabel metal2 24080 13944 24080 13944 0 chany_bottom_in[7]
rlabel metal2 2240 31920 2240 31920 0 chany_bottom_in[8]
rlabel metal2 18984 10360 18984 10360 0 chany_bottom_in[9]
rlabel metal2 2184 30576 2184 30576 0 chany_bottom_out[10]
rlabel metal2 31808 10360 31808 10360 0 chany_bottom_out[11]
rlabel metal3 5488 29960 5488 29960 0 chany_bottom_out[13]
rlabel metal2 27384 28728 27384 28728 0 chany_bottom_out[14]
rlabel metal2 6888 29008 6888 29008 0 chany_bottom_out[15]
rlabel metal2 31752 28112 31752 28112 0 chany_bottom_out[17]
rlabel metal2 17864 29456 17864 29456 0 chany_bottom_out[18]
rlabel metal2 27384 5152 27384 5152 0 chany_bottom_out[19]
rlabel metal2 5656 31920 5656 31920 0 chany_bottom_out[1]
rlabel metal3 27860 5320 27860 5320 0 chany_bottom_out[2]
rlabel metal2 3640 30464 3640 30464 0 chany_bottom_out[3]
rlabel metal2 25368 5040 25368 5040 0 chany_bottom_out[5]
rlabel metal2 3472 31920 3472 31920 0 chany_bottom_out[6]
rlabel metal2 3808 29400 3808 29400 0 chany_bottom_out[7]
rlabel metal2 12152 30730 12152 30730 0 chany_bottom_out[9]
rlabel metal2 3080 18256 3080 18256 0 chany_top_in[0]
rlabel metal3 28952 4088 28952 4088 0 chany_top_in[10]
rlabel metal3 4536 29064 4536 29064 0 chany_top_in[12]
rlabel metal2 26096 14616 26096 14616 0 chany_top_in[13]
rlabel metal2 10752 31920 10752 31920 0 chany_top_in[14]
rlabel metal3 30296 10696 30296 10696 0 chany_top_in[16]
rlabel metal3 19096 30184 19096 30184 0 chany_top_in[17]
rlabel metal3 28616 6608 28616 6608 0 chany_top_in[18]
rlabel metal3 24976 5208 24976 5208 0 chany_top_in[1]
rlabel metal3 2702 26936 2702 26936 0 chany_top_in[2]
rlabel metal2 22400 6440 22400 6440 0 chany_top_in[4]
rlabel metal2 4872 30268 4872 30268 0 chany_top_in[5]
rlabel metal2 18984 13328 18984 13328 0 chany_top_in[6]
rlabel metal2 11368 31920 11368 31920 0 chany_top_in[8]
rlabel metal3 1302 22904 1302 22904 0 chany_top_in[9]
rlabel metal3 1358 5432 1358 5432 0 chany_top_out[10]
rlabel metal2 28280 2310 28280 2310 0 chany_top_out[11]
rlabel metal3 12824 29624 12824 29624 0 chany_top_out[13]
rlabel metal2 7448 2058 7448 2058 0 chany_top_out[14]
rlabel metal3 2058 4760 2058 4760 0 chany_top_out[15]
rlabel metal3 854 32984 854 32984 0 chany_top_out[17]
rlabel metal2 28000 29624 28000 29624 0 chany_top_out[18]
rlabel metal3 1358 25592 1358 25592 0 chany_top_out[19]
rlabel metal2 14784 27160 14784 27160 0 chany_top_out[1]
rlabel metal2 21896 29288 21896 29288 0 chany_top_out[2]
rlabel metal2 27608 2422 27608 2422 0 chany_top_out[3]
rlabel metal3 30492 28616 30492 28616 0 chany_top_out[5]
rlabel metal3 1470 20888 1470 20888 0 chany_top_out[6]
rlabel metal3 1470 22232 1470 22232 0 chany_top_out[7]
rlabel metal2 1400 31066 1400 31066 0 chany_top_out[9]
rlabel metal2 26488 14168 26488 14168 0 clknet_0_prog_clk
rlabel metal2 1848 9296 1848 9296 0 clknet_3_0__leaf_prog_clk
rlabel metal2 20776 7840 20776 7840 0 clknet_3_1__leaf_prog_clk
rlabel metal2 8120 28224 8120 28224 0 clknet_3_2__leaf_prog_clk
rlabel metal3 12936 27048 12936 27048 0 clknet_3_3__leaf_prog_clk
rlabel metal3 22400 8232 22400 8232 0 clknet_3_4__leaf_prog_clk
rlabel metal2 29848 6776 29848 6776 0 clknet_3_5__leaf_prog_clk
rlabel metal2 18536 18480 18536 18480 0 clknet_3_6__leaf_prog_clk
rlabel metal2 28616 28168 28616 28168 0 clknet_3_7__leaf_prog_clk
rlabel metal2 11928 15064 11928 15064 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 2744 9072 2744 9072 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal2 3304 6664 3304 6664 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 3080 10024 3080 10024 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 3080 12376 3080 12376 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 3080 15344 3080 15344 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal3 7448 15400 7448 15400 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal2 10920 13552 10920 13552 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal2 17528 13160 17528 13160 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal2 29512 14616 29512 14616 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal2 31304 12936 31304 12936 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal2 25032 17472 25032 17472 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 14392 17864 14392 17864 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal2 20328 18984 20328 18984 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal2 31192 18648 31192 18648 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal2 31528 19768 31528 19768 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal3 28784 17528 28784 17528 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal3 29120 19208 29120 19208 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal3 29792 18312 29792 18312 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal3 31920 24920 31920 24920 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal2 29680 26936 29680 26936 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal2 31584 23800 31584 23800 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal2 22008 21840 22008 21840 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal2 21224 23408 21224 23408 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal2 31080 21112 31080 21112 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal2 25144 21840 25144 21840 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal2 31304 28560 31304 28560 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal2 20552 13552 20552 13552 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal3 22064 12264 22064 12264 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal2 27944 14728 27944 14728 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal3 28056 15960 28056 15960 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal2 25704 15176 25704 15176 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal2 31528 11816 31528 11816 0 mem_right_track_0.DFFR_0_.D
rlabel metal2 26600 26096 26600 26096 0 mem_right_track_0.DFFR_0_.Q
rlabel metal3 22512 25704 22512 25704 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 19656 23128 19656 23128 0 mem_right_track_10.DFFR_0_.D
rlabel metal2 21000 24136 21000 24136 0 mem_right_track_10.DFFR_0_.Q
rlabel metal3 18200 24920 18200 24920 0 mem_right_track_10.DFFR_1_.Q
rlabel metal2 3080 24136 3080 24136 0 mem_right_track_12.DFFR_0_.Q
rlabel metal2 8120 21784 8120 21784 0 mem_right_track_12.DFFR_1_.Q
rlabel metal2 2856 21056 2856 21056 0 mem_right_track_14.DFFR_0_.Q
rlabel metal2 3192 21616 3192 21616 0 mem_right_track_14.DFFR_1_.Q
rlabel metal2 12264 21560 12264 21560 0 mem_right_track_16.DFFR_0_.Q
rlabel metal2 10920 20048 10920 20048 0 mem_right_track_16.DFFR_1_.Q
rlabel metal3 17696 20104 17696 20104 0 mem_right_track_18.DFFR_0_.Q
rlabel metal2 14504 19600 14504 19600 0 mem_right_track_18.DFFR_1_.Q
rlabel metal2 17080 26488 17080 26488 0 mem_right_track_2.DFFR_0_.Q
rlabel metal2 19768 27944 19768 27944 0 mem_right_track_2.DFFR_1_.Q
rlabel metal3 24640 26376 24640 26376 0 mem_right_track_2.DFFR_2_.Q
rlabel metal3 25704 27944 25704 27944 0 mem_right_track_2.DFFR_3_.Q
rlabel metal2 30296 28392 30296 28392 0 mem_right_track_2.DFFR_4_.Q
rlabel metal2 22848 28392 22848 28392 0 mem_right_track_2.DFFR_5_.Q
rlabel metal2 2744 19432 2744 19432 0 mem_right_track_20.DFFR_0_.Q
rlabel metal2 9016 18984 9016 18984 0 mem_right_track_20.DFFR_1_.Q
rlabel metal2 1568 17080 1568 17080 0 mem_right_track_22.DFFR_0_.Q
rlabel metal2 1624 14728 1624 14728 0 mem_right_track_22.DFFR_1_.Q
rlabel metal2 7000 15960 7000 15960 0 mem_right_track_24.DFFR_0_.Q
rlabel metal2 5432 17304 5432 17304 0 mem_right_track_24.DFFR_1_.Q
rlabel metal2 11088 17416 11088 17416 0 mem_right_track_26.DFFR_0_.Q
rlabel metal2 9464 19376 9464 19376 0 mem_right_track_26.DFFR_1_.Q
rlabel metal2 15848 15512 15848 15512 0 mem_right_track_28.DFFR_0_.Q
rlabel metal2 8792 27608 8792 27608 0 mem_right_track_4.DFFR_0_.Q
rlabel metal3 10024 26992 10024 26992 0 mem_right_track_4.DFFR_1_.Q
rlabel metal2 10584 29456 10584 29456 0 mem_right_track_4.DFFR_2_.Q
rlabel metal2 17080 29176 17080 29176 0 mem_right_track_4.DFFR_3_.Q
rlabel metal3 21112 28840 21112 28840 0 mem_right_track_4.DFFR_4_.Q
rlabel metal2 8680 30016 8680 30016 0 mem_right_track_4.DFFR_5_.Q
rlabel metal2 3080 28840 3080 28840 0 mem_right_track_6.DFFR_0_.Q
rlabel metal2 3080 27272 3080 27272 0 mem_right_track_6.DFFR_1_.Q
rlabel metal3 6160 26376 6160 26376 0 mem_right_track_6.DFFR_2_.Q
rlabel metal2 7952 25592 7952 25592 0 mem_right_track_6.DFFR_3_.Q
rlabel metal2 12936 24136 12936 24136 0 mem_right_track_6.DFFR_4_.Q
rlabel metal3 15204 24808 15204 24808 0 mem_right_track_6.DFFR_5_.Q
rlabel metal2 17136 24136 17136 24136 0 mem_right_track_8.DFFR_0_.Q
rlabel metal3 2128 3416 2128 3416 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 18984 3976 18984 3976 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 3080 6440 3080 6440 0 mem_top_track_0.DFFR_2_.Q
rlabel metal2 10024 4928 10024 4928 0 mem_top_track_0.DFFR_3_.Q
rlabel metal2 10136 4648 10136 4648 0 mem_top_track_0.DFFR_4_.Q
rlabel metal2 14280 4536 14280 4536 0 mem_top_track_0.DFFR_5_.Q
rlabel metal3 17864 4424 17864 4424 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 18200 5936 18200 5936 0 mem_top_track_0.DFFR_7_.Q
rlabel metal2 12264 7336 12264 7336 0 mem_top_track_16.DFFR_0_.D
rlabel metal2 12936 8456 12936 8456 0 mem_top_track_16.DFFR_0_.Q
rlabel metal2 16408 6272 16408 6272 0 mem_top_track_16.DFFR_1_.Q
rlabel metal3 18200 8120 18200 8120 0 mem_top_track_16.DFFR_2_.Q
rlabel metal3 23464 8848 23464 8848 0 mem_top_track_16.DFFR_3_.Q
rlabel metal3 23072 7336 23072 7336 0 mem_top_track_16.DFFR_4_.Q
rlabel metal2 25032 8232 25032 8232 0 mem_top_track_16.DFFR_5_.Q
rlabel metal3 29176 8120 29176 8120 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 25032 7000 25032 7000 0 mem_top_track_24.DFFR_1_.Q
rlabel metal2 28168 4760 28168 4760 0 mem_top_track_24.DFFR_2_.Q
rlabel metal2 28392 6832 28392 6832 0 mem_top_track_24.DFFR_3_.Q
rlabel metal2 19040 10024 19040 10024 0 mem_top_track_24.DFFR_4_.Q
rlabel metal3 22792 10696 22792 10696 0 mem_top_track_24.DFFR_5_.Q
rlabel metal3 28112 9688 28112 9688 0 mem_top_track_32.DFFR_0_.Q
rlabel metal3 28168 11256 28168 11256 0 mem_top_track_32.DFFR_1_.Q
rlabel metal3 30520 5880 30520 5880 0 mem_top_track_32.DFFR_2_.Q
rlabel metal2 31528 6888 31528 6888 0 mem_top_track_32.DFFR_3_.Q
rlabel metal3 30296 6664 30296 6664 0 mem_top_track_32.DFFR_4_.Q
rlabel metal3 21672 5992 21672 5992 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 16744 6888 16744 6888 0 mem_top_track_8.DFFR_1_.Q
rlabel metal2 3976 8400 3976 8400 0 mem_top_track_8.DFFR_2_.Q
rlabel metal2 7560 4088 7560 4088 0 mem_top_track_8.DFFR_3_.Q
rlabel metal2 7784 5824 7784 5824 0 mem_top_track_8.DFFR_4_.Q
rlabel metal2 4760 4424 4760 4424 0 net1
rlabel metal2 22568 16352 22568 16352 0 net10
rlabel metal2 16632 27832 16632 27832 0 net100
rlabel metal2 15400 17696 15400 17696 0 net101
rlabel metal2 25816 16800 25816 16800 0 net102
rlabel metal2 4200 21112 4200 21112 0 net103
rlabel metal2 30296 8372 30296 8372 0 net104
rlabel metal2 2352 9016 2352 9016 0 net105
rlabel metal2 14840 14952 14840 14952 0 net106
rlabel metal2 16520 23968 16520 23968 0 net107
rlabel metal2 30632 19656 30632 19656 0 net108
rlabel metal2 17640 19544 17640 19544 0 net109
rlabel metal2 17752 13440 17752 13440 0 net11
rlabel metal2 11760 15288 11760 15288 0 net110
rlabel metal2 29064 29064 29064 29064 0 net111
rlabel metal2 28280 11480 28280 11480 0 net112
rlabel metal2 22568 29344 22568 29344 0 net113
rlabel metal2 9128 28784 9128 28784 0 net114
rlabel metal3 23352 17752 23352 17752 0 net115
rlabel metal2 17808 5880 17808 5880 0 net116
rlabel metal3 18984 8960 18984 8960 0 net117
rlabel metal2 23016 21728 23016 21728 0 net118
rlabel metal2 11144 5040 11144 5040 0 net119
rlabel metal2 8624 27944 8624 27944 0 net12
rlabel metal2 11704 8176 11704 8176 0 net120
rlabel metal2 22904 12880 22904 12880 0 net121
rlabel metal2 18648 11872 18648 11872 0 net122
rlabel metal3 8960 14840 8960 14840 0 net123
rlabel metal3 30016 25816 30016 25816 0 net124
rlabel metal2 4088 16520 4088 16520 0 net125
rlabel metal2 13832 27496 13832 27496 0 net126
rlabel metal2 24248 23968 24248 23968 0 net127
rlabel metal2 21896 7504 21896 7504 0 net128
rlabel metal3 4200 13048 4200 13048 0 net129
rlabel metal3 18368 3528 18368 3528 0 net13
rlabel metal2 21952 11368 21952 11368 0 net130
rlabel metal3 24388 19208 24388 19208 0 net131
rlabel metal3 24360 14952 24360 14952 0 net132
rlabel metal2 4200 25816 4200 25816 0 net133
rlabel metal2 28280 21504 28280 21504 0 net134
rlabel metal2 22904 25424 22904 25424 0 net135
rlabel metal2 3808 11480 3808 11480 0 net136
rlabel metal2 16296 7784 16296 7784 0 net137
rlabel metal2 4088 6720 4088 6720 0 net138
rlabel metal2 11928 13384 11928 13384 0 net139
rlabel metal2 3640 6328 3640 6328 0 net14
rlabel metal2 11816 25704 11816 25704 0 net140
rlabel metal3 20328 28280 20328 28280 0 net141
rlabel metal2 4088 19264 4088 19264 0 net142
rlabel metal2 9912 8064 9912 8064 0 net143
rlabel metal2 3976 17696 3976 17696 0 net144
rlabel metal2 5096 7336 5096 7336 0 net145
rlabel metal2 15176 4648 15176 4648 0 net146
rlabel metal3 29512 5208 29512 5208 0 net147
rlabel metal2 3976 16128 3976 16128 0 net148
rlabel metal2 25256 27384 25256 27384 0 net149
rlabel metal2 31752 9520 31752 9520 0 net15
rlabel metal2 19096 19152 19096 19152 0 net150
rlabel metal2 2184 7896 2184 7896 0 net151
rlabel metal2 11928 26040 11928 26040 0 net152
rlabel metal2 3192 27776 3192 27776 0 net153
rlabel metal2 4088 22008 4088 22008 0 net154
rlabel metal2 4088 9520 4088 9520 0 net155
rlabel metal3 5768 28728 5768 28728 0 net156
rlabel metal2 25816 18480 25816 18480 0 net157
rlabel metal2 4088 23576 4088 23576 0 net158
rlabel metal2 27776 25480 27776 25480 0 net159
rlabel metal2 16352 12376 16352 12376 0 net16
rlabel metal3 23688 26152 23688 26152 0 net160
rlabel metal2 13272 4200 13272 4200 0 net161
rlabel metal2 15400 6440 15400 6440 0 net162
rlabel metal3 24976 6776 24976 6776 0 net163
rlabel metal3 29288 7784 29288 7784 0 net164
rlabel metal2 8456 15988 8456 15988 0 net165
rlabel metal2 11144 3640 11144 3640 0 net166
rlabel metal3 29176 14056 29176 14056 0 net167
rlabel metal2 11032 19040 11032 19040 0 net168
rlabel metal2 18088 5432 18088 5432 0 net169
rlabel metal2 2072 7112 2072 7112 0 net17
rlabel metal2 16464 16072 16464 16072 0 net170
rlabel metal2 26824 10808 26824 10808 0 net171
rlabel metal2 17864 24752 17864 24752 0 net172
rlabel metal3 29904 14168 29904 14168 0 net173
rlabel metal2 6104 8904 6104 8904 0 net174
rlabel metal2 4088 20440 4088 20440 0 net175
rlabel metal3 5040 26264 5040 26264 0 net176
rlabel metal2 17416 14504 17416 14504 0 net177
rlabel metal2 11592 29456 11592 29456 0 net178
rlabel metal2 8120 23576 8120 23576 0 net179
rlabel metal2 23016 16856 23016 16856 0 net18
rlabel metal2 7448 29848 7448 29848 0 net180
rlabel metal2 23240 6608 23240 6608 0 net181
rlabel metal2 22680 15344 22680 15344 0 net182
rlabel metal2 28168 22400 28168 22400 0 net183
rlabel metal2 27160 5264 27160 5264 0 net184
rlabel metal3 16352 27720 16352 27720 0 net185
rlabel metal2 11928 19208 11928 19208 0 net186
rlabel metal2 28952 5432 28952 5432 0 net187
rlabel metal2 11928 28672 11928 28672 0 net188
rlabel metal2 15512 7896 15512 7896 0 net189
rlabel metal2 20776 14112 20776 14112 0 net19
rlabel metal2 23240 19880 23240 19880 0 net190
rlabel metal2 4760 20440 4760 20440 0 net191
rlabel metal2 29288 29288 29288 29288 0 net192
rlabel metal2 3976 11200 3976 11200 0 net193
rlabel metal2 30128 6776 30128 6776 0 net194
rlabel metal2 30184 27804 30184 27804 0 net195
rlabel metal2 4816 16856 4816 16856 0 net196
rlabel metal2 26712 24528 26712 24528 0 net197
rlabel metal2 3864 4648 3864 4648 0 net198
rlabel metal3 26264 7448 26264 7448 0 net199
rlabel metal2 2296 26992 2296 26992 0 net2
rlabel metal2 17752 9352 17752 9352 0 net20
rlabel metal2 15176 26068 15176 26068 0 net200
rlabel metal3 22932 21560 22932 21560 0 net201
rlabel metal2 24528 14616 24528 14616 0 net202
rlabel metal3 1792 15848 1792 15848 0 net21
rlabel metal2 18760 6216 18760 6216 0 net22
rlabel metal2 17584 12152 17584 12152 0 net23
rlabel metal2 17752 19376 17752 19376 0 net24
rlabel metal2 2632 21672 2632 21672 0 net25
rlabel metal3 22736 11256 22736 11256 0 net26
rlabel metal2 19656 29960 19656 29960 0 net27
rlabel metal2 28616 3640 28616 3640 0 net28
rlabel metal2 22792 4648 22792 4648 0 net29
rlabel metal3 23632 9576 23632 9576 0 net3
rlabel metal2 2296 7000 2296 7000 0 net30
rlabel metal2 26264 4872 26264 4872 0 net31
rlabel metal2 17416 16632 17416 16632 0 net32
rlabel metal3 2716 20776 2716 20776 0 net33
rlabel metal2 2184 26152 2184 26152 0 net34
rlabel metal2 2072 10248 2072 10248 0 net35
rlabel metal2 9016 29288 9016 29288 0 net36
rlabel metal2 32200 24136 32200 24136 0 net37
rlabel metal2 25592 3976 25592 3976 0 net38
rlabel metal2 6832 17416 6832 17416 0 net39
rlabel metal2 2296 11368 2296 11368 0 net4
rlabel metal3 22232 21784 22232 21784 0 net40
rlabel metal3 6944 16744 6944 16744 0 net41
rlabel metal2 2968 29848 2968 29848 0 net42
rlabel metal2 24584 7672 24584 7672 0 net43
rlabel metal2 7112 29960 7112 29960 0 net44
rlabel metal2 27104 28392 27104 28392 0 net45
rlabel metal2 7336 28784 7336 28784 0 net46
rlabel metal3 31584 29288 31584 29288 0 net47
rlabel metal2 17976 23772 17976 23772 0 net48
rlabel metal2 28392 3864 28392 3864 0 net49
rlabel metal2 2072 29456 2072 29456 0 net5
rlabel metal2 6888 23520 6888 23520 0 net50
rlabel metal2 23128 4816 23128 4816 0 net51
rlabel metal2 2688 21000 2688 21000 0 net52
rlabel metal2 26040 4704 26040 4704 0 net53
rlabel metal2 9520 17080 9520 17080 0 net54
rlabel metal2 2296 21336 2296 21336 0 net55
rlabel metal2 2408 26040 2408 26040 0 net56
rlabel metal2 17192 6804 17192 6804 0 net57
rlabel metal2 22792 3864 22792 3864 0 net58
rlabel metal2 2296 29008 2296 29008 0 net59
rlabel metal3 10920 3416 10920 3416 0 net6
rlabel metal2 8232 3416 8232 3416 0 net60
rlabel metal2 16296 10024 16296 10024 0 net61
rlabel metal2 4256 29288 4256 29288 0 net62
rlabel metal2 19208 19264 19208 19264 0 net63
rlabel metal2 17416 14112 17416 14112 0 net64
rlabel metal3 12320 26936 12320 26936 0 net65
rlabel metal2 8960 28056 8960 28056 0 net66
rlabel metal2 20272 3416 20272 3416 0 net67
rlabel metal3 24528 14392 24528 14392 0 net68
rlabel metal2 12096 15960 12096 15960 0 net69
rlabel metal2 16520 9744 16520 9744 0 net7
rlabel metal2 2968 24640 2968 24640 0 net70
rlabel metal2 20440 14672 20440 14672 0 net71
rlabel metal3 32690 30296 32690 30296 0 net72
rlabel metal3 8288 3304 8288 3304 0 net73
rlabel metal2 32200 3584 32200 3584 0 net74
rlabel metal2 7672 30772 7672 30772 0 net75
rlabel metal2 29176 30212 29176 30212 0 net76
rlabel metal3 5936 4872 5936 4872 0 net77
rlabel metal2 32088 7392 32088 7392 0 net78
rlabel metal2 27608 31738 27608 31738 0 net79
rlabel metal3 23856 3416 23856 3416 0 net8
rlabel metal2 6104 30506 6104 30506 0 net80
rlabel metal3 6510 2744 6510 2744 0 net81
rlabel metal3 31346 27608 31346 27608 0 net82
rlabel metal2 4984 21168 4984 21168 0 net83
rlabel metal3 2142 2072 2142 2072 0 net84
rlabel metal2 5768 29120 5768 29120 0 net85
rlabel metal2 4816 28392 4816 28392 0 net86
rlabel metal2 26936 2086 26936 2086 0 net87
rlabel metal2 28280 31682 28280 31682 0 net88
rlabel metal2 18984 29624 18984 29624 0 net89
rlabel metal2 2072 8624 2072 8624 0 net9
rlabel metal2 32200 25480 32200 25480 0 net90
rlabel metal3 6888 28280 6888 28280 0 net91
rlabel metal2 32144 6440 32144 6440 0 net92
rlabel metal2 32256 28952 32256 28952 0 net93
rlabel metal2 784 31920 784 31920 0 net94
rlabel metal2 3416 30128 3416 30128 0 net95
rlabel metal3 2478 28280 2478 28280 0 net96
rlabel metal2 22904 2030 22904 2030 0 net97
rlabel metal2 3080 21952 3080 21952 0 net98
rlabel metal2 17752 28952 17752 28952 0 net99
rlabel metal2 10136 28952 10136 28952 0 pReset
rlabel metal2 16800 17080 16800 17080 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 34000 34000
<< end >>
